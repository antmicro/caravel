magic
tech sky130A
magscale 1 2
timestamp 1612197717
<< obsli1 >>
rect 949 2159 398820 497777
<< obsm1 >>
rect 382 1232 398820 497808
<< metal2 >>
rect 1674 499200 1730 500000
rect 5078 499200 5134 500000
rect 8574 499200 8630 500000
rect 12070 499200 12126 500000
rect 15566 499200 15622 500000
rect 19062 499200 19118 500000
rect 22466 499200 22522 500000
rect 25962 499200 26018 500000
rect 29458 499200 29514 500000
rect 32954 499200 33010 500000
rect 36450 499200 36506 500000
rect 39854 499200 39910 500000
rect 43350 499200 43406 500000
rect 46846 499200 46902 500000
rect 50342 499200 50398 500000
rect 53838 499200 53894 500000
rect 57242 499200 57298 500000
rect 60738 499200 60794 500000
rect 64234 499200 64290 500000
rect 67730 499200 67786 500000
rect 71226 499200 71282 500000
rect 74630 499200 74686 500000
rect 78126 499200 78182 500000
rect 81622 499200 81678 500000
rect 85118 499200 85174 500000
rect 88614 499200 88670 500000
rect 92110 499200 92166 500000
rect 95514 499200 95570 500000
rect 99010 499200 99066 500000
rect 102506 499200 102562 500000
rect 106002 499200 106058 500000
rect 109498 499200 109554 500000
rect 112902 499200 112958 500000
rect 116398 499200 116454 500000
rect 119894 499200 119950 500000
rect 123390 499200 123446 500000
rect 126886 499200 126942 500000
rect 130290 499200 130346 500000
rect 133786 499200 133842 500000
rect 137282 499200 137338 500000
rect 140778 499200 140834 500000
rect 144274 499200 144330 500000
rect 147678 499200 147734 500000
rect 151174 499200 151230 500000
rect 154670 499200 154726 500000
rect 158166 499200 158222 500000
rect 161662 499200 161718 500000
rect 165158 499200 165214 500000
rect 168562 499200 168618 500000
rect 172058 499200 172114 500000
rect 175554 499200 175610 500000
rect 179050 499200 179106 500000
rect 182546 499200 182602 500000
rect 185950 499200 186006 500000
rect 189446 499200 189502 500000
rect 192942 499200 192998 500000
rect 196438 499200 196494 500000
rect 199934 499200 199990 500000
rect 203338 499200 203394 500000
rect 206834 499200 206890 500000
rect 210330 499200 210386 500000
rect 213826 499200 213882 500000
rect 217322 499200 217378 500000
rect 220726 499200 220782 500000
rect 224222 499200 224278 500000
rect 227718 499200 227774 500000
rect 231214 499200 231270 500000
rect 234710 499200 234766 500000
rect 238114 499200 238170 500000
rect 241610 499200 241666 500000
rect 245106 499200 245162 500000
rect 248602 499200 248658 500000
rect 252098 499200 252154 500000
rect 255594 499200 255650 500000
rect 258998 499200 259054 500000
rect 262494 499200 262550 500000
rect 265990 499200 266046 500000
rect 269486 499200 269542 500000
rect 272982 499200 273038 500000
rect 276386 499200 276442 500000
rect 279882 499200 279938 500000
rect 283378 499200 283434 500000
rect 286874 499200 286930 500000
rect 290370 499200 290426 500000
rect 293774 499200 293830 500000
rect 297270 499200 297326 500000
rect 300766 499200 300822 500000
rect 304262 499200 304318 500000
rect 307758 499200 307814 500000
rect 311162 499200 311218 500000
rect 314658 499200 314714 500000
rect 318154 499200 318210 500000
rect 321650 499200 321706 500000
rect 325146 499200 325202 500000
rect 328642 499200 328698 500000
rect 332046 499200 332102 500000
rect 335542 499200 335598 500000
rect 339038 499200 339094 500000
rect 342534 499200 342590 500000
rect 346030 499200 346086 500000
rect 349434 499200 349490 500000
rect 352930 499200 352986 500000
rect 356426 499200 356482 500000
rect 359922 499200 359978 500000
rect 363418 499200 363474 500000
rect 366822 499200 366878 500000
rect 370318 499200 370374 500000
rect 373814 499200 373870 500000
rect 377310 499200 377366 500000
rect 380806 499200 380862 500000
rect 384210 499200 384266 500000
rect 387706 499200 387762 500000
rect 391202 499200 391258 500000
rect 394698 499200 394754 500000
rect 398194 499200 398250 500000
rect 386 0 442 800
rect 1122 0 1178 800
rect 1950 0 2006 800
rect 2778 0 2834 800
rect 3606 0 3662 800
rect 4434 0 4490 800
rect 5170 0 5226 800
rect 5998 0 6054 800
rect 6826 0 6882 800
rect 7654 0 7710 800
rect 8482 0 8538 800
rect 9310 0 9366 800
rect 10046 0 10102 800
rect 10874 0 10930 800
rect 11702 0 11758 800
rect 12530 0 12586 800
rect 13358 0 13414 800
rect 14094 0 14150 800
rect 14922 0 14978 800
rect 15750 0 15806 800
rect 16578 0 16634 800
rect 17406 0 17462 800
rect 18234 0 18290 800
rect 18970 0 19026 800
rect 19798 0 19854 800
rect 20626 0 20682 800
rect 21454 0 21510 800
rect 22282 0 22338 800
rect 23018 0 23074 800
rect 23846 0 23902 800
rect 24674 0 24730 800
rect 25502 0 25558 800
rect 26330 0 26386 800
rect 27158 0 27214 800
rect 27894 0 27950 800
rect 28722 0 28778 800
rect 29550 0 29606 800
rect 30378 0 30434 800
rect 31206 0 31262 800
rect 31942 0 31998 800
rect 32770 0 32826 800
rect 33598 0 33654 800
rect 34426 0 34482 800
rect 35254 0 35310 800
rect 36082 0 36138 800
rect 36818 0 36874 800
rect 37646 0 37702 800
rect 38474 0 38530 800
rect 39302 0 39358 800
rect 40130 0 40186 800
rect 40866 0 40922 800
rect 41694 0 41750 800
rect 42522 0 42578 800
rect 43350 0 43406 800
rect 44178 0 44234 800
rect 45006 0 45062 800
rect 45742 0 45798 800
rect 46570 0 46626 800
rect 47398 0 47454 800
rect 48226 0 48282 800
rect 49054 0 49110 800
rect 49790 0 49846 800
rect 50618 0 50674 800
rect 51446 0 51502 800
rect 52274 0 52330 800
rect 53102 0 53158 800
rect 53930 0 53986 800
rect 54666 0 54722 800
rect 55494 0 55550 800
rect 56322 0 56378 800
rect 57150 0 57206 800
rect 57978 0 58034 800
rect 58806 0 58862 800
rect 59542 0 59598 800
rect 60370 0 60426 800
rect 61198 0 61254 800
rect 62026 0 62082 800
rect 62854 0 62910 800
rect 63590 0 63646 800
rect 64418 0 64474 800
rect 65246 0 65302 800
rect 66074 0 66130 800
rect 66902 0 66958 800
rect 67730 0 67786 800
rect 68466 0 68522 800
rect 69294 0 69350 800
rect 70122 0 70178 800
rect 70950 0 71006 800
rect 71778 0 71834 800
rect 72514 0 72570 800
rect 73342 0 73398 800
rect 74170 0 74226 800
rect 74998 0 75054 800
rect 75826 0 75882 800
rect 76654 0 76710 800
rect 77390 0 77446 800
rect 78218 0 78274 800
rect 79046 0 79102 800
rect 79874 0 79930 800
rect 80702 0 80758 800
rect 81438 0 81494 800
rect 82266 0 82322 800
rect 83094 0 83150 800
rect 83922 0 83978 800
rect 84750 0 84806 800
rect 85578 0 85634 800
rect 86314 0 86370 800
rect 87142 0 87198 800
rect 87970 0 88026 800
rect 88798 0 88854 800
rect 89626 0 89682 800
rect 90362 0 90418 800
rect 91190 0 91246 800
rect 92018 0 92074 800
rect 92846 0 92902 800
rect 93674 0 93730 800
rect 94502 0 94558 800
rect 95238 0 95294 800
rect 96066 0 96122 800
rect 96894 0 96950 800
rect 97722 0 97778 800
rect 98550 0 98606 800
rect 99286 0 99342 800
rect 100114 0 100170 800
rect 100942 0 100998 800
rect 101770 0 101826 800
rect 102598 0 102654 800
rect 103426 0 103482 800
rect 104162 0 104218 800
rect 104990 0 105046 800
rect 105818 0 105874 800
rect 106646 0 106702 800
rect 107474 0 107530 800
rect 108210 0 108266 800
rect 109038 0 109094 800
rect 109866 0 109922 800
rect 110694 0 110750 800
rect 111522 0 111578 800
rect 112350 0 112406 800
rect 113086 0 113142 800
rect 113914 0 113970 800
rect 114742 0 114798 800
rect 115570 0 115626 800
rect 116398 0 116454 800
rect 117226 0 117282 800
rect 117962 0 118018 800
rect 118790 0 118846 800
rect 119618 0 119674 800
rect 120446 0 120502 800
rect 121274 0 121330 800
rect 122010 0 122066 800
rect 122838 0 122894 800
rect 123666 0 123722 800
rect 124494 0 124550 800
rect 125322 0 125378 800
rect 126150 0 126206 800
rect 126886 0 126942 800
rect 127714 0 127770 800
rect 128542 0 128598 800
rect 129370 0 129426 800
rect 130198 0 130254 800
rect 130934 0 130990 800
rect 131762 0 131818 800
rect 132590 0 132646 800
rect 133418 0 133474 800
rect 134246 0 134302 800
rect 135074 0 135130 800
rect 135810 0 135866 800
rect 136638 0 136694 800
rect 137466 0 137522 800
rect 138294 0 138350 800
rect 139122 0 139178 800
rect 139858 0 139914 800
rect 140686 0 140742 800
rect 141514 0 141570 800
rect 142342 0 142398 800
rect 143170 0 143226 800
rect 143998 0 144054 800
rect 144734 0 144790 800
rect 145562 0 145618 800
rect 146390 0 146446 800
rect 147218 0 147274 800
rect 148046 0 148102 800
rect 148782 0 148838 800
rect 149610 0 149666 800
rect 150438 0 150494 800
rect 151266 0 151322 800
rect 152094 0 152150 800
rect 152922 0 152978 800
rect 153658 0 153714 800
rect 154486 0 154542 800
rect 155314 0 155370 800
rect 156142 0 156198 800
rect 156970 0 157026 800
rect 157706 0 157762 800
rect 158534 0 158590 800
rect 159362 0 159418 800
rect 160190 0 160246 800
rect 161018 0 161074 800
rect 161846 0 161902 800
rect 162582 0 162638 800
rect 163410 0 163466 800
rect 164238 0 164294 800
rect 165066 0 165122 800
rect 165894 0 165950 800
rect 166630 0 166686 800
rect 167458 0 167514 800
rect 168286 0 168342 800
rect 169114 0 169170 800
rect 169942 0 169998 800
rect 170770 0 170826 800
rect 171506 0 171562 800
rect 172334 0 172390 800
rect 173162 0 173218 800
rect 173990 0 174046 800
rect 174818 0 174874 800
rect 175646 0 175702 800
rect 176382 0 176438 800
rect 177210 0 177266 800
rect 178038 0 178094 800
rect 178866 0 178922 800
rect 179694 0 179750 800
rect 180430 0 180486 800
rect 181258 0 181314 800
rect 182086 0 182142 800
rect 182914 0 182970 800
rect 183742 0 183798 800
rect 184570 0 184626 800
rect 185306 0 185362 800
rect 186134 0 186190 800
rect 186962 0 187018 800
rect 187790 0 187846 800
rect 188618 0 188674 800
rect 189354 0 189410 800
rect 190182 0 190238 800
rect 191010 0 191066 800
rect 191838 0 191894 800
rect 192666 0 192722 800
rect 193494 0 193550 800
rect 194230 0 194286 800
rect 195058 0 195114 800
rect 195886 0 195942 800
rect 196714 0 196770 800
rect 197542 0 197598 800
rect 198278 0 198334 800
rect 199106 0 199162 800
rect 199934 0 199990 800
rect 200762 0 200818 800
rect 201590 0 201646 800
rect 202418 0 202474 800
rect 203154 0 203210 800
rect 203982 0 204038 800
rect 204810 0 204866 800
rect 205638 0 205694 800
rect 206466 0 206522 800
rect 207202 0 207258 800
rect 208030 0 208086 800
rect 208858 0 208914 800
rect 209686 0 209742 800
rect 210514 0 210570 800
rect 211342 0 211398 800
rect 212078 0 212134 800
rect 212906 0 212962 800
rect 213734 0 213790 800
rect 214562 0 214618 800
rect 215390 0 215446 800
rect 216126 0 216182 800
rect 216954 0 217010 800
rect 217782 0 217838 800
rect 218610 0 218666 800
rect 219438 0 219494 800
rect 220266 0 220322 800
rect 221002 0 221058 800
rect 221830 0 221886 800
rect 222658 0 222714 800
rect 223486 0 223542 800
rect 224314 0 224370 800
rect 225050 0 225106 800
rect 225878 0 225934 800
rect 226706 0 226762 800
rect 227534 0 227590 800
rect 228362 0 228418 800
rect 229190 0 229246 800
rect 229926 0 229982 800
rect 230754 0 230810 800
rect 231582 0 231638 800
rect 232410 0 232466 800
rect 233238 0 233294 800
rect 234066 0 234122 800
rect 234802 0 234858 800
rect 235630 0 235686 800
rect 236458 0 236514 800
rect 237286 0 237342 800
rect 238114 0 238170 800
rect 238850 0 238906 800
rect 239678 0 239734 800
rect 240506 0 240562 800
rect 241334 0 241390 800
rect 242162 0 242218 800
rect 242990 0 243046 800
rect 243726 0 243782 800
rect 244554 0 244610 800
rect 245382 0 245438 800
rect 246210 0 246266 800
rect 247038 0 247094 800
rect 247774 0 247830 800
rect 248602 0 248658 800
rect 249430 0 249486 800
rect 250258 0 250314 800
rect 251086 0 251142 800
rect 251914 0 251970 800
rect 252650 0 252706 800
rect 253478 0 253534 800
rect 254306 0 254362 800
rect 255134 0 255190 800
rect 255962 0 256018 800
rect 256698 0 256754 800
rect 257526 0 257582 800
rect 258354 0 258410 800
rect 259182 0 259238 800
rect 260010 0 260066 800
rect 260838 0 260894 800
rect 261574 0 261630 800
rect 262402 0 262458 800
rect 263230 0 263286 800
rect 264058 0 264114 800
rect 264886 0 264942 800
rect 265622 0 265678 800
rect 266450 0 266506 800
rect 267278 0 267334 800
rect 268106 0 268162 800
rect 268934 0 268990 800
rect 269762 0 269818 800
rect 270498 0 270554 800
rect 271326 0 271382 800
rect 272154 0 272210 800
rect 272982 0 273038 800
rect 273810 0 273866 800
rect 274546 0 274602 800
rect 275374 0 275430 800
rect 276202 0 276258 800
rect 277030 0 277086 800
rect 277858 0 277914 800
rect 278686 0 278742 800
rect 279422 0 279478 800
rect 280250 0 280306 800
rect 281078 0 281134 800
rect 281906 0 281962 800
rect 282734 0 282790 800
rect 283470 0 283526 800
rect 284298 0 284354 800
rect 285126 0 285182 800
rect 285954 0 286010 800
rect 286782 0 286838 800
rect 287610 0 287666 800
rect 288346 0 288402 800
rect 289174 0 289230 800
rect 290002 0 290058 800
rect 290830 0 290886 800
rect 291658 0 291714 800
rect 292486 0 292542 800
rect 293222 0 293278 800
rect 294050 0 294106 800
rect 294878 0 294934 800
rect 295706 0 295762 800
rect 296534 0 296590 800
rect 297270 0 297326 800
rect 298098 0 298154 800
rect 298926 0 298982 800
rect 299754 0 299810 800
rect 300582 0 300638 800
rect 301410 0 301466 800
rect 302146 0 302202 800
rect 302974 0 303030 800
rect 303802 0 303858 800
rect 304630 0 304686 800
rect 305458 0 305514 800
rect 306194 0 306250 800
rect 307022 0 307078 800
rect 307850 0 307906 800
rect 308678 0 308734 800
rect 309506 0 309562 800
rect 310334 0 310390 800
rect 311070 0 311126 800
rect 311898 0 311954 800
rect 312726 0 312782 800
rect 313554 0 313610 800
rect 314382 0 314438 800
rect 315118 0 315174 800
rect 315946 0 316002 800
rect 316774 0 316830 800
rect 317602 0 317658 800
rect 318430 0 318486 800
rect 319258 0 319314 800
rect 319994 0 320050 800
rect 320822 0 320878 800
rect 321650 0 321706 800
rect 322478 0 322534 800
rect 323306 0 323362 800
rect 324042 0 324098 800
rect 324870 0 324926 800
rect 325698 0 325754 800
rect 326526 0 326582 800
rect 327354 0 327410 800
rect 328182 0 328238 800
rect 328918 0 328974 800
rect 329746 0 329802 800
rect 330574 0 330630 800
rect 331402 0 331458 800
rect 332230 0 332286 800
rect 332966 0 333022 800
rect 333794 0 333850 800
rect 334622 0 334678 800
rect 335450 0 335506 800
rect 336278 0 336334 800
rect 337106 0 337162 800
rect 337842 0 337898 800
rect 338670 0 338726 800
rect 339498 0 339554 800
rect 340326 0 340382 800
rect 341154 0 341210 800
rect 341890 0 341946 800
rect 342718 0 342774 800
rect 343546 0 343602 800
rect 344374 0 344430 800
rect 345202 0 345258 800
rect 346030 0 346086 800
rect 346766 0 346822 800
rect 347594 0 347650 800
rect 348422 0 348478 800
rect 349250 0 349306 800
rect 350078 0 350134 800
rect 350906 0 350962 800
rect 351642 0 351698 800
rect 352470 0 352526 800
rect 353298 0 353354 800
rect 354126 0 354182 800
rect 354954 0 355010 800
rect 355690 0 355746 800
rect 356518 0 356574 800
rect 357346 0 357402 800
rect 358174 0 358230 800
rect 359002 0 359058 800
rect 359830 0 359886 800
rect 360566 0 360622 800
rect 361394 0 361450 800
rect 362222 0 362278 800
rect 363050 0 363106 800
rect 363878 0 363934 800
rect 364614 0 364670 800
rect 365442 0 365498 800
rect 366270 0 366326 800
rect 367098 0 367154 800
rect 367926 0 367982 800
rect 368754 0 368810 800
rect 369490 0 369546 800
rect 370318 0 370374 800
rect 371146 0 371202 800
rect 371974 0 372030 800
rect 372802 0 372858 800
rect 373538 0 373594 800
rect 374366 0 374422 800
rect 375194 0 375250 800
rect 376022 0 376078 800
rect 376850 0 376906 800
rect 377678 0 377734 800
rect 378414 0 378470 800
rect 379242 0 379298 800
rect 380070 0 380126 800
rect 380898 0 380954 800
rect 381726 0 381782 800
rect 382462 0 382518 800
rect 383290 0 383346 800
rect 384118 0 384174 800
rect 384946 0 385002 800
rect 385774 0 385830 800
rect 386602 0 386658 800
rect 387338 0 387394 800
rect 388166 0 388222 800
rect 388994 0 389050 800
rect 389822 0 389878 800
rect 390650 0 390706 800
rect 391386 0 391442 800
rect 392214 0 392270 800
rect 393042 0 393098 800
rect 393870 0 393926 800
rect 394698 0 394754 800
rect 395526 0 395582 800
rect 396262 0 396318 800
rect 397090 0 397146 800
rect 397918 0 397974 800
rect 398746 0 398802 800
rect 399574 0 399630 800
<< obsm2 >>
rect 388 499144 1618 499200
rect 1786 499144 5022 499200
rect 5190 499144 8518 499200
rect 8686 499144 12014 499200
rect 12182 499144 15510 499200
rect 15678 499144 19006 499200
rect 19174 499144 22410 499200
rect 22578 499144 25906 499200
rect 26074 499144 29402 499200
rect 29570 499144 32898 499200
rect 33066 499144 36394 499200
rect 36562 499144 39798 499200
rect 39966 499144 43294 499200
rect 43462 499144 46790 499200
rect 46958 499144 50286 499200
rect 50454 499144 53782 499200
rect 53950 499144 57186 499200
rect 57354 499144 60682 499200
rect 60850 499144 64178 499200
rect 64346 499144 67674 499200
rect 67842 499144 71170 499200
rect 71338 499144 74574 499200
rect 74742 499144 78070 499200
rect 78238 499144 81566 499200
rect 81734 499144 85062 499200
rect 85230 499144 88558 499200
rect 88726 499144 92054 499200
rect 92222 499144 95458 499200
rect 95626 499144 98954 499200
rect 99122 499144 102450 499200
rect 102618 499144 105946 499200
rect 106114 499144 109442 499200
rect 109610 499144 112846 499200
rect 113014 499144 116342 499200
rect 116510 499144 119838 499200
rect 120006 499144 123334 499200
rect 123502 499144 126830 499200
rect 126998 499144 130234 499200
rect 130402 499144 133730 499200
rect 133898 499144 137226 499200
rect 137394 499144 140722 499200
rect 140890 499144 144218 499200
rect 144386 499144 147622 499200
rect 147790 499144 151118 499200
rect 151286 499144 154614 499200
rect 154782 499144 158110 499200
rect 158278 499144 161606 499200
rect 161774 499144 165102 499200
rect 165270 499144 168506 499200
rect 168674 499144 172002 499200
rect 172170 499144 175498 499200
rect 175666 499144 178994 499200
rect 179162 499144 182490 499200
rect 182658 499144 185894 499200
rect 186062 499144 189390 499200
rect 189558 499144 192886 499200
rect 193054 499144 196382 499200
rect 196550 499144 199878 499200
rect 200046 499144 203282 499200
rect 203450 499144 206778 499200
rect 206946 499144 210274 499200
rect 210442 499144 213770 499200
rect 213938 499144 217266 499200
rect 217434 499144 220670 499200
rect 220838 499144 224166 499200
rect 224334 499144 227662 499200
rect 227830 499144 231158 499200
rect 231326 499144 234654 499200
rect 234822 499144 238058 499200
rect 238226 499144 241554 499200
rect 241722 499144 245050 499200
rect 245218 499144 248546 499200
rect 248714 499144 252042 499200
rect 252210 499144 255538 499200
rect 255706 499144 258942 499200
rect 259110 499144 262438 499200
rect 262606 499144 265934 499200
rect 266102 499144 269430 499200
rect 269598 499144 272926 499200
rect 273094 499144 276330 499200
rect 276498 499144 279826 499200
rect 279994 499144 283322 499200
rect 283490 499144 286818 499200
rect 286986 499144 290314 499200
rect 290482 499144 293718 499200
rect 293886 499144 297214 499200
rect 297382 499144 300710 499200
rect 300878 499144 304206 499200
rect 304374 499144 307702 499200
rect 307870 499144 311106 499200
rect 311274 499144 314602 499200
rect 314770 499144 318098 499200
rect 318266 499144 321594 499200
rect 321762 499144 325090 499200
rect 325258 499144 328586 499200
rect 328754 499144 331990 499200
rect 332158 499144 335486 499200
rect 335654 499144 338982 499200
rect 339150 499144 342478 499200
rect 342646 499144 345974 499200
rect 346142 499144 349378 499200
rect 349546 499144 352874 499200
rect 353042 499144 356370 499200
rect 356538 499144 359866 499200
rect 360034 499144 363362 499200
rect 363530 499144 366766 499200
rect 366934 499144 370262 499200
rect 370430 499144 373758 499200
rect 373926 499144 377254 499200
rect 377422 499144 380750 499200
rect 380918 499144 384154 499200
rect 384322 499144 387650 499200
rect 387818 499144 391146 499200
rect 391314 499144 394642 499200
rect 394810 499144 396316 499200
rect 388 856 396316 499144
rect 498 800 1066 856
rect 1234 800 1894 856
rect 2062 800 2722 856
rect 2890 800 3550 856
rect 3718 800 4378 856
rect 4546 800 5114 856
rect 5282 800 5942 856
rect 6110 800 6770 856
rect 6938 800 7598 856
rect 7766 800 8426 856
rect 8594 800 9254 856
rect 9422 800 9990 856
rect 10158 800 10818 856
rect 10986 800 11646 856
rect 11814 800 12474 856
rect 12642 800 13302 856
rect 13470 800 14038 856
rect 14206 800 14866 856
rect 15034 800 15694 856
rect 15862 800 16522 856
rect 16690 800 17350 856
rect 17518 800 18178 856
rect 18346 800 18914 856
rect 19082 800 19742 856
rect 19910 800 20570 856
rect 20738 800 21398 856
rect 21566 800 22226 856
rect 22394 800 22962 856
rect 23130 800 23790 856
rect 23958 800 24618 856
rect 24786 800 25446 856
rect 25614 800 26274 856
rect 26442 800 27102 856
rect 27270 800 27838 856
rect 28006 800 28666 856
rect 28834 800 29494 856
rect 29662 800 30322 856
rect 30490 800 31150 856
rect 31318 800 31886 856
rect 32054 800 32714 856
rect 32882 800 33542 856
rect 33710 800 34370 856
rect 34538 800 35198 856
rect 35366 800 36026 856
rect 36194 800 36762 856
rect 36930 800 37590 856
rect 37758 800 38418 856
rect 38586 800 39246 856
rect 39414 800 40074 856
rect 40242 800 40810 856
rect 40978 800 41638 856
rect 41806 800 42466 856
rect 42634 800 43294 856
rect 43462 800 44122 856
rect 44290 800 44950 856
rect 45118 800 45686 856
rect 45854 800 46514 856
rect 46682 800 47342 856
rect 47510 800 48170 856
rect 48338 800 48998 856
rect 49166 800 49734 856
rect 49902 800 50562 856
rect 50730 800 51390 856
rect 51558 800 52218 856
rect 52386 800 53046 856
rect 53214 800 53874 856
rect 54042 800 54610 856
rect 54778 800 55438 856
rect 55606 800 56266 856
rect 56434 800 57094 856
rect 57262 800 57922 856
rect 58090 800 58750 856
rect 58918 800 59486 856
rect 59654 800 60314 856
rect 60482 800 61142 856
rect 61310 800 61970 856
rect 62138 800 62798 856
rect 62966 800 63534 856
rect 63702 800 64362 856
rect 64530 800 65190 856
rect 65358 800 66018 856
rect 66186 800 66846 856
rect 67014 800 67674 856
rect 67842 800 68410 856
rect 68578 800 69238 856
rect 69406 800 70066 856
rect 70234 800 70894 856
rect 71062 800 71722 856
rect 71890 800 72458 856
rect 72626 800 73286 856
rect 73454 800 74114 856
rect 74282 800 74942 856
rect 75110 800 75770 856
rect 75938 800 76598 856
rect 76766 800 77334 856
rect 77502 800 78162 856
rect 78330 800 78990 856
rect 79158 800 79818 856
rect 79986 800 80646 856
rect 80814 800 81382 856
rect 81550 800 82210 856
rect 82378 800 83038 856
rect 83206 800 83866 856
rect 84034 800 84694 856
rect 84862 800 85522 856
rect 85690 800 86258 856
rect 86426 800 87086 856
rect 87254 800 87914 856
rect 88082 800 88742 856
rect 88910 800 89570 856
rect 89738 800 90306 856
rect 90474 800 91134 856
rect 91302 800 91962 856
rect 92130 800 92790 856
rect 92958 800 93618 856
rect 93786 800 94446 856
rect 94614 800 95182 856
rect 95350 800 96010 856
rect 96178 800 96838 856
rect 97006 800 97666 856
rect 97834 800 98494 856
rect 98662 800 99230 856
rect 99398 800 100058 856
rect 100226 800 100886 856
rect 101054 800 101714 856
rect 101882 800 102542 856
rect 102710 800 103370 856
rect 103538 800 104106 856
rect 104274 800 104934 856
rect 105102 800 105762 856
rect 105930 800 106590 856
rect 106758 800 107418 856
rect 107586 800 108154 856
rect 108322 800 108982 856
rect 109150 800 109810 856
rect 109978 800 110638 856
rect 110806 800 111466 856
rect 111634 800 112294 856
rect 112462 800 113030 856
rect 113198 800 113858 856
rect 114026 800 114686 856
rect 114854 800 115514 856
rect 115682 800 116342 856
rect 116510 800 117170 856
rect 117338 800 117906 856
rect 118074 800 118734 856
rect 118902 800 119562 856
rect 119730 800 120390 856
rect 120558 800 121218 856
rect 121386 800 121954 856
rect 122122 800 122782 856
rect 122950 800 123610 856
rect 123778 800 124438 856
rect 124606 800 125266 856
rect 125434 800 126094 856
rect 126262 800 126830 856
rect 126998 800 127658 856
rect 127826 800 128486 856
rect 128654 800 129314 856
rect 129482 800 130142 856
rect 130310 800 130878 856
rect 131046 800 131706 856
rect 131874 800 132534 856
rect 132702 800 133362 856
rect 133530 800 134190 856
rect 134358 800 135018 856
rect 135186 800 135754 856
rect 135922 800 136582 856
rect 136750 800 137410 856
rect 137578 800 138238 856
rect 138406 800 139066 856
rect 139234 800 139802 856
rect 139970 800 140630 856
rect 140798 800 141458 856
rect 141626 800 142286 856
rect 142454 800 143114 856
rect 143282 800 143942 856
rect 144110 800 144678 856
rect 144846 800 145506 856
rect 145674 800 146334 856
rect 146502 800 147162 856
rect 147330 800 147990 856
rect 148158 800 148726 856
rect 148894 800 149554 856
rect 149722 800 150382 856
rect 150550 800 151210 856
rect 151378 800 152038 856
rect 152206 800 152866 856
rect 153034 800 153602 856
rect 153770 800 154430 856
rect 154598 800 155258 856
rect 155426 800 156086 856
rect 156254 800 156914 856
rect 157082 800 157650 856
rect 157818 800 158478 856
rect 158646 800 159306 856
rect 159474 800 160134 856
rect 160302 800 160962 856
rect 161130 800 161790 856
rect 161958 800 162526 856
rect 162694 800 163354 856
rect 163522 800 164182 856
rect 164350 800 165010 856
rect 165178 800 165838 856
rect 166006 800 166574 856
rect 166742 800 167402 856
rect 167570 800 168230 856
rect 168398 800 169058 856
rect 169226 800 169886 856
rect 170054 800 170714 856
rect 170882 800 171450 856
rect 171618 800 172278 856
rect 172446 800 173106 856
rect 173274 800 173934 856
rect 174102 800 174762 856
rect 174930 800 175590 856
rect 175758 800 176326 856
rect 176494 800 177154 856
rect 177322 800 177982 856
rect 178150 800 178810 856
rect 178978 800 179638 856
rect 179806 800 180374 856
rect 180542 800 181202 856
rect 181370 800 182030 856
rect 182198 800 182858 856
rect 183026 800 183686 856
rect 183854 800 184514 856
rect 184682 800 185250 856
rect 185418 800 186078 856
rect 186246 800 186906 856
rect 187074 800 187734 856
rect 187902 800 188562 856
rect 188730 800 189298 856
rect 189466 800 190126 856
rect 190294 800 190954 856
rect 191122 800 191782 856
rect 191950 800 192610 856
rect 192778 800 193438 856
rect 193606 800 194174 856
rect 194342 800 195002 856
rect 195170 800 195830 856
rect 195998 800 196658 856
rect 196826 800 197486 856
rect 197654 800 198222 856
rect 198390 800 199050 856
rect 199218 800 199878 856
rect 200046 800 200706 856
rect 200874 800 201534 856
rect 201702 800 202362 856
rect 202530 800 203098 856
rect 203266 800 203926 856
rect 204094 800 204754 856
rect 204922 800 205582 856
rect 205750 800 206410 856
rect 206578 800 207146 856
rect 207314 800 207974 856
rect 208142 800 208802 856
rect 208970 800 209630 856
rect 209798 800 210458 856
rect 210626 800 211286 856
rect 211454 800 212022 856
rect 212190 800 212850 856
rect 213018 800 213678 856
rect 213846 800 214506 856
rect 214674 800 215334 856
rect 215502 800 216070 856
rect 216238 800 216898 856
rect 217066 800 217726 856
rect 217894 800 218554 856
rect 218722 800 219382 856
rect 219550 800 220210 856
rect 220378 800 220946 856
rect 221114 800 221774 856
rect 221942 800 222602 856
rect 222770 800 223430 856
rect 223598 800 224258 856
rect 224426 800 224994 856
rect 225162 800 225822 856
rect 225990 800 226650 856
rect 226818 800 227478 856
rect 227646 800 228306 856
rect 228474 800 229134 856
rect 229302 800 229870 856
rect 230038 800 230698 856
rect 230866 800 231526 856
rect 231694 800 232354 856
rect 232522 800 233182 856
rect 233350 800 234010 856
rect 234178 800 234746 856
rect 234914 800 235574 856
rect 235742 800 236402 856
rect 236570 800 237230 856
rect 237398 800 238058 856
rect 238226 800 238794 856
rect 238962 800 239622 856
rect 239790 800 240450 856
rect 240618 800 241278 856
rect 241446 800 242106 856
rect 242274 800 242934 856
rect 243102 800 243670 856
rect 243838 800 244498 856
rect 244666 800 245326 856
rect 245494 800 246154 856
rect 246322 800 246982 856
rect 247150 800 247718 856
rect 247886 800 248546 856
rect 248714 800 249374 856
rect 249542 800 250202 856
rect 250370 800 251030 856
rect 251198 800 251858 856
rect 252026 800 252594 856
rect 252762 800 253422 856
rect 253590 800 254250 856
rect 254418 800 255078 856
rect 255246 800 255906 856
rect 256074 800 256642 856
rect 256810 800 257470 856
rect 257638 800 258298 856
rect 258466 800 259126 856
rect 259294 800 259954 856
rect 260122 800 260782 856
rect 260950 800 261518 856
rect 261686 800 262346 856
rect 262514 800 263174 856
rect 263342 800 264002 856
rect 264170 800 264830 856
rect 264998 800 265566 856
rect 265734 800 266394 856
rect 266562 800 267222 856
rect 267390 800 268050 856
rect 268218 800 268878 856
rect 269046 800 269706 856
rect 269874 800 270442 856
rect 270610 800 271270 856
rect 271438 800 272098 856
rect 272266 800 272926 856
rect 273094 800 273754 856
rect 273922 800 274490 856
rect 274658 800 275318 856
rect 275486 800 276146 856
rect 276314 800 276974 856
rect 277142 800 277802 856
rect 277970 800 278630 856
rect 278798 800 279366 856
rect 279534 800 280194 856
rect 280362 800 281022 856
rect 281190 800 281850 856
rect 282018 800 282678 856
rect 282846 800 283414 856
rect 283582 800 284242 856
rect 284410 800 285070 856
rect 285238 800 285898 856
rect 286066 800 286726 856
rect 286894 800 287554 856
rect 287722 800 288290 856
rect 288458 800 289118 856
rect 289286 800 289946 856
rect 290114 800 290774 856
rect 290942 800 291602 856
rect 291770 800 292430 856
rect 292598 800 293166 856
rect 293334 800 293994 856
rect 294162 800 294822 856
rect 294990 800 295650 856
rect 295818 800 296478 856
rect 296646 800 297214 856
rect 297382 800 298042 856
rect 298210 800 298870 856
rect 299038 800 299698 856
rect 299866 800 300526 856
rect 300694 800 301354 856
rect 301522 800 302090 856
rect 302258 800 302918 856
rect 303086 800 303746 856
rect 303914 800 304574 856
rect 304742 800 305402 856
rect 305570 800 306138 856
rect 306306 800 306966 856
rect 307134 800 307794 856
rect 307962 800 308622 856
rect 308790 800 309450 856
rect 309618 800 310278 856
rect 310446 800 311014 856
rect 311182 800 311842 856
rect 312010 800 312670 856
rect 312838 800 313498 856
rect 313666 800 314326 856
rect 314494 800 315062 856
rect 315230 800 315890 856
rect 316058 800 316718 856
rect 316886 800 317546 856
rect 317714 800 318374 856
rect 318542 800 319202 856
rect 319370 800 319938 856
rect 320106 800 320766 856
rect 320934 800 321594 856
rect 321762 800 322422 856
rect 322590 800 323250 856
rect 323418 800 323986 856
rect 324154 800 324814 856
rect 324982 800 325642 856
rect 325810 800 326470 856
rect 326638 800 327298 856
rect 327466 800 328126 856
rect 328294 800 328862 856
rect 329030 800 329690 856
rect 329858 800 330518 856
rect 330686 800 331346 856
rect 331514 800 332174 856
rect 332342 800 332910 856
rect 333078 800 333738 856
rect 333906 800 334566 856
rect 334734 800 335394 856
rect 335562 800 336222 856
rect 336390 800 337050 856
rect 337218 800 337786 856
rect 337954 800 338614 856
rect 338782 800 339442 856
rect 339610 800 340270 856
rect 340438 800 341098 856
rect 341266 800 341834 856
rect 342002 800 342662 856
rect 342830 800 343490 856
rect 343658 800 344318 856
rect 344486 800 345146 856
rect 345314 800 345974 856
rect 346142 800 346710 856
rect 346878 800 347538 856
rect 347706 800 348366 856
rect 348534 800 349194 856
rect 349362 800 350022 856
rect 350190 800 350850 856
rect 351018 800 351586 856
rect 351754 800 352414 856
rect 352582 800 353242 856
rect 353410 800 354070 856
rect 354238 800 354898 856
rect 355066 800 355634 856
rect 355802 800 356462 856
rect 356630 800 357290 856
rect 357458 800 358118 856
rect 358286 800 358946 856
rect 359114 800 359774 856
rect 359942 800 360510 856
rect 360678 800 361338 856
rect 361506 800 362166 856
rect 362334 800 362994 856
rect 363162 800 363822 856
rect 363990 800 364558 856
rect 364726 800 365386 856
rect 365554 800 366214 856
rect 366382 800 367042 856
rect 367210 800 367870 856
rect 368038 800 368698 856
rect 368866 800 369434 856
rect 369602 800 370262 856
rect 370430 800 371090 856
rect 371258 800 371918 856
rect 372086 800 372746 856
rect 372914 800 373482 856
rect 373650 800 374310 856
rect 374478 800 375138 856
rect 375306 800 375966 856
rect 376134 800 376794 856
rect 376962 800 377622 856
rect 377790 800 378358 856
rect 378526 800 379186 856
rect 379354 800 380014 856
rect 380182 800 380842 856
rect 381010 800 381670 856
rect 381838 800 382406 856
rect 382574 800 383234 856
rect 383402 800 384062 856
rect 384230 800 384890 856
rect 385058 800 385718 856
rect 385886 800 386546 856
rect 386714 800 387282 856
rect 387450 800 388110 856
rect 388278 800 388938 856
rect 389106 800 389766 856
rect 389934 800 390594 856
rect 390762 800 391330 856
rect 391498 800 392158 856
rect 392326 800 392986 856
rect 393154 800 393814 856
rect 393982 800 394642 856
rect 394810 800 395470 856
rect 395638 800 396206 856
<< metal3 >>
rect 0 416440 800 416560
rect 0 249840 800 249960
rect 0 83240 800 83360
rect 399200 249976 400000 250096
<< obsm3 >>
rect 2037 2143 388528 497793
<< metal4 >>
rect 4208 2128 4528 497808
rect 19568 2128 19888 497808
rect 34928 2128 35248 497808
rect 50288 2128 50608 497808
rect 65648 2128 65968 497808
rect 81008 2128 81328 497808
rect 96368 2128 96688 497808
rect 111728 2128 112048 497808
rect 127088 2128 127408 497808
rect 142448 2128 142768 497808
rect 157808 2128 158128 497808
rect 173168 2128 173488 497808
rect 188528 2128 188848 497808
rect 203888 2128 204208 497808
rect 219248 2128 219568 497808
rect 234608 2128 234928 497808
rect 249968 2128 250288 497808
rect 265328 2128 265648 497808
rect 280688 2128 281008 497808
rect 296048 2128 296368 497808
rect 311408 2128 311728 497808
rect 326768 2128 327088 497808
rect 342128 2128 342448 497808
rect 357488 2128 357808 497808
rect 372848 2128 373168 497808
rect 388208 2128 388528 497808
<< labels >>
rlabel metal2 s 1674 499200 1730 500000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 106002 499200 106058 500000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 116398 499200 116454 500000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 126886 499200 126942 500000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 137282 499200 137338 500000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 147678 499200 147734 500000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 158166 499200 158222 500000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 168562 499200 168618 500000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 179050 499200 179106 500000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 189446 499200 189502 500000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 199934 499200 199990 500000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 12070 499200 12126 500000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 210330 499200 210386 500000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 220726 499200 220782 500000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 231214 499200 231270 500000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 241610 499200 241666 500000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 252098 499200 252154 500000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 262494 499200 262550 500000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 272982 499200 273038 500000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 283378 499200 283434 500000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 293774 499200 293830 500000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 304262 499200 304318 500000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 22466 499200 22522 500000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 314658 499200 314714 500000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 325146 499200 325202 500000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 335542 499200 335598 500000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 346030 499200 346086 500000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 356426 499200 356482 500000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 366822 499200 366878 500000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 377310 499200 377366 500000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 387706 499200 387762 500000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 32954 499200 33010 500000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 43350 499200 43406 500000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 53838 499200 53894 500000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 64234 499200 64290 500000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 74630 499200 74686 500000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 85118 499200 85174 500000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 95514 499200 95570 500000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 5078 499200 5134 500000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 109498 499200 109554 500000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 119894 499200 119950 500000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 130290 499200 130346 500000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 140778 499200 140834 500000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 151174 499200 151230 500000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 161662 499200 161718 500000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 172058 499200 172114 500000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 182546 499200 182602 500000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 192942 499200 192998 500000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 203338 499200 203394 500000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 15566 499200 15622 500000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 213826 499200 213882 500000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 224222 499200 224278 500000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 234710 499200 234766 500000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 245106 499200 245162 500000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 255594 499200 255650 500000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 265990 499200 266046 500000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 276386 499200 276442 500000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 286874 499200 286930 500000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 297270 499200 297326 500000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 307758 499200 307814 500000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 25962 499200 26018 500000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 318154 499200 318210 500000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 328642 499200 328698 500000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 339038 499200 339094 500000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 349434 499200 349490 500000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 359922 499200 359978 500000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 370318 499200 370374 500000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 380806 499200 380862 500000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 391202 499200 391258 500000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 36450 499200 36506 500000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 46846 499200 46902 500000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 57242 499200 57298 500000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 67730 499200 67786 500000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 78126 499200 78182 500000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 88614 499200 88670 500000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 99010 499200 99066 500000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 8574 499200 8630 500000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 112902 499200 112958 500000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 123390 499200 123446 500000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 133786 499200 133842 500000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 144274 499200 144330 500000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 154670 499200 154726 500000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 165158 499200 165214 500000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 175554 499200 175610 500000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 185950 499200 186006 500000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 196438 499200 196494 500000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 206834 499200 206890 500000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 19062 499200 19118 500000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 217322 499200 217378 500000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 227718 499200 227774 500000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 238114 499200 238170 500000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 248602 499200 248658 500000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 258998 499200 259054 500000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 269486 499200 269542 500000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 279882 499200 279938 500000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 290370 499200 290426 500000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 300766 499200 300822 500000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 311162 499200 311218 500000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 29458 499200 29514 500000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 321650 499200 321706 500000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 332046 499200 332102 500000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 342534 499200 342590 500000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 352930 499200 352986 500000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 363418 499200 363474 500000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 373814 499200 373870 500000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 384210 499200 384266 500000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 394698 499200 394754 500000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 39854 499200 39910 500000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 50342 499200 50398 500000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 60738 499200 60794 500000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 71226 499200 71282 500000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 81622 499200 81678 500000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 92110 499200 92166 500000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 102506 499200 102562 500000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 86314 0 86370 800 6 la_data_in[0]
port 115 nsew signal input
rlabel metal2 s 329746 0 329802 800 6 la_data_in[100]
port 116 nsew signal input
rlabel metal2 s 332230 0 332286 800 6 la_data_in[101]
port 117 nsew signal input
rlabel metal2 s 334622 0 334678 800 6 la_data_in[102]
port 118 nsew signal input
rlabel metal2 s 337106 0 337162 800 6 la_data_in[103]
port 119 nsew signal input
rlabel metal2 s 339498 0 339554 800 6 la_data_in[104]
port 120 nsew signal input
rlabel metal2 s 341890 0 341946 800 6 la_data_in[105]
port 121 nsew signal input
rlabel metal2 s 344374 0 344430 800 6 la_data_in[106]
port 122 nsew signal input
rlabel metal2 s 346766 0 346822 800 6 la_data_in[107]
port 123 nsew signal input
rlabel metal2 s 349250 0 349306 800 6 la_data_in[108]
port 124 nsew signal input
rlabel metal2 s 351642 0 351698 800 6 la_data_in[109]
port 125 nsew signal input
rlabel metal2 s 110694 0 110750 800 6 la_data_in[10]
port 126 nsew signal input
rlabel metal2 s 354126 0 354182 800 6 la_data_in[110]
port 127 nsew signal input
rlabel metal2 s 356518 0 356574 800 6 la_data_in[111]
port 128 nsew signal input
rlabel metal2 s 359002 0 359058 800 6 la_data_in[112]
port 129 nsew signal input
rlabel metal2 s 361394 0 361450 800 6 la_data_in[113]
port 130 nsew signal input
rlabel metal2 s 363878 0 363934 800 6 la_data_in[114]
port 131 nsew signal input
rlabel metal2 s 366270 0 366326 800 6 la_data_in[115]
port 132 nsew signal input
rlabel metal2 s 368754 0 368810 800 6 la_data_in[116]
port 133 nsew signal input
rlabel metal2 s 371146 0 371202 800 6 la_data_in[117]
port 134 nsew signal input
rlabel metal2 s 373538 0 373594 800 6 la_data_in[118]
port 135 nsew signal input
rlabel metal2 s 376022 0 376078 800 6 la_data_in[119]
port 136 nsew signal input
rlabel metal2 s 113086 0 113142 800 6 la_data_in[11]
port 137 nsew signal input
rlabel metal2 s 378414 0 378470 800 6 la_data_in[120]
port 138 nsew signal input
rlabel metal2 s 380898 0 380954 800 6 la_data_in[121]
port 139 nsew signal input
rlabel metal2 s 383290 0 383346 800 6 la_data_in[122]
port 140 nsew signal input
rlabel metal2 s 385774 0 385830 800 6 la_data_in[123]
port 141 nsew signal input
rlabel metal2 s 388166 0 388222 800 6 la_data_in[124]
port 142 nsew signal input
rlabel metal2 s 390650 0 390706 800 6 la_data_in[125]
port 143 nsew signal input
rlabel metal2 s 393042 0 393098 800 6 la_data_in[126]
port 144 nsew signal input
rlabel metal2 s 395526 0 395582 800 6 la_data_in[127]
port 145 nsew signal input
rlabel metal2 s 115570 0 115626 800 6 la_data_in[12]
port 146 nsew signal input
rlabel metal2 s 117962 0 118018 800 6 la_data_in[13]
port 147 nsew signal input
rlabel metal2 s 120446 0 120502 800 6 la_data_in[14]
port 148 nsew signal input
rlabel metal2 s 122838 0 122894 800 6 la_data_in[15]
port 149 nsew signal input
rlabel metal2 s 125322 0 125378 800 6 la_data_in[16]
port 150 nsew signal input
rlabel metal2 s 127714 0 127770 800 6 la_data_in[17]
port 151 nsew signal input
rlabel metal2 s 130198 0 130254 800 6 la_data_in[18]
port 152 nsew signal input
rlabel metal2 s 132590 0 132646 800 6 la_data_in[19]
port 153 nsew signal input
rlabel metal2 s 88798 0 88854 800 6 la_data_in[1]
port 154 nsew signal input
rlabel metal2 s 135074 0 135130 800 6 la_data_in[20]
port 155 nsew signal input
rlabel metal2 s 137466 0 137522 800 6 la_data_in[21]
port 156 nsew signal input
rlabel metal2 s 139858 0 139914 800 6 la_data_in[22]
port 157 nsew signal input
rlabel metal2 s 142342 0 142398 800 6 la_data_in[23]
port 158 nsew signal input
rlabel metal2 s 144734 0 144790 800 6 la_data_in[24]
port 159 nsew signal input
rlabel metal2 s 147218 0 147274 800 6 la_data_in[25]
port 160 nsew signal input
rlabel metal2 s 149610 0 149666 800 6 la_data_in[26]
port 161 nsew signal input
rlabel metal2 s 152094 0 152150 800 6 la_data_in[27]
port 162 nsew signal input
rlabel metal2 s 154486 0 154542 800 6 la_data_in[28]
port 163 nsew signal input
rlabel metal2 s 156970 0 157026 800 6 la_data_in[29]
port 164 nsew signal input
rlabel metal2 s 91190 0 91246 800 6 la_data_in[2]
port 165 nsew signal input
rlabel metal2 s 159362 0 159418 800 6 la_data_in[30]
port 166 nsew signal input
rlabel metal2 s 161846 0 161902 800 6 la_data_in[31]
port 167 nsew signal input
rlabel metal2 s 164238 0 164294 800 6 la_data_in[32]
port 168 nsew signal input
rlabel metal2 s 166630 0 166686 800 6 la_data_in[33]
port 169 nsew signal input
rlabel metal2 s 169114 0 169170 800 6 la_data_in[34]
port 170 nsew signal input
rlabel metal2 s 171506 0 171562 800 6 la_data_in[35]
port 171 nsew signal input
rlabel metal2 s 173990 0 174046 800 6 la_data_in[36]
port 172 nsew signal input
rlabel metal2 s 176382 0 176438 800 6 la_data_in[37]
port 173 nsew signal input
rlabel metal2 s 178866 0 178922 800 6 la_data_in[38]
port 174 nsew signal input
rlabel metal2 s 181258 0 181314 800 6 la_data_in[39]
port 175 nsew signal input
rlabel metal2 s 93674 0 93730 800 6 la_data_in[3]
port 176 nsew signal input
rlabel metal2 s 183742 0 183798 800 6 la_data_in[40]
port 177 nsew signal input
rlabel metal2 s 186134 0 186190 800 6 la_data_in[41]
port 178 nsew signal input
rlabel metal2 s 188618 0 188674 800 6 la_data_in[42]
port 179 nsew signal input
rlabel metal2 s 191010 0 191066 800 6 la_data_in[43]
port 180 nsew signal input
rlabel metal2 s 193494 0 193550 800 6 la_data_in[44]
port 181 nsew signal input
rlabel metal2 s 195886 0 195942 800 6 la_data_in[45]
port 182 nsew signal input
rlabel metal2 s 198278 0 198334 800 6 la_data_in[46]
port 183 nsew signal input
rlabel metal2 s 200762 0 200818 800 6 la_data_in[47]
port 184 nsew signal input
rlabel metal2 s 203154 0 203210 800 6 la_data_in[48]
port 185 nsew signal input
rlabel metal2 s 205638 0 205694 800 6 la_data_in[49]
port 186 nsew signal input
rlabel metal2 s 96066 0 96122 800 6 la_data_in[4]
port 187 nsew signal input
rlabel metal2 s 208030 0 208086 800 6 la_data_in[50]
port 188 nsew signal input
rlabel metal2 s 210514 0 210570 800 6 la_data_in[51]
port 189 nsew signal input
rlabel metal2 s 212906 0 212962 800 6 la_data_in[52]
port 190 nsew signal input
rlabel metal2 s 215390 0 215446 800 6 la_data_in[53]
port 191 nsew signal input
rlabel metal2 s 217782 0 217838 800 6 la_data_in[54]
port 192 nsew signal input
rlabel metal2 s 220266 0 220322 800 6 la_data_in[55]
port 193 nsew signal input
rlabel metal2 s 222658 0 222714 800 6 la_data_in[56]
port 194 nsew signal input
rlabel metal2 s 225050 0 225106 800 6 la_data_in[57]
port 195 nsew signal input
rlabel metal2 s 227534 0 227590 800 6 la_data_in[58]
port 196 nsew signal input
rlabel metal2 s 229926 0 229982 800 6 la_data_in[59]
port 197 nsew signal input
rlabel metal2 s 98550 0 98606 800 6 la_data_in[5]
port 198 nsew signal input
rlabel metal2 s 232410 0 232466 800 6 la_data_in[60]
port 199 nsew signal input
rlabel metal2 s 234802 0 234858 800 6 la_data_in[61]
port 200 nsew signal input
rlabel metal2 s 237286 0 237342 800 6 la_data_in[62]
port 201 nsew signal input
rlabel metal2 s 239678 0 239734 800 6 la_data_in[63]
port 202 nsew signal input
rlabel metal2 s 242162 0 242218 800 6 la_data_in[64]
port 203 nsew signal input
rlabel metal2 s 244554 0 244610 800 6 la_data_in[65]
port 204 nsew signal input
rlabel metal2 s 247038 0 247094 800 6 la_data_in[66]
port 205 nsew signal input
rlabel metal2 s 249430 0 249486 800 6 la_data_in[67]
port 206 nsew signal input
rlabel metal2 s 251914 0 251970 800 6 la_data_in[68]
port 207 nsew signal input
rlabel metal2 s 254306 0 254362 800 6 la_data_in[69]
port 208 nsew signal input
rlabel metal2 s 100942 0 100998 800 6 la_data_in[6]
port 209 nsew signal input
rlabel metal2 s 256698 0 256754 800 6 la_data_in[70]
port 210 nsew signal input
rlabel metal2 s 259182 0 259238 800 6 la_data_in[71]
port 211 nsew signal input
rlabel metal2 s 261574 0 261630 800 6 la_data_in[72]
port 212 nsew signal input
rlabel metal2 s 264058 0 264114 800 6 la_data_in[73]
port 213 nsew signal input
rlabel metal2 s 266450 0 266506 800 6 la_data_in[74]
port 214 nsew signal input
rlabel metal2 s 268934 0 268990 800 6 la_data_in[75]
port 215 nsew signal input
rlabel metal2 s 271326 0 271382 800 6 la_data_in[76]
port 216 nsew signal input
rlabel metal2 s 273810 0 273866 800 6 la_data_in[77]
port 217 nsew signal input
rlabel metal2 s 276202 0 276258 800 6 la_data_in[78]
port 218 nsew signal input
rlabel metal2 s 278686 0 278742 800 6 la_data_in[79]
port 219 nsew signal input
rlabel metal2 s 103426 0 103482 800 6 la_data_in[7]
port 220 nsew signal input
rlabel metal2 s 281078 0 281134 800 6 la_data_in[80]
port 221 nsew signal input
rlabel metal2 s 283470 0 283526 800 6 la_data_in[81]
port 222 nsew signal input
rlabel metal2 s 285954 0 286010 800 6 la_data_in[82]
port 223 nsew signal input
rlabel metal2 s 288346 0 288402 800 6 la_data_in[83]
port 224 nsew signal input
rlabel metal2 s 290830 0 290886 800 6 la_data_in[84]
port 225 nsew signal input
rlabel metal2 s 293222 0 293278 800 6 la_data_in[85]
port 226 nsew signal input
rlabel metal2 s 295706 0 295762 800 6 la_data_in[86]
port 227 nsew signal input
rlabel metal2 s 298098 0 298154 800 6 la_data_in[87]
port 228 nsew signal input
rlabel metal2 s 300582 0 300638 800 6 la_data_in[88]
port 229 nsew signal input
rlabel metal2 s 302974 0 303030 800 6 la_data_in[89]
port 230 nsew signal input
rlabel metal2 s 105818 0 105874 800 6 la_data_in[8]
port 231 nsew signal input
rlabel metal2 s 305458 0 305514 800 6 la_data_in[90]
port 232 nsew signal input
rlabel metal2 s 307850 0 307906 800 6 la_data_in[91]
port 233 nsew signal input
rlabel metal2 s 310334 0 310390 800 6 la_data_in[92]
port 234 nsew signal input
rlabel metal2 s 312726 0 312782 800 6 la_data_in[93]
port 235 nsew signal input
rlabel metal2 s 315118 0 315174 800 6 la_data_in[94]
port 236 nsew signal input
rlabel metal2 s 317602 0 317658 800 6 la_data_in[95]
port 237 nsew signal input
rlabel metal2 s 319994 0 320050 800 6 la_data_in[96]
port 238 nsew signal input
rlabel metal2 s 322478 0 322534 800 6 la_data_in[97]
port 239 nsew signal input
rlabel metal2 s 324870 0 324926 800 6 la_data_in[98]
port 240 nsew signal input
rlabel metal2 s 327354 0 327410 800 6 la_data_in[99]
port 241 nsew signal input
rlabel metal2 s 108210 0 108266 800 6 la_data_in[9]
port 242 nsew signal input
rlabel metal2 s 87142 0 87198 800 6 la_data_out[0]
port 243 nsew signal output
rlabel metal2 s 330574 0 330630 800 6 la_data_out[100]
port 244 nsew signal output
rlabel metal2 s 332966 0 333022 800 6 la_data_out[101]
port 245 nsew signal output
rlabel metal2 s 335450 0 335506 800 6 la_data_out[102]
port 246 nsew signal output
rlabel metal2 s 337842 0 337898 800 6 la_data_out[103]
port 247 nsew signal output
rlabel metal2 s 340326 0 340382 800 6 la_data_out[104]
port 248 nsew signal output
rlabel metal2 s 342718 0 342774 800 6 la_data_out[105]
port 249 nsew signal output
rlabel metal2 s 345202 0 345258 800 6 la_data_out[106]
port 250 nsew signal output
rlabel metal2 s 347594 0 347650 800 6 la_data_out[107]
port 251 nsew signal output
rlabel metal2 s 350078 0 350134 800 6 la_data_out[108]
port 252 nsew signal output
rlabel metal2 s 352470 0 352526 800 6 la_data_out[109]
port 253 nsew signal output
rlabel metal2 s 111522 0 111578 800 6 la_data_out[10]
port 254 nsew signal output
rlabel metal2 s 354954 0 355010 800 6 la_data_out[110]
port 255 nsew signal output
rlabel metal2 s 357346 0 357402 800 6 la_data_out[111]
port 256 nsew signal output
rlabel metal2 s 359830 0 359886 800 6 la_data_out[112]
port 257 nsew signal output
rlabel metal2 s 362222 0 362278 800 6 la_data_out[113]
port 258 nsew signal output
rlabel metal2 s 364614 0 364670 800 6 la_data_out[114]
port 259 nsew signal output
rlabel metal2 s 367098 0 367154 800 6 la_data_out[115]
port 260 nsew signal output
rlabel metal2 s 369490 0 369546 800 6 la_data_out[116]
port 261 nsew signal output
rlabel metal2 s 371974 0 372030 800 6 la_data_out[117]
port 262 nsew signal output
rlabel metal2 s 374366 0 374422 800 6 la_data_out[118]
port 263 nsew signal output
rlabel metal2 s 376850 0 376906 800 6 la_data_out[119]
port 264 nsew signal output
rlabel metal2 s 113914 0 113970 800 6 la_data_out[11]
port 265 nsew signal output
rlabel metal2 s 379242 0 379298 800 6 la_data_out[120]
port 266 nsew signal output
rlabel metal2 s 381726 0 381782 800 6 la_data_out[121]
port 267 nsew signal output
rlabel metal2 s 384118 0 384174 800 6 la_data_out[122]
port 268 nsew signal output
rlabel metal2 s 386602 0 386658 800 6 la_data_out[123]
port 269 nsew signal output
rlabel metal2 s 388994 0 389050 800 6 la_data_out[124]
port 270 nsew signal output
rlabel metal2 s 391386 0 391442 800 6 la_data_out[125]
port 271 nsew signal output
rlabel metal2 s 393870 0 393926 800 6 la_data_out[126]
port 272 nsew signal output
rlabel metal2 s 396262 0 396318 800 6 la_data_out[127]
port 273 nsew signal output
rlabel metal2 s 116398 0 116454 800 6 la_data_out[12]
port 274 nsew signal output
rlabel metal2 s 118790 0 118846 800 6 la_data_out[13]
port 275 nsew signal output
rlabel metal2 s 121274 0 121330 800 6 la_data_out[14]
port 276 nsew signal output
rlabel metal2 s 123666 0 123722 800 6 la_data_out[15]
port 277 nsew signal output
rlabel metal2 s 126150 0 126206 800 6 la_data_out[16]
port 278 nsew signal output
rlabel metal2 s 128542 0 128598 800 6 la_data_out[17]
port 279 nsew signal output
rlabel metal2 s 130934 0 130990 800 6 la_data_out[18]
port 280 nsew signal output
rlabel metal2 s 133418 0 133474 800 6 la_data_out[19]
port 281 nsew signal output
rlabel metal2 s 89626 0 89682 800 6 la_data_out[1]
port 282 nsew signal output
rlabel metal2 s 135810 0 135866 800 6 la_data_out[20]
port 283 nsew signal output
rlabel metal2 s 138294 0 138350 800 6 la_data_out[21]
port 284 nsew signal output
rlabel metal2 s 140686 0 140742 800 6 la_data_out[22]
port 285 nsew signal output
rlabel metal2 s 143170 0 143226 800 6 la_data_out[23]
port 286 nsew signal output
rlabel metal2 s 145562 0 145618 800 6 la_data_out[24]
port 287 nsew signal output
rlabel metal2 s 148046 0 148102 800 6 la_data_out[25]
port 288 nsew signal output
rlabel metal2 s 150438 0 150494 800 6 la_data_out[26]
port 289 nsew signal output
rlabel metal2 s 152922 0 152978 800 6 la_data_out[27]
port 290 nsew signal output
rlabel metal2 s 155314 0 155370 800 6 la_data_out[28]
port 291 nsew signal output
rlabel metal2 s 157706 0 157762 800 6 la_data_out[29]
port 292 nsew signal output
rlabel metal2 s 92018 0 92074 800 6 la_data_out[2]
port 293 nsew signal output
rlabel metal2 s 160190 0 160246 800 6 la_data_out[30]
port 294 nsew signal output
rlabel metal2 s 162582 0 162638 800 6 la_data_out[31]
port 295 nsew signal output
rlabel metal2 s 165066 0 165122 800 6 la_data_out[32]
port 296 nsew signal output
rlabel metal2 s 167458 0 167514 800 6 la_data_out[33]
port 297 nsew signal output
rlabel metal2 s 169942 0 169998 800 6 la_data_out[34]
port 298 nsew signal output
rlabel metal2 s 172334 0 172390 800 6 la_data_out[35]
port 299 nsew signal output
rlabel metal2 s 174818 0 174874 800 6 la_data_out[36]
port 300 nsew signal output
rlabel metal2 s 177210 0 177266 800 6 la_data_out[37]
port 301 nsew signal output
rlabel metal2 s 179694 0 179750 800 6 la_data_out[38]
port 302 nsew signal output
rlabel metal2 s 182086 0 182142 800 6 la_data_out[39]
port 303 nsew signal output
rlabel metal2 s 94502 0 94558 800 6 la_data_out[3]
port 304 nsew signal output
rlabel metal2 s 184570 0 184626 800 6 la_data_out[40]
port 305 nsew signal output
rlabel metal2 s 186962 0 187018 800 6 la_data_out[41]
port 306 nsew signal output
rlabel metal2 s 189354 0 189410 800 6 la_data_out[42]
port 307 nsew signal output
rlabel metal2 s 191838 0 191894 800 6 la_data_out[43]
port 308 nsew signal output
rlabel metal2 s 194230 0 194286 800 6 la_data_out[44]
port 309 nsew signal output
rlabel metal2 s 196714 0 196770 800 6 la_data_out[45]
port 310 nsew signal output
rlabel metal2 s 199106 0 199162 800 6 la_data_out[46]
port 311 nsew signal output
rlabel metal2 s 201590 0 201646 800 6 la_data_out[47]
port 312 nsew signal output
rlabel metal2 s 203982 0 204038 800 6 la_data_out[48]
port 313 nsew signal output
rlabel metal2 s 206466 0 206522 800 6 la_data_out[49]
port 314 nsew signal output
rlabel metal2 s 96894 0 96950 800 6 la_data_out[4]
port 315 nsew signal output
rlabel metal2 s 208858 0 208914 800 6 la_data_out[50]
port 316 nsew signal output
rlabel metal2 s 211342 0 211398 800 6 la_data_out[51]
port 317 nsew signal output
rlabel metal2 s 213734 0 213790 800 6 la_data_out[52]
port 318 nsew signal output
rlabel metal2 s 216126 0 216182 800 6 la_data_out[53]
port 319 nsew signal output
rlabel metal2 s 218610 0 218666 800 6 la_data_out[54]
port 320 nsew signal output
rlabel metal2 s 221002 0 221058 800 6 la_data_out[55]
port 321 nsew signal output
rlabel metal2 s 223486 0 223542 800 6 la_data_out[56]
port 322 nsew signal output
rlabel metal2 s 225878 0 225934 800 6 la_data_out[57]
port 323 nsew signal output
rlabel metal2 s 228362 0 228418 800 6 la_data_out[58]
port 324 nsew signal output
rlabel metal2 s 230754 0 230810 800 6 la_data_out[59]
port 325 nsew signal output
rlabel metal2 s 99286 0 99342 800 6 la_data_out[5]
port 326 nsew signal output
rlabel metal2 s 233238 0 233294 800 6 la_data_out[60]
port 327 nsew signal output
rlabel metal2 s 235630 0 235686 800 6 la_data_out[61]
port 328 nsew signal output
rlabel metal2 s 238114 0 238170 800 6 la_data_out[62]
port 329 nsew signal output
rlabel metal2 s 240506 0 240562 800 6 la_data_out[63]
port 330 nsew signal output
rlabel metal2 s 242990 0 243046 800 6 la_data_out[64]
port 331 nsew signal output
rlabel metal2 s 245382 0 245438 800 6 la_data_out[65]
port 332 nsew signal output
rlabel metal2 s 247774 0 247830 800 6 la_data_out[66]
port 333 nsew signal output
rlabel metal2 s 250258 0 250314 800 6 la_data_out[67]
port 334 nsew signal output
rlabel metal2 s 252650 0 252706 800 6 la_data_out[68]
port 335 nsew signal output
rlabel metal2 s 255134 0 255190 800 6 la_data_out[69]
port 336 nsew signal output
rlabel metal2 s 101770 0 101826 800 6 la_data_out[6]
port 337 nsew signal output
rlabel metal2 s 257526 0 257582 800 6 la_data_out[70]
port 338 nsew signal output
rlabel metal2 s 260010 0 260066 800 6 la_data_out[71]
port 339 nsew signal output
rlabel metal2 s 262402 0 262458 800 6 la_data_out[72]
port 340 nsew signal output
rlabel metal2 s 264886 0 264942 800 6 la_data_out[73]
port 341 nsew signal output
rlabel metal2 s 267278 0 267334 800 6 la_data_out[74]
port 342 nsew signal output
rlabel metal2 s 269762 0 269818 800 6 la_data_out[75]
port 343 nsew signal output
rlabel metal2 s 272154 0 272210 800 6 la_data_out[76]
port 344 nsew signal output
rlabel metal2 s 274546 0 274602 800 6 la_data_out[77]
port 345 nsew signal output
rlabel metal2 s 277030 0 277086 800 6 la_data_out[78]
port 346 nsew signal output
rlabel metal2 s 279422 0 279478 800 6 la_data_out[79]
port 347 nsew signal output
rlabel metal2 s 104162 0 104218 800 6 la_data_out[7]
port 348 nsew signal output
rlabel metal2 s 281906 0 281962 800 6 la_data_out[80]
port 349 nsew signal output
rlabel metal2 s 284298 0 284354 800 6 la_data_out[81]
port 350 nsew signal output
rlabel metal2 s 286782 0 286838 800 6 la_data_out[82]
port 351 nsew signal output
rlabel metal2 s 289174 0 289230 800 6 la_data_out[83]
port 352 nsew signal output
rlabel metal2 s 291658 0 291714 800 6 la_data_out[84]
port 353 nsew signal output
rlabel metal2 s 294050 0 294106 800 6 la_data_out[85]
port 354 nsew signal output
rlabel metal2 s 296534 0 296590 800 6 la_data_out[86]
port 355 nsew signal output
rlabel metal2 s 298926 0 298982 800 6 la_data_out[87]
port 356 nsew signal output
rlabel metal2 s 301410 0 301466 800 6 la_data_out[88]
port 357 nsew signal output
rlabel metal2 s 303802 0 303858 800 6 la_data_out[89]
port 358 nsew signal output
rlabel metal2 s 106646 0 106702 800 6 la_data_out[8]
port 359 nsew signal output
rlabel metal2 s 306194 0 306250 800 6 la_data_out[90]
port 360 nsew signal output
rlabel metal2 s 308678 0 308734 800 6 la_data_out[91]
port 361 nsew signal output
rlabel metal2 s 311070 0 311126 800 6 la_data_out[92]
port 362 nsew signal output
rlabel metal2 s 313554 0 313610 800 6 la_data_out[93]
port 363 nsew signal output
rlabel metal2 s 315946 0 316002 800 6 la_data_out[94]
port 364 nsew signal output
rlabel metal2 s 318430 0 318486 800 6 la_data_out[95]
port 365 nsew signal output
rlabel metal2 s 320822 0 320878 800 6 la_data_out[96]
port 366 nsew signal output
rlabel metal2 s 323306 0 323362 800 6 la_data_out[97]
port 367 nsew signal output
rlabel metal2 s 325698 0 325754 800 6 la_data_out[98]
port 368 nsew signal output
rlabel metal2 s 328182 0 328238 800 6 la_data_out[99]
port 369 nsew signal output
rlabel metal2 s 109038 0 109094 800 6 la_data_out[9]
port 370 nsew signal output
rlabel metal2 s 87970 0 88026 800 6 la_oen[0]
port 371 nsew signal input
rlabel metal2 s 331402 0 331458 800 6 la_oen[100]
port 372 nsew signal input
rlabel metal2 s 333794 0 333850 800 6 la_oen[101]
port 373 nsew signal input
rlabel metal2 s 336278 0 336334 800 6 la_oen[102]
port 374 nsew signal input
rlabel metal2 s 338670 0 338726 800 6 la_oen[103]
port 375 nsew signal input
rlabel metal2 s 341154 0 341210 800 6 la_oen[104]
port 376 nsew signal input
rlabel metal2 s 343546 0 343602 800 6 la_oen[105]
port 377 nsew signal input
rlabel metal2 s 346030 0 346086 800 6 la_oen[106]
port 378 nsew signal input
rlabel metal2 s 348422 0 348478 800 6 la_oen[107]
port 379 nsew signal input
rlabel metal2 s 350906 0 350962 800 6 la_oen[108]
port 380 nsew signal input
rlabel metal2 s 353298 0 353354 800 6 la_oen[109]
port 381 nsew signal input
rlabel metal2 s 112350 0 112406 800 6 la_oen[10]
port 382 nsew signal input
rlabel metal2 s 355690 0 355746 800 6 la_oen[110]
port 383 nsew signal input
rlabel metal2 s 358174 0 358230 800 6 la_oen[111]
port 384 nsew signal input
rlabel metal2 s 360566 0 360622 800 6 la_oen[112]
port 385 nsew signal input
rlabel metal2 s 363050 0 363106 800 6 la_oen[113]
port 386 nsew signal input
rlabel metal2 s 365442 0 365498 800 6 la_oen[114]
port 387 nsew signal input
rlabel metal2 s 367926 0 367982 800 6 la_oen[115]
port 388 nsew signal input
rlabel metal2 s 370318 0 370374 800 6 la_oen[116]
port 389 nsew signal input
rlabel metal2 s 372802 0 372858 800 6 la_oen[117]
port 390 nsew signal input
rlabel metal2 s 375194 0 375250 800 6 la_oen[118]
port 391 nsew signal input
rlabel metal2 s 377678 0 377734 800 6 la_oen[119]
port 392 nsew signal input
rlabel metal2 s 114742 0 114798 800 6 la_oen[11]
port 393 nsew signal input
rlabel metal2 s 380070 0 380126 800 6 la_oen[120]
port 394 nsew signal input
rlabel metal2 s 382462 0 382518 800 6 la_oen[121]
port 395 nsew signal input
rlabel metal2 s 384946 0 385002 800 6 la_oen[122]
port 396 nsew signal input
rlabel metal2 s 387338 0 387394 800 6 la_oen[123]
port 397 nsew signal input
rlabel metal2 s 389822 0 389878 800 6 la_oen[124]
port 398 nsew signal input
rlabel metal2 s 392214 0 392270 800 6 la_oen[125]
port 399 nsew signal input
rlabel metal2 s 394698 0 394754 800 6 la_oen[126]
port 400 nsew signal input
rlabel metal2 s 397090 0 397146 800 6 la_oen[127]
port 401 nsew signal input
rlabel metal2 s 117226 0 117282 800 6 la_oen[12]
port 402 nsew signal input
rlabel metal2 s 119618 0 119674 800 6 la_oen[13]
port 403 nsew signal input
rlabel metal2 s 122010 0 122066 800 6 la_oen[14]
port 404 nsew signal input
rlabel metal2 s 124494 0 124550 800 6 la_oen[15]
port 405 nsew signal input
rlabel metal2 s 126886 0 126942 800 6 la_oen[16]
port 406 nsew signal input
rlabel metal2 s 129370 0 129426 800 6 la_oen[17]
port 407 nsew signal input
rlabel metal2 s 131762 0 131818 800 6 la_oen[18]
port 408 nsew signal input
rlabel metal2 s 134246 0 134302 800 6 la_oen[19]
port 409 nsew signal input
rlabel metal2 s 90362 0 90418 800 6 la_oen[1]
port 410 nsew signal input
rlabel metal2 s 136638 0 136694 800 6 la_oen[20]
port 411 nsew signal input
rlabel metal2 s 139122 0 139178 800 6 la_oen[21]
port 412 nsew signal input
rlabel metal2 s 141514 0 141570 800 6 la_oen[22]
port 413 nsew signal input
rlabel metal2 s 143998 0 144054 800 6 la_oen[23]
port 414 nsew signal input
rlabel metal2 s 146390 0 146446 800 6 la_oen[24]
port 415 nsew signal input
rlabel metal2 s 148782 0 148838 800 6 la_oen[25]
port 416 nsew signal input
rlabel metal2 s 151266 0 151322 800 6 la_oen[26]
port 417 nsew signal input
rlabel metal2 s 153658 0 153714 800 6 la_oen[27]
port 418 nsew signal input
rlabel metal2 s 156142 0 156198 800 6 la_oen[28]
port 419 nsew signal input
rlabel metal2 s 158534 0 158590 800 6 la_oen[29]
port 420 nsew signal input
rlabel metal2 s 92846 0 92902 800 6 la_oen[2]
port 421 nsew signal input
rlabel metal2 s 161018 0 161074 800 6 la_oen[30]
port 422 nsew signal input
rlabel metal2 s 163410 0 163466 800 6 la_oen[31]
port 423 nsew signal input
rlabel metal2 s 165894 0 165950 800 6 la_oen[32]
port 424 nsew signal input
rlabel metal2 s 168286 0 168342 800 6 la_oen[33]
port 425 nsew signal input
rlabel metal2 s 170770 0 170826 800 6 la_oen[34]
port 426 nsew signal input
rlabel metal2 s 173162 0 173218 800 6 la_oen[35]
port 427 nsew signal input
rlabel metal2 s 175646 0 175702 800 6 la_oen[36]
port 428 nsew signal input
rlabel metal2 s 178038 0 178094 800 6 la_oen[37]
port 429 nsew signal input
rlabel metal2 s 180430 0 180486 800 6 la_oen[38]
port 430 nsew signal input
rlabel metal2 s 182914 0 182970 800 6 la_oen[39]
port 431 nsew signal input
rlabel metal2 s 95238 0 95294 800 6 la_oen[3]
port 432 nsew signal input
rlabel metal2 s 185306 0 185362 800 6 la_oen[40]
port 433 nsew signal input
rlabel metal2 s 187790 0 187846 800 6 la_oen[41]
port 434 nsew signal input
rlabel metal2 s 190182 0 190238 800 6 la_oen[42]
port 435 nsew signal input
rlabel metal2 s 192666 0 192722 800 6 la_oen[43]
port 436 nsew signal input
rlabel metal2 s 195058 0 195114 800 6 la_oen[44]
port 437 nsew signal input
rlabel metal2 s 197542 0 197598 800 6 la_oen[45]
port 438 nsew signal input
rlabel metal2 s 199934 0 199990 800 6 la_oen[46]
port 439 nsew signal input
rlabel metal2 s 202418 0 202474 800 6 la_oen[47]
port 440 nsew signal input
rlabel metal2 s 204810 0 204866 800 6 la_oen[48]
port 441 nsew signal input
rlabel metal2 s 207202 0 207258 800 6 la_oen[49]
port 442 nsew signal input
rlabel metal2 s 97722 0 97778 800 6 la_oen[4]
port 443 nsew signal input
rlabel metal2 s 209686 0 209742 800 6 la_oen[50]
port 444 nsew signal input
rlabel metal2 s 212078 0 212134 800 6 la_oen[51]
port 445 nsew signal input
rlabel metal2 s 214562 0 214618 800 6 la_oen[52]
port 446 nsew signal input
rlabel metal2 s 216954 0 217010 800 6 la_oen[53]
port 447 nsew signal input
rlabel metal2 s 219438 0 219494 800 6 la_oen[54]
port 448 nsew signal input
rlabel metal2 s 221830 0 221886 800 6 la_oen[55]
port 449 nsew signal input
rlabel metal2 s 224314 0 224370 800 6 la_oen[56]
port 450 nsew signal input
rlabel metal2 s 226706 0 226762 800 6 la_oen[57]
port 451 nsew signal input
rlabel metal2 s 229190 0 229246 800 6 la_oen[58]
port 452 nsew signal input
rlabel metal2 s 231582 0 231638 800 6 la_oen[59]
port 453 nsew signal input
rlabel metal2 s 100114 0 100170 800 6 la_oen[5]
port 454 nsew signal input
rlabel metal2 s 234066 0 234122 800 6 la_oen[60]
port 455 nsew signal input
rlabel metal2 s 236458 0 236514 800 6 la_oen[61]
port 456 nsew signal input
rlabel metal2 s 238850 0 238906 800 6 la_oen[62]
port 457 nsew signal input
rlabel metal2 s 241334 0 241390 800 6 la_oen[63]
port 458 nsew signal input
rlabel metal2 s 243726 0 243782 800 6 la_oen[64]
port 459 nsew signal input
rlabel metal2 s 246210 0 246266 800 6 la_oen[65]
port 460 nsew signal input
rlabel metal2 s 248602 0 248658 800 6 la_oen[66]
port 461 nsew signal input
rlabel metal2 s 251086 0 251142 800 6 la_oen[67]
port 462 nsew signal input
rlabel metal2 s 253478 0 253534 800 6 la_oen[68]
port 463 nsew signal input
rlabel metal2 s 255962 0 256018 800 6 la_oen[69]
port 464 nsew signal input
rlabel metal2 s 102598 0 102654 800 6 la_oen[6]
port 465 nsew signal input
rlabel metal2 s 258354 0 258410 800 6 la_oen[70]
port 466 nsew signal input
rlabel metal2 s 260838 0 260894 800 6 la_oen[71]
port 467 nsew signal input
rlabel metal2 s 263230 0 263286 800 6 la_oen[72]
port 468 nsew signal input
rlabel metal2 s 265622 0 265678 800 6 la_oen[73]
port 469 nsew signal input
rlabel metal2 s 268106 0 268162 800 6 la_oen[74]
port 470 nsew signal input
rlabel metal2 s 270498 0 270554 800 6 la_oen[75]
port 471 nsew signal input
rlabel metal2 s 272982 0 273038 800 6 la_oen[76]
port 472 nsew signal input
rlabel metal2 s 275374 0 275430 800 6 la_oen[77]
port 473 nsew signal input
rlabel metal2 s 277858 0 277914 800 6 la_oen[78]
port 474 nsew signal input
rlabel metal2 s 280250 0 280306 800 6 la_oen[79]
port 475 nsew signal input
rlabel metal2 s 104990 0 105046 800 6 la_oen[7]
port 476 nsew signal input
rlabel metal2 s 282734 0 282790 800 6 la_oen[80]
port 477 nsew signal input
rlabel metal2 s 285126 0 285182 800 6 la_oen[81]
port 478 nsew signal input
rlabel metal2 s 287610 0 287666 800 6 la_oen[82]
port 479 nsew signal input
rlabel metal2 s 290002 0 290058 800 6 la_oen[83]
port 480 nsew signal input
rlabel metal2 s 292486 0 292542 800 6 la_oen[84]
port 481 nsew signal input
rlabel metal2 s 294878 0 294934 800 6 la_oen[85]
port 482 nsew signal input
rlabel metal2 s 297270 0 297326 800 6 la_oen[86]
port 483 nsew signal input
rlabel metal2 s 299754 0 299810 800 6 la_oen[87]
port 484 nsew signal input
rlabel metal2 s 302146 0 302202 800 6 la_oen[88]
port 485 nsew signal input
rlabel metal2 s 304630 0 304686 800 6 la_oen[89]
port 486 nsew signal input
rlabel metal2 s 107474 0 107530 800 6 la_oen[8]
port 487 nsew signal input
rlabel metal2 s 307022 0 307078 800 6 la_oen[90]
port 488 nsew signal input
rlabel metal2 s 309506 0 309562 800 6 la_oen[91]
port 489 nsew signal input
rlabel metal2 s 311898 0 311954 800 6 la_oen[92]
port 490 nsew signal input
rlabel metal2 s 314382 0 314438 800 6 la_oen[93]
port 491 nsew signal input
rlabel metal2 s 316774 0 316830 800 6 la_oen[94]
port 492 nsew signal input
rlabel metal2 s 319258 0 319314 800 6 la_oen[95]
port 493 nsew signal input
rlabel metal2 s 321650 0 321706 800 6 la_oen[96]
port 494 nsew signal input
rlabel metal2 s 324042 0 324098 800 6 la_oen[97]
port 495 nsew signal input
rlabel metal2 s 326526 0 326582 800 6 la_oen[98]
port 496 nsew signal input
rlabel metal2 s 328918 0 328974 800 6 la_oen[99]
port 497 nsew signal input
rlabel metal2 s 109866 0 109922 800 6 la_oen[9]
port 498 nsew signal input
rlabel metal3 s 0 83240 800 83360 6 vccd1
port 499 nsew signal bidirectional
rlabel metal3 s 0 249840 800 249960 6 vccd2
port 500 nsew signal bidirectional
rlabel metal2 s 397918 0 397974 800 6 vdda1
port 501 nsew signal bidirectional
rlabel metal2 s 398194 499200 398250 500000 6 vdda2
port 502 nsew signal bidirectional
rlabel metal3 s 399200 249976 400000 250096 6 vssa1
port 503 nsew signal bidirectional
rlabel metal3 s 0 416440 800 416560 6 vssa2
port 504 nsew signal bidirectional
rlabel metal2 s 398746 0 398802 800 6 vssd1
port 505 nsew signal bidirectional
rlabel metal2 s 399574 0 399630 800 6 vssd2
port 506 nsew signal bidirectional
rlabel metal2 s 386 0 442 800 6 wb_clk_i
port 507 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 wb_rst_i
port 508 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 wbs_ack_o
port 509 nsew signal output
rlabel metal2 s 5170 0 5226 800 6 wbs_adr_i[0]
port 510 nsew signal input
rlabel metal2 s 32770 0 32826 800 6 wbs_adr_i[10]
port 511 nsew signal input
rlabel metal2 s 35254 0 35310 800 6 wbs_adr_i[11]
port 512 nsew signal input
rlabel metal2 s 37646 0 37702 800 6 wbs_adr_i[12]
port 513 nsew signal input
rlabel metal2 s 40130 0 40186 800 6 wbs_adr_i[13]
port 514 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 wbs_adr_i[14]
port 515 nsew signal input
rlabel metal2 s 45006 0 45062 800 6 wbs_adr_i[15]
port 516 nsew signal input
rlabel metal2 s 47398 0 47454 800 6 wbs_adr_i[16]
port 517 nsew signal input
rlabel metal2 s 49790 0 49846 800 6 wbs_adr_i[17]
port 518 nsew signal input
rlabel metal2 s 52274 0 52330 800 6 wbs_adr_i[18]
port 519 nsew signal input
rlabel metal2 s 54666 0 54722 800 6 wbs_adr_i[19]
port 520 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 wbs_adr_i[1]
port 521 nsew signal input
rlabel metal2 s 57150 0 57206 800 6 wbs_adr_i[20]
port 522 nsew signal input
rlabel metal2 s 59542 0 59598 800 6 wbs_adr_i[21]
port 523 nsew signal input
rlabel metal2 s 62026 0 62082 800 6 wbs_adr_i[22]
port 524 nsew signal input
rlabel metal2 s 64418 0 64474 800 6 wbs_adr_i[23]
port 525 nsew signal input
rlabel metal2 s 66902 0 66958 800 6 wbs_adr_i[24]
port 526 nsew signal input
rlabel metal2 s 69294 0 69350 800 6 wbs_adr_i[25]
port 527 nsew signal input
rlabel metal2 s 71778 0 71834 800 6 wbs_adr_i[26]
port 528 nsew signal input
rlabel metal2 s 74170 0 74226 800 6 wbs_adr_i[27]
port 529 nsew signal input
rlabel metal2 s 76654 0 76710 800 6 wbs_adr_i[28]
port 530 nsew signal input
rlabel metal2 s 79046 0 79102 800 6 wbs_adr_i[29]
port 531 nsew signal input
rlabel metal2 s 11702 0 11758 800 6 wbs_adr_i[2]
port 532 nsew signal input
rlabel metal2 s 81438 0 81494 800 6 wbs_adr_i[30]
port 533 nsew signal input
rlabel metal2 s 83922 0 83978 800 6 wbs_adr_i[31]
port 534 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 wbs_adr_i[3]
port 535 nsew signal input
rlabel metal2 s 18234 0 18290 800 6 wbs_adr_i[4]
port 536 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 wbs_adr_i[5]
port 537 nsew signal input
rlabel metal2 s 23018 0 23074 800 6 wbs_adr_i[6]
port 538 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 wbs_adr_i[7]
port 539 nsew signal input
rlabel metal2 s 27894 0 27950 800 6 wbs_adr_i[8]
port 540 nsew signal input
rlabel metal2 s 30378 0 30434 800 6 wbs_adr_i[9]
port 541 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 wbs_cyc_i
port 542 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 wbs_dat_i[0]
port 543 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 wbs_dat_i[10]
port 544 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 wbs_dat_i[11]
port 545 nsew signal input
rlabel metal2 s 38474 0 38530 800 6 wbs_dat_i[12]
port 546 nsew signal input
rlabel metal2 s 40866 0 40922 800 6 wbs_dat_i[13]
port 547 nsew signal input
rlabel metal2 s 43350 0 43406 800 6 wbs_dat_i[14]
port 548 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 wbs_dat_i[15]
port 549 nsew signal input
rlabel metal2 s 48226 0 48282 800 6 wbs_dat_i[16]
port 550 nsew signal input
rlabel metal2 s 50618 0 50674 800 6 wbs_dat_i[17]
port 551 nsew signal input
rlabel metal2 s 53102 0 53158 800 6 wbs_dat_i[18]
port 552 nsew signal input
rlabel metal2 s 55494 0 55550 800 6 wbs_dat_i[19]
port 553 nsew signal input
rlabel metal2 s 9310 0 9366 800 6 wbs_dat_i[1]
port 554 nsew signal input
rlabel metal2 s 57978 0 58034 800 6 wbs_dat_i[20]
port 555 nsew signal input
rlabel metal2 s 60370 0 60426 800 6 wbs_dat_i[21]
port 556 nsew signal input
rlabel metal2 s 62854 0 62910 800 6 wbs_dat_i[22]
port 557 nsew signal input
rlabel metal2 s 65246 0 65302 800 6 wbs_dat_i[23]
port 558 nsew signal input
rlabel metal2 s 67730 0 67786 800 6 wbs_dat_i[24]
port 559 nsew signal input
rlabel metal2 s 70122 0 70178 800 6 wbs_dat_i[25]
port 560 nsew signal input
rlabel metal2 s 72514 0 72570 800 6 wbs_dat_i[26]
port 561 nsew signal input
rlabel metal2 s 74998 0 75054 800 6 wbs_dat_i[27]
port 562 nsew signal input
rlabel metal2 s 77390 0 77446 800 6 wbs_dat_i[28]
port 563 nsew signal input
rlabel metal2 s 79874 0 79930 800 6 wbs_dat_i[29]
port 564 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 wbs_dat_i[2]
port 565 nsew signal input
rlabel metal2 s 82266 0 82322 800 6 wbs_dat_i[30]
port 566 nsew signal input
rlabel metal2 s 84750 0 84806 800 6 wbs_dat_i[31]
port 567 nsew signal input
rlabel metal2 s 15750 0 15806 800 6 wbs_dat_i[3]
port 568 nsew signal input
rlabel metal2 s 18970 0 19026 800 6 wbs_dat_i[4]
port 569 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 wbs_dat_i[5]
port 570 nsew signal input
rlabel metal2 s 23846 0 23902 800 6 wbs_dat_i[6]
port 571 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 wbs_dat_i[7]
port 572 nsew signal input
rlabel metal2 s 28722 0 28778 800 6 wbs_dat_i[8]
port 573 nsew signal input
rlabel metal2 s 31206 0 31262 800 6 wbs_dat_i[9]
port 574 nsew signal input
rlabel metal2 s 6826 0 6882 800 6 wbs_dat_o[0]
port 575 nsew signal output
rlabel metal2 s 34426 0 34482 800 6 wbs_dat_o[10]
port 576 nsew signal output
rlabel metal2 s 36818 0 36874 800 6 wbs_dat_o[11]
port 577 nsew signal output
rlabel metal2 s 39302 0 39358 800 6 wbs_dat_o[12]
port 578 nsew signal output
rlabel metal2 s 41694 0 41750 800 6 wbs_dat_o[13]
port 579 nsew signal output
rlabel metal2 s 44178 0 44234 800 6 wbs_dat_o[14]
port 580 nsew signal output
rlabel metal2 s 46570 0 46626 800 6 wbs_dat_o[15]
port 581 nsew signal output
rlabel metal2 s 49054 0 49110 800 6 wbs_dat_o[16]
port 582 nsew signal output
rlabel metal2 s 51446 0 51502 800 6 wbs_dat_o[17]
port 583 nsew signal output
rlabel metal2 s 53930 0 53986 800 6 wbs_dat_o[18]
port 584 nsew signal output
rlabel metal2 s 56322 0 56378 800 6 wbs_dat_o[19]
port 585 nsew signal output
rlabel metal2 s 10046 0 10102 800 6 wbs_dat_o[1]
port 586 nsew signal output
rlabel metal2 s 58806 0 58862 800 6 wbs_dat_o[20]
port 587 nsew signal output
rlabel metal2 s 61198 0 61254 800 6 wbs_dat_o[21]
port 588 nsew signal output
rlabel metal2 s 63590 0 63646 800 6 wbs_dat_o[22]
port 589 nsew signal output
rlabel metal2 s 66074 0 66130 800 6 wbs_dat_o[23]
port 590 nsew signal output
rlabel metal2 s 68466 0 68522 800 6 wbs_dat_o[24]
port 591 nsew signal output
rlabel metal2 s 70950 0 71006 800 6 wbs_dat_o[25]
port 592 nsew signal output
rlabel metal2 s 73342 0 73398 800 6 wbs_dat_o[26]
port 593 nsew signal output
rlabel metal2 s 75826 0 75882 800 6 wbs_dat_o[27]
port 594 nsew signal output
rlabel metal2 s 78218 0 78274 800 6 wbs_dat_o[28]
port 595 nsew signal output
rlabel metal2 s 80702 0 80758 800 6 wbs_dat_o[29]
port 596 nsew signal output
rlabel metal2 s 13358 0 13414 800 6 wbs_dat_o[2]
port 597 nsew signal output
rlabel metal2 s 83094 0 83150 800 6 wbs_dat_o[30]
port 598 nsew signal output
rlabel metal2 s 85578 0 85634 800 6 wbs_dat_o[31]
port 599 nsew signal output
rlabel metal2 s 16578 0 16634 800 6 wbs_dat_o[3]
port 600 nsew signal output
rlabel metal2 s 19798 0 19854 800 6 wbs_dat_o[4]
port 601 nsew signal output
rlabel metal2 s 22282 0 22338 800 6 wbs_dat_o[5]
port 602 nsew signal output
rlabel metal2 s 24674 0 24730 800 6 wbs_dat_o[6]
port 603 nsew signal output
rlabel metal2 s 27158 0 27214 800 6 wbs_dat_o[7]
port 604 nsew signal output
rlabel metal2 s 29550 0 29606 800 6 wbs_dat_o[8]
port 605 nsew signal output
rlabel metal2 s 31942 0 31998 800 6 wbs_dat_o[9]
port 606 nsew signal output
rlabel metal2 s 7654 0 7710 800 6 wbs_sel_i[0]
port 607 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 wbs_sel_i[1]
port 608 nsew signal input
rlabel metal2 s 14094 0 14150 800 6 wbs_sel_i[2]
port 609 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 wbs_sel_i[3]
port 610 nsew signal input
rlabel metal2 s 3606 0 3662 800 6 wbs_stb_i
port 611 nsew signal input
rlabel metal2 s 4434 0 4490 800 6 wbs_we_i
port 612 nsew signal input
rlabel metal4 s 372848 2128 373168 497808 6 VPWR
port 613 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 497808 6 VPWR
port 614 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 497808 6 VPWR
port 615 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 497808 6 VPWR
port 616 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 497808 6 VPWR
port 617 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 497808 6 VPWR
port 618 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 497808 6 VPWR
port 619 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 497808 6 VPWR
port 620 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 497808 6 VPWR
port 621 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 497808 6 VPWR
port 622 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 497808 6 VPWR
port 623 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 497808 6 VPWR
port 624 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 497808 6 VPWR
port 625 nsew power bidirectional
rlabel metal4 s 388208 2128 388528 497808 6 VGND
port 626 nsew ground bidirectional
rlabel metal4 s 357488 2128 357808 497808 6 VGND
port 627 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 497808 6 VGND
port 628 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 497808 6 VGND
port 629 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 497808 6 VGND
port 630 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 497808 6 VGND
port 631 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 497808 6 VGND
port 632 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 497808 6 VGND
port 633 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 497808 6 VGND
port 634 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 497808 6 VGND
port 635 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 497808 6 VGND
port 636 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 497808 6 VGND
port 637 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 497808 6 VGND
port 638 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 400000 500000
string LEFview TRUE
<< end >>
