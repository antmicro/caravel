VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2918.000 28.980 2924.000 30.180 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2918.000 2374.980 2924.000 2376.180 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2918.000 2609.580 2924.000 2610.780 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2918.000 2844.180 2924.000 2845.380 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2918.000 3078.780 2924.000 3079.980 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2918.000 3313.380 2924.000 3314.580 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3518.000 2879.650 3524.000 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3518.000 2555.350 3524.000 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3518.000 2231.050 3524.000 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3518.000 1906.290 3524.000 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3518.000 1581.990 3524.000 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2918.000 263.580 2924.000 264.780 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3518.000 1257.690 3524.000 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 932.370 3518.000 932.930 3524.000 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 608.070 3518.000 608.630 3524.000 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 283.770 3518.000 284.330 3524.000 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.000 3482.700 2.000 3483.900 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.000 3195.060 2.000 3196.260 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.000 2908.100 2.000 2909.300 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.000 2620.460 2.000 2621.660 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.000 2333.500 2.000 2334.700 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.000 2045.860 2.000 2047.060 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2918.000 498.180 2924.000 499.380 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.000 1758.900 2.000 1760.100 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2918.000 732.780 2924.000 733.980 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2918.000 967.380 2924.000 968.580 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2918.000 1201.980 2924.000 1203.180 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2918.000 1436.580 2924.000 1437.780 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2918.000 1671.180 2924.000 1672.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2918.000 1905.780 2924.000 1906.980 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2918.000 2140.380 2924.000 2141.580 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1140.485 89.505 1141.575 89.675 ;
      LAYER mcon ;
        RECT 1141.405 89.505 1141.575 89.675 ;
      LAYER met1 ;
        RECT 848.770 89.660 849.090 89.720 ;
        RECT 1140.425 89.660 1140.715 89.705 ;
        RECT 848.770 89.520 911.100 89.660 ;
        RECT 848.770 89.460 849.090 89.520 ;
        RECT 910.960 89.320 911.100 89.520 ;
        RECT 923.380 89.520 1140.715 89.660 ;
        RECT 923.380 89.320 923.520 89.520 ;
        RECT 1140.425 89.475 1140.715 89.520 ;
        RECT 1141.345 89.660 1141.635 89.705 ;
        RECT 2898.070 89.660 2898.390 89.720 ;
        RECT 1141.345 89.520 2898.390 89.660 ;
        RECT 1141.345 89.475 1141.635 89.520 ;
        RECT 2898.070 89.460 2898.390 89.520 ;
        RECT 910.960 89.180 923.520 89.320 ;
      LAYER via ;
        RECT 848.800 89.460 849.060 89.720 ;
        RECT 2898.100 89.460 2898.360 89.720 ;
      LAYER met2 ;
        RECT 854.230 2596.650 854.510 2600.000 ;
        RECT 848.860 2596.510 854.510 2596.650 ;
        RECT 848.860 89.750 849.000 2596.510 ;
        RECT 854.230 2596.000 854.510 2596.510 ;
        RECT 848.800 89.430 849.060 89.750 ;
        RECT 2898.100 89.430 2898.360 89.750 ;
        RECT 2898.160 88.245 2898.300 89.430 ;
        RECT 2898.090 87.875 2898.370 88.245 ;
      LAYER via2 ;
        RECT 2898.090 87.920 2898.370 88.200 ;
      LAYER met3 ;
        RECT 2898.065 88.210 2898.395 88.225 ;
        RECT 2918.000 88.210 2924.000 88.660 ;
        RECT 2898.065 87.910 2924.000 88.210 ;
        RECT 2898.065 87.895 2898.395 87.910 ;
        RECT 2918.000 87.460 2924.000 87.910 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1993.710 2430.220 1994.030 2430.280 ;
        RECT 2028.210 2430.220 2028.530 2430.280 ;
        RECT 1993.710 2430.080 2028.530 2430.220 ;
        RECT 1993.710 2430.020 1994.030 2430.080 ;
        RECT 2028.210 2430.020 2028.530 2430.080 ;
      LAYER via ;
        RECT 1993.740 2430.020 1994.000 2430.280 ;
        RECT 2028.240 2430.020 2028.500 2430.280 ;
      LAYER met2 ;
        RECT 1110.070 2614.755 1110.350 2615.125 ;
        RECT 1110.140 2600.050 1110.280 2614.755 ;
        RECT 1110.140 2600.000 1110.670 2600.050 ;
        RECT 1110.140 2599.910 1110.730 2600.000 ;
        RECT 1110.450 2596.000 1110.730 2599.910 ;
        RECT 2884.290 2434.555 2884.570 2434.925 ;
        RECT 2916.950 2434.555 2917.230 2434.925 ;
        RECT 1859.410 2431.835 1859.690 2432.205 ;
        RECT 1859.480 2429.485 1859.620 2431.835 ;
        RECT 1973.030 2431.155 1973.310 2431.525 ;
        RECT 1898.050 2430.050 1898.330 2430.165 ;
        RECT 1897.200 2429.910 1898.330 2430.050 ;
        RECT 1897.200 2429.485 1897.340 2429.910 ;
        RECT 1898.050 2429.795 1898.330 2429.910 ;
        RECT 1973.100 2429.485 1973.240 2431.155 ;
        RECT 2028.230 2430.475 2028.510 2430.845 ;
        RECT 2028.300 2430.310 2028.440 2430.475 ;
        RECT 1993.740 2430.165 1994.000 2430.310 ;
        RECT 1993.730 2429.795 1994.010 2430.165 ;
        RECT 2028.240 2429.990 2028.500 2430.310 ;
        RECT 2884.360 2429.485 2884.500 2434.555 ;
        RECT 2917.020 2434.245 2917.160 2434.555 ;
        RECT 2916.950 2433.875 2917.230 2434.245 ;
        RECT 1859.410 2429.115 1859.690 2429.485 ;
        RECT 1897.130 2429.115 1897.410 2429.485 ;
        RECT 1973.030 2429.115 1973.310 2429.485 ;
        RECT 2884.290 2429.115 2884.570 2429.485 ;
      LAYER via2 ;
        RECT 1110.070 2614.800 1110.350 2615.080 ;
        RECT 2884.290 2434.600 2884.570 2434.880 ;
        RECT 2916.950 2434.600 2917.230 2434.880 ;
        RECT 1859.410 2431.880 1859.690 2432.160 ;
        RECT 1973.030 2431.200 1973.310 2431.480 ;
        RECT 1898.050 2429.840 1898.330 2430.120 ;
        RECT 2028.230 2430.520 2028.510 2430.800 ;
        RECT 1993.730 2429.840 1994.010 2430.120 ;
        RECT 2916.950 2433.920 2917.230 2434.200 ;
        RECT 1859.410 2429.160 1859.690 2429.440 ;
        RECT 1897.130 2429.160 1897.410 2429.440 ;
        RECT 1973.030 2429.160 1973.310 2429.440 ;
        RECT 2884.290 2429.160 2884.570 2429.440 ;
      LAYER met3 ;
        RECT 1110.045 2615.090 1110.375 2615.105 ;
        RECT 1798.870 2615.090 1799.250 2615.100 ;
        RECT 1110.045 2614.790 1799.250 2615.090 ;
        RECT 1110.045 2614.775 1110.375 2614.790 ;
        RECT 1798.870 2614.780 1799.250 2614.790 ;
        RECT 2884.265 2434.890 2884.595 2434.905 ;
        RECT 2916.925 2434.890 2917.255 2434.905 ;
        RECT 2884.265 2434.590 2917.255 2434.890 ;
        RECT 2884.265 2434.575 2884.595 2434.590 ;
        RECT 2916.925 2434.575 2917.255 2434.590 ;
        RECT 2916.925 2434.210 2917.255 2434.225 ;
        RECT 2918.000 2434.210 2924.000 2434.660 ;
        RECT 2916.925 2433.910 2924.000 2434.210 ;
        RECT 2916.925 2433.895 2917.255 2433.910 ;
        RECT 2918.000 2433.460 2924.000 2433.910 ;
        RECT 1835.670 2432.170 1836.050 2432.180 ;
        RECT 1859.385 2432.170 1859.715 2432.185 ;
        RECT 1835.670 2431.870 1859.715 2432.170 ;
        RECT 1835.670 2431.860 1836.050 2431.870 ;
        RECT 1859.385 2431.855 1859.715 2431.870 ;
        RECT 1924.910 2431.490 1925.290 2431.500 ;
        RECT 1973.005 2431.490 1973.335 2431.505 ;
        RECT 1924.910 2431.190 1973.335 2431.490 ;
        RECT 1924.910 2431.180 1925.290 2431.190 ;
        RECT 1973.005 2431.175 1973.335 2431.190 ;
        RECT 1835.670 2430.810 1836.050 2430.820 ;
        RECT 1800.750 2430.510 1836.050 2430.810 ;
        RECT 1798.870 2429.450 1799.250 2429.460 ;
        RECT 1800.750 2429.450 1801.050 2430.510 ;
        RECT 1835.670 2430.500 1836.050 2430.510 ;
        RECT 2028.205 2430.810 2028.535 2430.825 ;
        RECT 2028.205 2430.510 2063.250 2430.810 ;
        RECT 2028.205 2430.495 2028.535 2430.510 ;
        RECT 1898.025 2430.130 1898.355 2430.145 ;
        RECT 1924.910 2430.130 1925.290 2430.140 ;
        RECT 1993.705 2430.130 1994.035 2430.145 ;
        RECT 1898.025 2429.830 1925.290 2430.130 ;
        RECT 1898.025 2429.815 1898.355 2429.830 ;
        RECT 1924.910 2429.820 1925.290 2429.830 ;
        RECT 1980.150 2429.830 1994.035 2430.130 ;
        RECT 2062.950 2430.130 2063.250 2430.510 ;
        RECT 2111.710 2430.510 2159.850 2430.810 ;
        RECT 2062.950 2429.830 2111.090 2430.130 ;
        RECT 1798.870 2429.150 1801.050 2429.450 ;
        RECT 1859.385 2429.450 1859.715 2429.465 ;
        RECT 1897.105 2429.450 1897.435 2429.465 ;
        RECT 1859.385 2429.150 1897.435 2429.450 ;
        RECT 1798.870 2429.140 1799.250 2429.150 ;
        RECT 1859.385 2429.135 1859.715 2429.150 ;
        RECT 1897.105 2429.135 1897.435 2429.150 ;
        RECT 1973.005 2429.450 1973.335 2429.465 ;
        RECT 1980.150 2429.450 1980.450 2429.830 ;
        RECT 1993.705 2429.815 1994.035 2429.830 ;
        RECT 1973.005 2429.150 1980.450 2429.450 ;
        RECT 2110.790 2429.450 2111.090 2429.830 ;
        RECT 2111.710 2429.450 2112.010 2430.510 ;
        RECT 2159.550 2430.130 2159.850 2430.510 ;
        RECT 2208.310 2430.510 2256.450 2430.810 ;
        RECT 2159.550 2429.830 2207.690 2430.130 ;
        RECT 2110.790 2429.150 2112.010 2429.450 ;
        RECT 2207.390 2429.450 2207.690 2429.830 ;
        RECT 2208.310 2429.450 2208.610 2430.510 ;
        RECT 2256.150 2430.130 2256.450 2430.510 ;
        RECT 2304.910 2430.510 2353.050 2430.810 ;
        RECT 2256.150 2429.830 2304.290 2430.130 ;
        RECT 2207.390 2429.150 2208.610 2429.450 ;
        RECT 2303.990 2429.450 2304.290 2429.830 ;
        RECT 2304.910 2429.450 2305.210 2430.510 ;
        RECT 2352.750 2430.130 2353.050 2430.510 ;
        RECT 2401.510 2430.510 2449.650 2430.810 ;
        RECT 2352.750 2429.830 2400.890 2430.130 ;
        RECT 2303.990 2429.150 2305.210 2429.450 ;
        RECT 2400.590 2429.450 2400.890 2429.830 ;
        RECT 2401.510 2429.450 2401.810 2430.510 ;
        RECT 2449.350 2430.130 2449.650 2430.510 ;
        RECT 2498.110 2430.510 2546.250 2430.810 ;
        RECT 2449.350 2429.830 2497.490 2430.130 ;
        RECT 2400.590 2429.150 2401.810 2429.450 ;
        RECT 2497.190 2429.450 2497.490 2429.830 ;
        RECT 2498.110 2429.450 2498.410 2430.510 ;
        RECT 2545.950 2430.130 2546.250 2430.510 ;
        RECT 2594.710 2430.510 2642.850 2430.810 ;
        RECT 2545.950 2429.830 2594.090 2430.130 ;
        RECT 2497.190 2429.150 2498.410 2429.450 ;
        RECT 2593.790 2429.450 2594.090 2429.830 ;
        RECT 2594.710 2429.450 2595.010 2430.510 ;
        RECT 2642.550 2430.130 2642.850 2430.510 ;
        RECT 2691.310 2430.510 2739.450 2430.810 ;
        RECT 2642.550 2429.830 2690.690 2430.130 ;
        RECT 2593.790 2429.150 2595.010 2429.450 ;
        RECT 2690.390 2429.450 2690.690 2429.830 ;
        RECT 2691.310 2429.450 2691.610 2430.510 ;
        RECT 2739.150 2430.130 2739.450 2430.510 ;
        RECT 2787.910 2430.510 2836.050 2430.810 ;
        RECT 2739.150 2429.830 2787.290 2430.130 ;
        RECT 2690.390 2429.150 2691.610 2429.450 ;
        RECT 2786.990 2429.450 2787.290 2429.830 ;
        RECT 2787.910 2429.450 2788.210 2430.510 ;
        RECT 2835.750 2430.130 2836.050 2430.510 ;
        RECT 2835.750 2429.830 2883.890 2430.130 ;
        RECT 2786.990 2429.150 2788.210 2429.450 ;
        RECT 2883.590 2429.450 2883.890 2429.830 ;
        RECT 2884.265 2429.450 2884.595 2429.465 ;
        RECT 2883.590 2429.150 2884.595 2429.450 ;
        RECT 1973.005 2429.135 1973.335 2429.150 ;
        RECT 2884.265 2429.135 2884.595 2429.150 ;
      LAYER via3 ;
        RECT 1798.900 2614.780 1799.220 2615.100 ;
        RECT 1835.700 2431.860 1836.020 2432.180 ;
        RECT 1924.940 2431.180 1925.260 2431.500 ;
        RECT 1798.900 2429.140 1799.220 2429.460 ;
        RECT 1835.700 2430.500 1836.020 2430.820 ;
        RECT 1924.940 2429.820 1925.260 2430.140 ;
      LAYER met4 ;
        RECT 1798.895 2614.775 1799.225 2615.105 ;
        RECT 1798.910 2429.465 1799.210 2614.775 ;
        RECT 1835.695 2431.855 1836.025 2432.185 ;
        RECT 1835.710 2430.825 1836.010 2431.855 ;
        RECT 1924.935 2431.175 1925.265 2431.505 ;
        RECT 1835.695 2430.495 1836.025 2430.825 ;
        RECT 1924.950 2430.145 1925.250 2431.175 ;
        RECT 1924.935 2429.815 1925.265 2430.145 ;
        RECT 1798.895 2429.135 1799.225 2429.465 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1138.110 2663.800 1138.430 2663.860 ;
        RECT 2901.290 2663.800 2901.610 2663.860 ;
        RECT 1138.110 2663.660 2901.610 2663.800 ;
        RECT 1138.110 2663.600 1138.430 2663.660 ;
        RECT 2901.290 2663.600 2901.610 2663.660 ;
      LAYER via ;
        RECT 1138.140 2663.600 1138.400 2663.860 ;
        RECT 2901.320 2663.600 2901.580 2663.860 ;
      LAYER met2 ;
        RECT 2901.310 2669.155 2901.590 2669.525 ;
        RECT 2901.380 2663.890 2901.520 2669.155 ;
        RECT 1138.140 2663.570 1138.400 2663.890 ;
        RECT 2901.320 2663.570 2901.580 2663.890 ;
        RECT 1136.210 2599.370 1136.490 2600.000 ;
        RECT 1138.200 2599.370 1138.340 2663.570 ;
        RECT 1136.210 2599.230 1138.340 2599.370 ;
        RECT 1136.210 2596.000 1136.490 2599.230 ;
      LAYER via2 ;
        RECT 2901.310 2669.200 2901.590 2669.480 ;
      LAYER met3 ;
        RECT 2901.285 2669.490 2901.615 2669.505 ;
        RECT 2918.000 2669.490 2924.000 2669.940 ;
        RECT 2901.285 2669.190 2924.000 2669.490 ;
        RECT 2901.285 2669.175 2901.615 2669.190 ;
        RECT 2918.000 2668.740 2924.000 2669.190 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1165.710 2898.400 1166.030 2898.460 ;
        RECT 2901.290 2898.400 2901.610 2898.460 ;
        RECT 1165.710 2898.260 2901.610 2898.400 ;
        RECT 1165.710 2898.200 1166.030 2898.260 ;
        RECT 2901.290 2898.200 2901.610 2898.260 ;
        RECT 1159.270 2632.520 1159.590 2632.580 ;
        RECT 1165.710 2632.520 1166.030 2632.580 ;
        RECT 1159.270 2632.380 1166.030 2632.520 ;
        RECT 1159.270 2632.320 1159.590 2632.380 ;
        RECT 1165.710 2632.320 1166.030 2632.380 ;
      LAYER via ;
        RECT 1165.740 2898.200 1166.000 2898.460 ;
        RECT 2901.320 2898.200 2901.580 2898.460 ;
        RECT 1159.300 2632.320 1159.560 2632.580 ;
        RECT 1165.740 2632.320 1166.000 2632.580 ;
      LAYER met2 ;
        RECT 2901.310 2903.755 2901.590 2904.125 ;
        RECT 2901.380 2898.490 2901.520 2903.755 ;
        RECT 1165.740 2898.170 1166.000 2898.490 ;
        RECT 2901.320 2898.170 2901.580 2898.490 ;
        RECT 1165.800 2632.610 1165.940 2898.170 ;
        RECT 1159.300 2632.290 1159.560 2632.610 ;
        RECT 1165.740 2632.290 1166.000 2632.610 ;
        RECT 1159.360 2599.370 1159.500 2632.290 ;
        RECT 1161.510 2599.370 1161.790 2600.000 ;
        RECT 1159.360 2599.230 1161.790 2599.370 ;
        RECT 1161.510 2596.000 1161.790 2599.230 ;
      LAYER via2 ;
        RECT 2901.310 2903.800 2901.590 2904.080 ;
      LAYER met3 ;
        RECT 2901.285 2904.090 2901.615 2904.105 ;
        RECT 2918.000 2904.090 2924.000 2904.540 ;
        RECT 2901.285 2903.790 2924.000 2904.090 ;
        RECT 2901.285 2903.775 2901.615 2903.790 ;
        RECT 2918.000 2903.340 2924.000 2903.790 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1193.310 3133.000 1193.630 3133.060 ;
        RECT 2901.290 3133.000 2901.610 3133.060 ;
        RECT 1193.310 3132.860 2901.610 3133.000 ;
        RECT 1193.310 3132.800 1193.630 3132.860 ;
        RECT 2901.290 3132.800 2901.610 3132.860 ;
        RECT 1186.870 2632.520 1187.190 2632.580 ;
        RECT 1193.310 2632.520 1193.630 2632.580 ;
        RECT 1186.870 2632.380 1193.630 2632.520 ;
        RECT 1186.870 2632.320 1187.190 2632.380 ;
        RECT 1193.310 2632.320 1193.630 2632.380 ;
      LAYER via ;
        RECT 1193.340 3132.800 1193.600 3133.060 ;
        RECT 2901.320 3132.800 2901.580 3133.060 ;
        RECT 1186.900 2632.320 1187.160 2632.580 ;
        RECT 1193.340 2632.320 1193.600 2632.580 ;
      LAYER met2 ;
        RECT 2901.310 3138.355 2901.590 3138.725 ;
        RECT 2901.380 3133.090 2901.520 3138.355 ;
        RECT 1193.340 3132.770 1193.600 3133.090 ;
        RECT 2901.320 3132.770 2901.580 3133.090 ;
        RECT 1193.400 2632.610 1193.540 3132.770 ;
        RECT 1186.900 2632.290 1187.160 2632.610 ;
        RECT 1193.340 2632.290 1193.600 2632.610 ;
        RECT 1186.960 2600.050 1187.100 2632.290 ;
        RECT 1186.960 2600.000 1187.490 2600.050 ;
        RECT 1186.960 2599.910 1187.550 2600.000 ;
        RECT 1187.270 2596.000 1187.550 2599.910 ;
      LAYER via2 ;
        RECT 2901.310 3138.400 2901.590 3138.680 ;
      LAYER met3 ;
        RECT 2901.285 3138.690 2901.615 3138.705 ;
        RECT 2918.000 3138.690 2924.000 3139.140 ;
        RECT 2901.285 3138.390 2924.000 3138.690 ;
        RECT 2901.285 3138.375 2901.615 3138.390 ;
        RECT 2918.000 3137.940 2924.000 3138.390 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1214.010 3367.600 1214.330 3367.660 ;
        RECT 2901.290 3367.600 2901.610 3367.660 ;
        RECT 1214.010 3367.460 2901.610 3367.600 ;
        RECT 1214.010 3367.400 1214.330 3367.460 ;
        RECT 2901.290 3367.400 2901.610 3367.460 ;
      LAYER via ;
        RECT 1214.040 3367.400 1214.300 3367.660 ;
        RECT 2901.320 3367.400 2901.580 3367.660 ;
      LAYER met2 ;
        RECT 2901.310 3372.955 2901.590 3373.325 ;
        RECT 2901.380 3367.690 2901.520 3372.955 ;
        RECT 1214.040 3367.370 1214.300 3367.690 ;
        RECT 2901.320 3367.370 2901.580 3367.690 ;
        RECT 1213.030 2599.370 1213.310 2600.000 ;
        RECT 1214.100 2599.370 1214.240 3367.370 ;
        RECT 1213.030 2599.230 1214.240 2599.370 ;
        RECT 1213.030 2596.000 1213.310 2599.230 ;
      LAYER via2 ;
        RECT 2901.310 3373.000 2901.590 3373.280 ;
      LAYER met3 ;
        RECT 2901.285 3373.290 2901.615 3373.305 ;
        RECT 2918.000 3373.290 2924.000 3373.740 ;
        RECT 2901.285 3372.990 2924.000 3373.290 ;
        RECT 2901.285 3372.975 2901.615 3372.990 ;
        RECT 2918.000 3372.540 2924.000 3372.990 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2796.485 3332.765 2796.655 3422.355 ;
        RECT 2795.565 3008.405 2795.735 3042.915 ;
        RECT 2796.485 2946.525 2796.655 2994.635 ;
        RECT 2795.105 2753.065 2795.275 2801.175 ;
      LAYER mcon ;
        RECT 2796.485 3422.185 2796.655 3422.355 ;
        RECT 2795.565 3042.745 2795.735 3042.915 ;
        RECT 2796.485 2994.465 2796.655 2994.635 ;
        RECT 2795.105 2801.005 2795.275 2801.175 ;
      LAYER met1 ;
        RECT 2795.490 3443.080 2795.810 3443.140 ;
        RECT 2798.250 3443.080 2798.570 3443.140 ;
        RECT 2795.490 3442.940 2798.570 3443.080 ;
        RECT 2795.490 3442.880 2795.810 3442.940 ;
        RECT 2798.250 3442.880 2798.570 3442.940 ;
        RECT 2795.030 3422.340 2795.350 3422.400 ;
        RECT 2796.425 3422.340 2796.715 3422.385 ;
        RECT 2795.030 3422.200 2796.715 3422.340 ;
        RECT 2795.030 3422.140 2795.350 3422.200 ;
        RECT 2796.425 3422.155 2796.715 3422.200 ;
        RECT 2796.425 3332.920 2796.715 3332.965 ;
        RECT 2796.870 3332.920 2797.190 3332.980 ;
        RECT 2796.425 3332.780 2797.190 3332.920 ;
        RECT 2796.425 3332.735 2796.715 3332.780 ;
        RECT 2796.870 3332.720 2797.190 3332.780 ;
        RECT 2795.490 3236.360 2795.810 3236.420 ;
        RECT 2795.950 3236.360 2796.270 3236.420 ;
        RECT 2795.490 3236.220 2796.270 3236.360 ;
        RECT 2795.490 3236.160 2795.810 3236.220 ;
        RECT 2795.950 3236.160 2796.270 3236.220 ;
        RECT 2795.490 3202.020 2795.810 3202.080 ;
        RECT 2795.950 3202.020 2796.270 3202.080 ;
        RECT 2795.490 3201.880 2796.270 3202.020 ;
        RECT 2795.490 3201.820 2795.810 3201.880 ;
        RECT 2795.950 3201.820 2796.270 3201.880 ;
        RECT 2795.030 3153.400 2795.350 3153.460 ;
        RECT 2795.950 3153.400 2796.270 3153.460 ;
        RECT 2795.030 3153.260 2796.270 3153.400 ;
        RECT 2795.030 3153.200 2795.350 3153.260 ;
        RECT 2795.950 3153.200 2796.270 3153.260 ;
        RECT 2795.030 3056.840 2795.350 3056.900 ;
        RECT 2795.950 3056.840 2796.270 3056.900 ;
        RECT 2795.030 3056.700 2796.270 3056.840 ;
        RECT 2795.030 3056.640 2795.350 3056.700 ;
        RECT 2795.950 3056.640 2796.270 3056.700 ;
        RECT 2795.490 3042.900 2795.810 3042.960 ;
        RECT 2795.295 3042.760 2795.810 3042.900 ;
        RECT 2795.490 3042.700 2795.810 3042.760 ;
        RECT 2795.505 3008.560 2795.795 3008.605 ;
        RECT 2796.410 3008.560 2796.730 3008.620 ;
        RECT 2795.505 3008.420 2796.730 3008.560 ;
        RECT 2795.505 3008.375 2795.795 3008.420 ;
        RECT 2796.410 3008.360 2796.730 3008.420 ;
        RECT 2796.410 2994.620 2796.730 2994.680 ;
        RECT 2796.215 2994.480 2796.730 2994.620 ;
        RECT 2796.410 2994.420 2796.730 2994.480 ;
        RECT 2796.425 2946.680 2796.715 2946.725 ;
        RECT 2796.870 2946.680 2797.190 2946.740 ;
        RECT 2796.425 2946.540 2797.190 2946.680 ;
        RECT 2796.425 2946.495 2796.715 2946.540 ;
        RECT 2796.870 2946.480 2797.190 2946.540 ;
        RECT 2796.870 2912.340 2797.190 2912.400 ;
        RECT 2796.500 2912.200 2797.190 2912.340 ;
        RECT 2796.500 2911.720 2796.640 2912.200 ;
        RECT 2796.870 2912.140 2797.190 2912.200 ;
        RECT 2796.410 2911.460 2796.730 2911.720 ;
        RECT 2795.030 2815.580 2795.350 2815.840 ;
        RECT 2795.120 2815.160 2795.260 2815.580 ;
        RECT 2795.030 2814.900 2795.350 2815.160 ;
        RECT 2795.030 2801.160 2795.350 2801.220 ;
        RECT 2794.835 2801.020 2795.350 2801.160 ;
        RECT 2795.030 2800.960 2795.350 2801.020 ;
        RECT 2795.045 2753.220 2795.335 2753.265 ;
        RECT 2795.950 2753.220 2796.270 2753.280 ;
        RECT 2795.045 2753.080 2796.270 2753.220 ;
        RECT 2795.045 2753.035 2795.335 2753.080 ;
        RECT 2795.950 2753.020 2796.270 2753.080 ;
        RECT 2795.030 2718.200 2795.350 2718.260 ;
        RECT 2795.950 2718.200 2796.270 2718.260 ;
        RECT 2795.030 2718.060 2796.270 2718.200 ;
        RECT 2795.030 2718.000 2795.350 2718.060 ;
        RECT 2795.950 2718.000 2796.270 2718.060 ;
        RECT 1240.690 2618.580 1241.010 2618.640 ;
        RECT 2795.950 2618.580 2796.270 2618.640 ;
        RECT 1240.690 2618.440 2796.270 2618.580 ;
        RECT 1240.690 2618.380 1241.010 2618.440 ;
        RECT 2795.950 2618.380 2796.270 2618.440 ;
      LAYER via ;
        RECT 2795.520 3442.880 2795.780 3443.140 ;
        RECT 2798.280 3442.880 2798.540 3443.140 ;
        RECT 2795.060 3422.140 2795.320 3422.400 ;
        RECT 2796.900 3332.720 2797.160 3332.980 ;
        RECT 2795.520 3236.160 2795.780 3236.420 ;
        RECT 2795.980 3236.160 2796.240 3236.420 ;
        RECT 2795.520 3201.820 2795.780 3202.080 ;
        RECT 2795.980 3201.820 2796.240 3202.080 ;
        RECT 2795.060 3153.200 2795.320 3153.460 ;
        RECT 2795.980 3153.200 2796.240 3153.460 ;
        RECT 2795.060 3056.640 2795.320 3056.900 ;
        RECT 2795.980 3056.640 2796.240 3056.900 ;
        RECT 2795.520 3042.700 2795.780 3042.960 ;
        RECT 2796.440 3008.360 2796.700 3008.620 ;
        RECT 2796.440 2994.420 2796.700 2994.680 ;
        RECT 2796.900 2946.480 2797.160 2946.740 ;
        RECT 2796.900 2912.140 2797.160 2912.400 ;
        RECT 2796.440 2911.460 2796.700 2911.720 ;
        RECT 2795.060 2815.580 2795.320 2815.840 ;
        RECT 2795.060 2814.900 2795.320 2815.160 ;
        RECT 2795.060 2800.960 2795.320 2801.220 ;
        RECT 2795.980 2753.020 2796.240 2753.280 ;
        RECT 2795.060 2718.000 2795.320 2718.260 ;
        RECT 2795.980 2718.000 2796.240 2718.260 ;
        RECT 1240.720 2618.380 1240.980 2618.640 ;
        RECT 2795.980 2618.380 2796.240 2618.640 ;
      LAYER met2 ;
        RECT 2798.130 3518.000 2798.690 3524.000 ;
        RECT 2798.340 3443.170 2798.480 3518.000 ;
        RECT 2795.520 3442.850 2795.780 3443.170 ;
        RECT 2798.280 3442.850 2798.540 3443.170 ;
        RECT 2795.580 3429.650 2795.720 3442.850 ;
        RECT 2795.120 3429.510 2795.720 3429.650 ;
        RECT 2795.120 3422.430 2795.260 3429.510 ;
        RECT 2795.060 3422.110 2795.320 3422.430 ;
        RECT 2796.900 3332.690 2797.160 3333.010 ;
        RECT 2796.960 3298.410 2797.100 3332.690 ;
        RECT 2796.040 3298.270 2797.100 3298.410 ;
        RECT 2796.040 3236.450 2796.180 3298.270 ;
        RECT 2795.520 3236.130 2795.780 3236.450 ;
        RECT 2795.980 3236.130 2796.240 3236.450 ;
        RECT 2795.580 3202.110 2795.720 3236.130 ;
        RECT 2795.520 3201.790 2795.780 3202.110 ;
        RECT 2795.980 3201.790 2796.240 3202.110 ;
        RECT 2796.040 3153.490 2796.180 3201.790 ;
        RECT 2795.060 3153.170 2795.320 3153.490 ;
        RECT 2795.980 3153.170 2796.240 3153.490 ;
        RECT 2795.120 3152.890 2795.260 3153.170 ;
        RECT 2795.120 3152.750 2795.720 3152.890 ;
        RECT 2795.580 3105.290 2795.720 3152.750 ;
        RECT 2795.580 3105.150 2796.180 3105.290 ;
        RECT 2796.040 3056.930 2796.180 3105.150 ;
        RECT 2795.060 3056.610 2795.320 3056.930 ;
        RECT 2795.980 3056.610 2796.240 3056.930 ;
        RECT 2795.120 3056.330 2795.260 3056.610 ;
        RECT 2795.120 3056.190 2795.720 3056.330 ;
        RECT 2795.580 3042.990 2795.720 3056.190 ;
        RECT 2795.520 3042.670 2795.780 3042.990 ;
        RECT 2796.440 3008.330 2796.700 3008.650 ;
        RECT 2796.500 2994.710 2796.640 3008.330 ;
        RECT 2796.440 2994.390 2796.700 2994.710 ;
        RECT 2796.900 2946.450 2797.160 2946.770 ;
        RECT 2796.960 2912.430 2797.100 2946.450 ;
        RECT 2796.900 2912.110 2797.160 2912.430 ;
        RECT 2796.440 2911.430 2796.700 2911.750 ;
        RECT 2796.500 2863.210 2796.640 2911.430 ;
        RECT 2795.580 2863.070 2796.640 2863.210 ;
        RECT 2795.580 2849.610 2795.720 2863.070 ;
        RECT 2795.120 2849.470 2795.720 2849.610 ;
        RECT 2795.120 2815.870 2795.260 2849.470 ;
        RECT 2795.060 2815.550 2795.320 2815.870 ;
        RECT 2795.060 2814.870 2795.320 2815.190 ;
        RECT 2795.120 2801.250 2795.260 2814.870 ;
        RECT 2795.060 2800.930 2795.320 2801.250 ;
        RECT 2795.980 2752.990 2796.240 2753.310 ;
        RECT 2796.040 2718.290 2796.180 2752.990 ;
        RECT 2795.060 2717.970 2795.320 2718.290 ;
        RECT 2795.980 2717.970 2796.240 2718.290 ;
        RECT 2795.120 2670.090 2795.260 2717.970 ;
        RECT 2795.120 2669.950 2795.720 2670.090 ;
        RECT 2795.580 2622.490 2795.720 2669.950 ;
        RECT 2795.580 2622.350 2796.180 2622.490 ;
        RECT 2796.040 2618.670 2796.180 2622.350 ;
        RECT 1240.720 2618.350 1240.980 2618.670 ;
        RECT 2795.980 2618.350 2796.240 2618.670 ;
        RECT 1238.790 2599.370 1239.070 2600.000 ;
        RECT 1240.780 2599.370 1240.920 2618.350 ;
        RECT 1238.790 2599.230 1240.920 2599.370 ;
        RECT 1238.790 2596.000 1239.070 2599.230 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2470.345 3332.765 2470.515 3380.875 ;
        RECT 2470.805 2815.285 2470.975 2849.455 ;
      LAYER mcon ;
        RECT 2470.345 3380.705 2470.515 3380.875 ;
        RECT 2470.805 2849.285 2470.975 2849.455 ;
      LAYER met1 ;
        RECT 2470.270 3380.860 2470.590 3380.920 ;
        RECT 2470.075 3380.720 2470.590 3380.860 ;
        RECT 2470.270 3380.660 2470.590 3380.720 ;
        RECT 2470.285 3332.920 2470.575 3332.965 ;
        RECT 2470.730 3332.920 2471.050 3332.980 ;
        RECT 2470.285 3332.780 2471.050 3332.920 ;
        RECT 2470.285 3332.735 2470.575 3332.780 ;
        RECT 2470.730 3332.720 2471.050 3332.780 ;
        RECT 2470.270 3270.700 2470.590 3270.760 ;
        RECT 2471.190 3270.700 2471.510 3270.760 ;
        RECT 2470.270 3270.560 2471.510 3270.700 ;
        RECT 2470.270 3270.500 2470.590 3270.560 ;
        RECT 2471.190 3270.500 2471.510 3270.560 ;
        RECT 2470.270 3174.140 2470.590 3174.200 ;
        RECT 2471.190 3174.140 2471.510 3174.200 ;
        RECT 2470.270 3174.000 2471.510 3174.140 ;
        RECT 2470.270 3173.940 2470.590 3174.000 ;
        RECT 2471.190 3173.940 2471.510 3174.000 ;
        RECT 2470.270 3077.580 2470.590 3077.640 ;
        RECT 2471.190 3077.580 2471.510 3077.640 ;
        RECT 2470.270 3077.440 2471.510 3077.580 ;
        RECT 2470.270 3077.380 2470.590 3077.440 ;
        RECT 2471.190 3077.380 2471.510 3077.440 ;
        RECT 2470.270 2981.020 2470.590 2981.080 ;
        RECT 2471.190 2981.020 2471.510 2981.080 ;
        RECT 2470.270 2980.880 2471.510 2981.020 ;
        RECT 2470.270 2980.820 2470.590 2980.880 ;
        RECT 2471.190 2980.820 2471.510 2980.880 ;
        RECT 2469.350 2946.340 2469.670 2946.400 ;
        RECT 2470.730 2946.340 2471.050 2946.400 ;
        RECT 2469.350 2946.200 2471.050 2946.340 ;
        RECT 2469.350 2946.140 2469.670 2946.200 ;
        RECT 2470.730 2946.140 2471.050 2946.200 ;
        RECT 2470.730 2849.440 2471.050 2849.500 ;
        RECT 2470.535 2849.300 2471.050 2849.440 ;
        RECT 2470.730 2849.240 2471.050 2849.300 ;
        RECT 2470.745 2815.440 2471.035 2815.485 ;
        RECT 2471.650 2815.440 2471.970 2815.500 ;
        RECT 2470.745 2815.300 2471.970 2815.440 ;
        RECT 2470.745 2815.255 2471.035 2815.300 ;
        RECT 2471.650 2815.240 2471.970 2815.300 ;
        RECT 2470.730 2753.220 2471.050 2753.280 ;
        RECT 2472.110 2753.220 2472.430 2753.280 ;
        RECT 2470.730 2753.080 2472.430 2753.220 ;
        RECT 2470.730 2753.020 2471.050 2753.080 ;
        RECT 2472.110 2753.020 2472.430 2753.080 ;
        RECT 2472.110 2719.220 2472.430 2719.280 ;
        RECT 2471.740 2719.080 2472.430 2719.220 ;
        RECT 2471.740 2718.600 2471.880 2719.080 ;
        RECT 2472.110 2719.020 2472.430 2719.080 ;
        RECT 2471.650 2718.340 2471.970 2718.600 ;
        RECT 2470.730 2656.660 2471.050 2656.720 ;
        RECT 2472.110 2656.660 2472.430 2656.720 ;
        RECT 2470.730 2656.520 2472.430 2656.660 ;
        RECT 2470.730 2656.460 2471.050 2656.520 ;
        RECT 2472.110 2656.460 2472.430 2656.520 ;
        RECT 1265.530 2618.920 1265.850 2618.980 ;
        RECT 2472.110 2618.920 2472.430 2618.980 ;
        RECT 1265.530 2618.780 2472.430 2618.920 ;
        RECT 1265.530 2618.720 1265.850 2618.780 ;
        RECT 2472.110 2618.720 2472.430 2618.780 ;
      LAYER via ;
        RECT 2470.300 3380.660 2470.560 3380.920 ;
        RECT 2470.760 3332.720 2471.020 3332.980 ;
        RECT 2470.300 3270.500 2470.560 3270.760 ;
        RECT 2471.220 3270.500 2471.480 3270.760 ;
        RECT 2470.300 3173.940 2470.560 3174.200 ;
        RECT 2471.220 3173.940 2471.480 3174.200 ;
        RECT 2470.300 3077.380 2470.560 3077.640 ;
        RECT 2471.220 3077.380 2471.480 3077.640 ;
        RECT 2470.300 2980.820 2470.560 2981.080 ;
        RECT 2471.220 2980.820 2471.480 2981.080 ;
        RECT 2469.380 2946.140 2469.640 2946.400 ;
        RECT 2470.760 2946.140 2471.020 2946.400 ;
        RECT 2470.760 2849.240 2471.020 2849.500 ;
        RECT 2471.680 2815.240 2471.940 2815.500 ;
        RECT 2470.760 2753.020 2471.020 2753.280 ;
        RECT 2472.140 2753.020 2472.400 2753.280 ;
        RECT 2472.140 2719.020 2472.400 2719.280 ;
        RECT 2471.680 2718.340 2471.940 2718.600 ;
        RECT 2470.760 2656.460 2471.020 2656.720 ;
        RECT 2472.140 2656.460 2472.400 2656.720 ;
        RECT 1265.560 2618.720 1265.820 2618.980 ;
        RECT 2472.140 2618.720 2472.400 2618.980 ;
      LAYER met2 ;
        RECT 2473.830 3518.050 2474.390 3524.000 ;
        RECT 2473.830 3518.000 2474.640 3518.050 ;
        RECT 2474.040 3517.910 2474.640 3518.000 ;
        RECT 2474.500 3430.445 2474.640 3517.910 ;
        RECT 2474.430 3430.075 2474.710 3430.445 ;
        RECT 2471.210 3429.395 2471.490 3429.765 ;
        RECT 2471.280 3394.970 2471.420 3429.395 ;
        RECT 2470.360 3394.830 2471.420 3394.970 ;
        RECT 2470.360 3380.950 2470.500 3394.830 ;
        RECT 2470.300 3380.630 2470.560 3380.950 ;
        RECT 2470.760 3332.690 2471.020 3333.010 ;
        RECT 2470.820 3298.410 2470.960 3332.690 ;
        RECT 2470.820 3298.270 2471.420 3298.410 ;
        RECT 2471.280 3270.790 2471.420 3298.270 ;
        RECT 2470.300 3270.470 2470.560 3270.790 ;
        RECT 2471.220 3270.470 2471.480 3270.790 ;
        RECT 2470.360 3222.250 2470.500 3270.470 ;
        RECT 2470.360 3222.110 2471.420 3222.250 ;
        RECT 2471.280 3174.230 2471.420 3222.110 ;
        RECT 2470.300 3173.910 2470.560 3174.230 ;
        RECT 2471.220 3173.910 2471.480 3174.230 ;
        RECT 2470.360 3125.690 2470.500 3173.910 ;
        RECT 2470.360 3125.550 2471.420 3125.690 ;
        RECT 2471.280 3077.670 2471.420 3125.550 ;
        RECT 2470.300 3077.350 2470.560 3077.670 ;
        RECT 2471.220 3077.350 2471.480 3077.670 ;
        RECT 2470.360 3029.130 2470.500 3077.350 ;
        RECT 2470.360 3028.990 2471.420 3029.130 ;
        RECT 2471.280 2981.110 2471.420 3028.990 ;
        RECT 2470.300 2980.850 2470.560 2981.110 ;
        RECT 2470.300 2980.790 2470.960 2980.850 ;
        RECT 2471.220 2980.790 2471.480 2981.110 ;
        RECT 2470.360 2980.710 2470.960 2980.790 ;
        RECT 2470.820 2980.170 2470.960 2980.710 ;
        RECT 2470.820 2980.030 2471.420 2980.170 ;
        RECT 2471.280 2959.770 2471.420 2980.030 ;
        RECT 2470.820 2959.630 2471.420 2959.770 ;
        RECT 2470.820 2946.430 2470.960 2959.630 ;
        RECT 2469.380 2946.110 2469.640 2946.430 ;
        RECT 2470.760 2946.110 2471.020 2946.430 ;
        RECT 2469.440 2898.685 2469.580 2946.110 ;
        RECT 2469.370 2898.315 2469.650 2898.685 ;
        RECT 2470.290 2898.315 2470.570 2898.685 ;
        RECT 2470.360 2863.210 2470.500 2898.315 ;
        RECT 2470.360 2863.070 2470.960 2863.210 ;
        RECT 2470.820 2849.530 2470.960 2863.070 ;
        RECT 2470.760 2849.210 2471.020 2849.530 ;
        RECT 2471.680 2815.210 2471.940 2815.530 ;
        RECT 2471.740 2801.445 2471.880 2815.210 ;
        RECT 2470.750 2801.075 2471.030 2801.445 ;
        RECT 2471.670 2801.075 2471.950 2801.445 ;
        RECT 2470.820 2753.310 2470.960 2801.075 ;
        RECT 2470.760 2752.990 2471.020 2753.310 ;
        RECT 2472.140 2752.990 2472.400 2753.310 ;
        RECT 2472.200 2719.310 2472.340 2752.990 ;
        RECT 2472.140 2718.990 2472.400 2719.310 ;
        RECT 2471.680 2718.310 2471.940 2718.630 ;
        RECT 2471.740 2704.885 2471.880 2718.310 ;
        RECT 2470.750 2704.515 2471.030 2704.885 ;
        RECT 2471.670 2704.515 2471.950 2704.885 ;
        RECT 2470.820 2656.750 2470.960 2704.515 ;
        RECT 2470.760 2656.430 2471.020 2656.750 ;
        RECT 2472.140 2656.430 2472.400 2656.750 ;
        RECT 2472.200 2619.010 2472.340 2656.430 ;
        RECT 1265.560 2618.690 1265.820 2619.010 ;
        RECT 2472.140 2618.690 2472.400 2619.010 ;
        RECT 1264.090 2599.370 1264.370 2600.000 ;
        RECT 1265.620 2599.370 1265.760 2618.690 ;
        RECT 1264.090 2599.230 1265.760 2599.370 ;
        RECT 1264.090 2596.000 1264.370 2599.230 ;
      LAYER via2 ;
        RECT 2474.430 3430.120 2474.710 3430.400 ;
        RECT 2471.210 3429.440 2471.490 3429.720 ;
        RECT 2469.370 2898.360 2469.650 2898.640 ;
        RECT 2470.290 2898.360 2470.570 2898.640 ;
        RECT 2470.750 2801.120 2471.030 2801.400 ;
        RECT 2471.670 2801.120 2471.950 2801.400 ;
        RECT 2470.750 2704.560 2471.030 2704.840 ;
        RECT 2471.670 2704.560 2471.950 2704.840 ;
      LAYER met3 ;
        RECT 2474.405 3430.410 2474.735 3430.425 ;
        RECT 2470.510 3430.110 2474.735 3430.410 ;
        RECT 2470.510 3429.730 2470.810 3430.110 ;
        RECT 2474.405 3430.095 2474.735 3430.110 ;
        RECT 2471.185 3429.730 2471.515 3429.745 ;
        RECT 2470.510 3429.430 2471.515 3429.730 ;
        RECT 2471.185 3429.415 2471.515 3429.430 ;
        RECT 2469.345 2898.650 2469.675 2898.665 ;
        RECT 2470.265 2898.650 2470.595 2898.665 ;
        RECT 2469.345 2898.350 2470.595 2898.650 ;
        RECT 2469.345 2898.335 2469.675 2898.350 ;
        RECT 2470.265 2898.335 2470.595 2898.350 ;
        RECT 2470.725 2801.410 2471.055 2801.425 ;
        RECT 2471.645 2801.410 2471.975 2801.425 ;
        RECT 2470.725 2801.110 2471.975 2801.410 ;
        RECT 2470.725 2801.095 2471.055 2801.110 ;
        RECT 2471.645 2801.095 2471.975 2801.110 ;
        RECT 2470.725 2704.850 2471.055 2704.865 ;
        RECT 2471.645 2704.850 2471.975 2704.865 ;
        RECT 2470.725 2704.550 2471.975 2704.850 ;
        RECT 2470.725 2704.535 2471.055 2704.550 ;
        RECT 2471.645 2704.535 2471.975 2704.550 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1679.990 3501.560 1680.310 3501.620 ;
        RECT 2149.190 3501.560 2149.510 3501.620 ;
        RECT 1679.990 3501.420 2149.510 3501.560 ;
        RECT 1679.990 3501.360 1680.310 3501.420 ;
        RECT 2149.190 3501.360 2149.510 3501.420 ;
        RECT 1289.910 3087.780 1290.230 3087.840 ;
        RECT 1679.990 3087.780 1680.310 3087.840 ;
        RECT 1289.910 3087.640 1680.310 3087.780 ;
        RECT 1289.910 3087.580 1290.230 3087.640 ;
        RECT 1679.990 3087.580 1680.310 3087.640 ;
      LAYER via ;
        RECT 1680.020 3501.360 1680.280 3501.620 ;
        RECT 2149.220 3501.360 2149.480 3501.620 ;
        RECT 1289.940 3087.580 1290.200 3087.840 ;
        RECT 1680.020 3087.580 1680.280 3087.840 ;
      LAYER met2 ;
        RECT 2149.070 3518.000 2149.630 3524.000 ;
        RECT 2149.280 3501.650 2149.420 3518.000 ;
        RECT 1680.020 3501.330 1680.280 3501.650 ;
        RECT 2149.220 3501.330 2149.480 3501.650 ;
        RECT 1680.080 3087.870 1680.220 3501.330 ;
        RECT 1289.940 3087.550 1290.200 3087.870 ;
        RECT 1680.020 3087.550 1680.280 3087.870 ;
        RECT 1290.000 2600.730 1290.140 3087.550 ;
        RECT 1290.000 2600.590 1290.600 2600.730 ;
        RECT 1289.850 2599.370 1290.130 2600.000 ;
        RECT 1290.460 2599.370 1290.600 2600.590 ;
        RECT 1289.850 2599.230 1290.600 2599.370 ;
        RECT 1289.850 2596.000 1290.130 2599.230 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1397.090 3500.540 1397.410 3500.600 ;
        RECT 1824.890 3500.540 1825.210 3500.600 ;
        RECT 1397.090 3500.400 1825.210 3500.540 ;
        RECT 1397.090 3500.340 1397.410 3500.400 ;
        RECT 1824.890 3500.340 1825.210 3500.400 ;
        RECT 1316.590 2619.600 1316.910 2619.660 ;
        RECT 1397.090 2619.600 1397.410 2619.660 ;
        RECT 1316.590 2619.460 1397.410 2619.600 ;
        RECT 1316.590 2619.400 1316.910 2619.460 ;
        RECT 1397.090 2619.400 1397.410 2619.460 ;
      LAYER via ;
        RECT 1397.120 3500.340 1397.380 3500.600 ;
        RECT 1824.920 3500.340 1825.180 3500.600 ;
        RECT 1316.620 2619.400 1316.880 2619.660 ;
        RECT 1397.120 2619.400 1397.380 2619.660 ;
      LAYER met2 ;
        RECT 1824.770 3518.000 1825.330 3524.000 ;
        RECT 1824.980 3500.630 1825.120 3518.000 ;
        RECT 1397.120 3500.310 1397.380 3500.630 ;
        RECT 1824.920 3500.310 1825.180 3500.630 ;
        RECT 1397.180 2619.690 1397.320 3500.310 ;
        RECT 1316.620 2619.370 1316.880 2619.690 ;
        RECT 1397.120 2619.370 1397.380 2619.690 ;
        RECT 1315.610 2599.370 1315.890 2600.000 ;
        RECT 1316.680 2599.370 1316.820 2619.370 ;
        RECT 1315.610 2599.230 1316.820 2599.370 ;
        RECT 1315.610 2596.000 1315.890 2599.230 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1499.285 3332.765 1499.455 3422.355 ;
        RECT 1498.365 3008.405 1498.535 3042.915 ;
        RECT 1498.825 2946.525 1498.995 2994.635 ;
      LAYER mcon ;
        RECT 1499.285 3422.185 1499.455 3422.355 ;
        RECT 1498.365 3042.745 1498.535 3042.915 ;
        RECT 1498.825 2994.465 1498.995 2994.635 ;
      LAYER met1 ;
        RECT 1498.290 3443.080 1498.610 3443.140 ;
        RECT 1500.590 3443.080 1500.910 3443.140 ;
        RECT 1498.290 3442.940 1500.910 3443.080 ;
        RECT 1498.290 3442.880 1498.610 3442.940 ;
        RECT 1500.590 3442.880 1500.910 3442.940 ;
        RECT 1497.830 3422.340 1498.150 3422.400 ;
        RECT 1499.225 3422.340 1499.515 3422.385 ;
        RECT 1497.830 3422.200 1499.515 3422.340 ;
        RECT 1497.830 3422.140 1498.150 3422.200 ;
        RECT 1499.225 3422.155 1499.515 3422.200 ;
        RECT 1499.225 3332.920 1499.515 3332.965 ;
        RECT 1499.670 3332.920 1499.990 3332.980 ;
        RECT 1499.225 3332.780 1499.990 3332.920 ;
        RECT 1499.225 3332.735 1499.515 3332.780 ;
        RECT 1499.670 3332.720 1499.990 3332.780 ;
        RECT 1498.290 3236.360 1498.610 3236.420 ;
        RECT 1498.750 3236.360 1499.070 3236.420 ;
        RECT 1498.290 3236.220 1499.070 3236.360 ;
        RECT 1498.290 3236.160 1498.610 3236.220 ;
        RECT 1498.750 3236.160 1499.070 3236.220 ;
        RECT 1498.290 3202.020 1498.610 3202.080 ;
        RECT 1498.750 3202.020 1499.070 3202.080 ;
        RECT 1498.290 3201.880 1499.070 3202.020 ;
        RECT 1498.290 3201.820 1498.610 3201.880 ;
        RECT 1498.750 3201.820 1499.070 3201.880 ;
        RECT 1497.830 3153.400 1498.150 3153.460 ;
        RECT 1498.750 3153.400 1499.070 3153.460 ;
        RECT 1497.830 3153.260 1499.070 3153.400 ;
        RECT 1497.830 3153.200 1498.150 3153.260 ;
        RECT 1498.750 3153.200 1499.070 3153.260 ;
        RECT 1497.830 3056.840 1498.150 3056.900 ;
        RECT 1498.750 3056.840 1499.070 3056.900 ;
        RECT 1497.830 3056.700 1499.070 3056.840 ;
        RECT 1497.830 3056.640 1498.150 3056.700 ;
        RECT 1498.750 3056.640 1499.070 3056.700 ;
        RECT 1498.290 3042.900 1498.610 3042.960 ;
        RECT 1498.095 3042.760 1498.610 3042.900 ;
        RECT 1498.290 3042.700 1498.610 3042.760 ;
        RECT 1498.305 3008.560 1498.595 3008.605 ;
        RECT 1499.210 3008.560 1499.530 3008.620 ;
        RECT 1498.305 3008.420 1499.530 3008.560 ;
        RECT 1498.305 3008.375 1498.595 3008.420 ;
        RECT 1499.210 3008.360 1499.530 3008.420 ;
        RECT 1498.765 2994.620 1499.055 2994.665 ;
        RECT 1499.210 2994.620 1499.530 2994.680 ;
        RECT 1498.765 2994.480 1499.530 2994.620 ;
        RECT 1498.765 2994.435 1499.055 2994.480 ;
        RECT 1499.210 2994.420 1499.530 2994.480 ;
        RECT 1498.750 2946.680 1499.070 2946.740 ;
        RECT 1498.555 2946.540 1499.070 2946.680 ;
        RECT 1498.750 2946.480 1499.070 2946.540 ;
        RECT 1498.750 2911.800 1499.070 2912.060 ;
        RECT 1498.840 2911.320 1498.980 2911.800 ;
        RECT 1499.210 2911.320 1499.530 2911.380 ;
        RECT 1498.840 2911.180 1499.530 2911.320 ;
        RECT 1499.210 2911.120 1499.530 2911.180 ;
        RECT 1497.370 2863.720 1497.690 2863.780 ;
        RECT 1499.210 2863.720 1499.530 2863.780 ;
        RECT 1497.370 2863.580 1499.530 2863.720 ;
        RECT 1497.370 2863.520 1497.690 2863.580 ;
        RECT 1499.210 2863.520 1499.530 2863.580 ;
        RECT 1497.370 2766.820 1497.690 2766.880 ;
        RECT 1499.670 2766.820 1499.990 2766.880 ;
        RECT 1497.370 2766.680 1499.990 2766.820 ;
        RECT 1497.370 2766.620 1497.690 2766.680 ;
        RECT 1499.670 2766.620 1499.990 2766.680 ;
        RECT 1499.670 2719.220 1499.990 2719.280 ;
        RECT 1499.300 2719.080 1499.990 2719.220 ;
        RECT 1499.300 2718.600 1499.440 2719.080 ;
        RECT 1499.670 2719.020 1499.990 2719.080 ;
        RECT 1499.210 2718.340 1499.530 2718.600 ;
        RECT 1498.290 2656.660 1498.610 2656.720 ;
        RECT 1499.670 2656.660 1499.990 2656.720 ;
        RECT 1498.290 2656.520 1499.990 2656.660 ;
        RECT 1498.290 2656.460 1498.610 2656.520 ;
        RECT 1499.670 2656.460 1499.990 2656.520 ;
        RECT 1342.810 2619.260 1343.130 2619.320 ;
        RECT 1499.670 2619.260 1499.990 2619.320 ;
        RECT 1342.810 2619.120 1499.990 2619.260 ;
        RECT 1342.810 2619.060 1343.130 2619.120 ;
        RECT 1499.670 2619.060 1499.990 2619.120 ;
      LAYER via ;
        RECT 1498.320 3442.880 1498.580 3443.140 ;
        RECT 1500.620 3442.880 1500.880 3443.140 ;
        RECT 1497.860 3422.140 1498.120 3422.400 ;
        RECT 1499.700 3332.720 1499.960 3332.980 ;
        RECT 1498.320 3236.160 1498.580 3236.420 ;
        RECT 1498.780 3236.160 1499.040 3236.420 ;
        RECT 1498.320 3201.820 1498.580 3202.080 ;
        RECT 1498.780 3201.820 1499.040 3202.080 ;
        RECT 1497.860 3153.200 1498.120 3153.460 ;
        RECT 1498.780 3153.200 1499.040 3153.460 ;
        RECT 1497.860 3056.640 1498.120 3056.900 ;
        RECT 1498.780 3056.640 1499.040 3056.900 ;
        RECT 1498.320 3042.700 1498.580 3042.960 ;
        RECT 1499.240 3008.360 1499.500 3008.620 ;
        RECT 1499.240 2994.420 1499.500 2994.680 ;
        RECT 1498.780 2946.480 1499.040 2946.740 ;
        RECT 1498.780 2911.800 1499.040 2912.060 ;
        RECT 1499.240 2911.120 1499.500 2911.380 ;
        RECT 1497.400 2863.520 1497.660 2863.780 ;
        RECT 1499.240 2863.520 1499.500 2863.780 ;
        RECT 1497.400 2766.620 1497.660 2766.880 ;
        RECT 1499.700 2766.620 1499.960 2766.880 ;
        RECT 1499.700 2719.020 1499.960 2719.280 ;
        RECT 1499.240 2718.340 1499.500 2718.600 ;
        RECT 1498.320 2656.460 1498.580 2656.720 ;
        RECT 1499.700 2656.460 1499.960 2656.720 ;
        RECT 1342.840 2619.060 1343.100 2619.320 ;
        RECT 1499.700 2619.060 1499.960 2619.320 ;
      LAYER met2 ;
        RECT 1500.470 3518.000 1501.030 3524.000 ;
        RECT 1500.680 3443.170 1500.820 3518.000 ;
        RECT 1498.320 3442.850 1498.580 3443.170 ;
        RECT 1500.620 3442.850 1500.880 3443.170 ;
        RECT 1498.380 3429.650 1498.520 3442.850 ;
        RECT 1497.920 3429.510 1498.520 3429.650 ;
        RECT 1497.920 3422.430 1498.060 3429.510 ;
        RECT 1497.860 3422.110 1498.120 3422.430 ;
        RECT 1499.700 3332.690 1499.960 3333.010 ;
        RECT 1499.760 3298.410 1499.900 3332.690 ;
        RECT 1498.840 3298.270 1499.900 3298.410 ;
        RECT 1498.840 3236.450 1498.980 3298.270 ;
        RECT 1498.320 3236.130 1498.580 3236.450 ;
        RECT 1498.780 3236.130 1499.040 3236.450 ;
        RECT 1498.380 3202.110 1498.520 3236.130 ;
        RECT 1498.320 3201.790 1498.580 3202.110 ;
        RECT 1498.780 3201.790 1499.040 3202.110 ;
        RECT 1498.840 3153.490 1498.980 3201.790 ;
        RECT 1497.860 3153.170 1498.120 3153.490 ;
        RECT 1498.780 3153.170 1499.040 3153.490 ;
        RECT 1497.920 3152.890 1498.060 3153.170 ;
        RECT 1497.920 3152.750 1498.520 3152.890 ;
        RECT 1498.380 3105.290 1498.520 3152.750 ;
        RECT 1498.380 3105.150 1498.980 3105.290 ;
        RECT 1498.840 3056.930 1498.980 3105.150 ;
        RECT 1497.860 3056.610 1498.120 3056.930 ;
        RECT 1498.780 3056.610 1499.040 3056.930 ;
        RECT 1497.920 3056.330 1498.060 3056.610 ;
        RECT 1497.920 3056.190 1498.520 3056.330 ;
        RECT 1498.380 3042.990 1498.520 3056.190 ;
        RECT 1498.320 3042.670 1498.580 3042.990 ;
        RECT 1499.240 3008.330 1499.500 3008.650 ;
        RECT 1499.300 2994.710 1499.440 3008.330 ;
        RECT 1499.240 2994.390 1499.500 2994.710 ;
        RECT 1498.780 2946.450 1499.040 2946.770 ;
        RECT 1498.840 2912.090 1498.980 2946.450 ;
        RECT 1498.780 2911.770 1499.040 2912.090 ;
        RECT 1499.240 2911.090 1499.500 2911.410 ;
        RECT 1499.300 2863.810 1499.440 2911.090 ;
        RECT 1497.400 2863.490 1497.660 2863.810 ;
        RECT 1499.240 2863.490 1499.500 2863.810 ;
        RECT 1497.460 2766.910 1497.600 2863.490 ;
        RECT 1497.400 2766.590 1497.660 2766.910 ;
        RECT 1499.700 2766.590 1499.960 2766.910 ;
        RECT 1499.760 2719.310 1499.900 2766.590 ;
        RECT 1499.700 2718.990 1499.960 2719.310 ;
        RECT 1499.240 2718.310 1499.500 2718.630 ;
        RECT 1499.300 2704.885 1499.440 2718.310 ;
        RECT 1498.310 2704.515 1498.590 2704.885 ;
        RECT 1499.230 2704.515 1499.510 2704.885 ;
        RECT 1498.380 2656.750 1498.520 2704.515 ;
        RECT 1498.320 2656.430 1498.580 2656.750 ;
        RECT 1499.700 2656.430 1499.960 2656.750 ;
        RECT 1499.760 2619.350 1499.900 2656.430 ;
        RECT 1342.840 2619.030 1343.100 2619.350 ;
        RECT 1499.700 2619.030 1499.960 2619.350 ;
        RECT 1341.370 2599.370 1341.650 2600.000 ;
        RECT 1342.900 2599.370 1343.040 2619.030 ;
        RECT 1341.370 2599.230 1343.040 2599.370 ;
        RECT 1341.370 2596.000 1341.650 2599.230 ;
      LAYER via2 ;
        RECT 1498.310 2704.560 1498.590 2704.840 ;
        RECT 1499.230 2704.560 1499.510 2704.840 ;
      LAYER met3 ;
        RECT 1498.285 2704.850 1498.615 2704.865 ;
        RECT 1499.205 2704.850 1499.535 2704.865 ;
        RECT 1498.285 2704.550 1499.535 2704.850 ;
        RECT 1498.285 2704.535 1498.615 2704.550 ;
        RECT 1499.205 2704.535 1499.535 2704.550 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 880.990 2608.635 881.270 2609.005 ;
        RECT 2901.310 2608.635 2901.590 2609.005 ;
        RECT 879.530 2599.370 879.810 2600.000 ;
        RECT 881.060 2599.370 881.200 2608.635 ;
        RECT 879.530 2599.230 881.200 2599.370 ;
        RECT 879.530 2596.000 879.810 2599.230 ;
        RECT 2901.380 322.845 2901.520 2608.635 ;
        RECT 2901.310 322.475 2901.590 322.845 ;
      LAYER via2 ;
        RECT 880.990 2608.680 881.270 2608.960 ;
        RECT 2901.310 2608.680 2901.590 2608.960 ;
        RECT 2901.310 322.520 2901.590 322.800 ;
      LAYER met3 ;
        RECT 880.965 2608.970 881.295 2608.985 ;
        RECT 2901.285 2608.970 2901.615 2608.985 ;
        RECT 880.965 2608.670 2901.615 2608.970 ;
        RECT 880.965 2608.655 881.295 2608.670 ;
        RECT 2901.285 2608.655 2901.615 2608.670 ;
        RECT 2901.285 322.810 2901.615 322.825 ;
        RECT 2918.000 322.810 2924.000 323.260 ;
        RECT 2901.285 322.510 2924.000 322.810 ;
        RECT 2901.285 322.495 2901.615 322.510 ;
        RECT 2918.000 322.060 2924.000 322.510 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1175.830 3498.840 1176.150 3498.900 ;
        RECT 1366.270 3498.840 1366.590 3498.900 ;
        RECT 1175.830 3498.700 1366.590 3498.840 ;
        RECT 1175.830 3498.640 1176.150 3498.700 ;
        RECT 1366.270 3498.640 1366.590 3498.700 ;
      LAYER via ;
        RECT 1175.860 3498.640 1176.120 3498.900 ;
        RECT 1366.300 3498.640 1366.560 3498.900 ;
      LAYER met2 ;
        RECT 1175.710 3518.000 1176.270 3524.000 ;
        RECT 1175.920 3498.930 1176.060 3518.000 ;
        RECT 1175.860 3498.610 1176.120 3498.930 ;
        RECT 1366.300 3498.610 1366.560 3498.930 ;
        RECT 1366.360 2600.050 1366.500 3498.610 ;
        RECT 1366.360 2600.000 1366.890 2600.050 ;
        RECT 1366.360 2599.910 1366.950 2600.000 ;
        RECT 1366.670 2596.000 1366.950 2599.910 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 851.530 3500.540 851.850 3500.600 ;
        RECT 1386.970 3500.540 1387.290 3500.600 ;
        RECT 851.530 3500.400 1387.290 3500.540 ;
        RECT 851.530 3500.340 851.850 3500.400 ;
        RECT 1386.970 3500.340 1387.290 3500.400 ;
      LAYER via ;
        RECT 851.560 3500.340 851.820 3500.600 ;
        RECT 1387.000 3500.340 1387.260 3500.600 ;
      LAYER met2 ;
        RECT 851.410 3518.000 851.970 3524.000 ;
        RECT 851.620 3500.630 851.760 3518.000 ;
        RECT 851.560 3500.310 851.820 3500.630 ;
        RECT 1387.000 3500.310 1387.260 3500.630 ;
        RECT 1387.060 2600.730 1387.200 3500.310 ;
        RECT 1387.060 2600.590 1391.340 2600.730 ;
        RECT 1391.200 2600.050 1391.340 2600.590 ;
        RECT 1391.200 2600.000 1392.650 2600.050 ;
        RECT 1391.200 2599.910 1392.710 2600.000 ;
        RECT 1392.430 2596.000 1392.710 2599.910 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 527.230 3504.280 527.550 3504.340 ;
        RECT 1415.030 3504.280 1415.350 3504.340 ;
        RECT 527.230 3504.140 1415.350 3504.280 ;
        RECT 527.230 3504.080 527.550 3504.140 ;
        RECT 1415.030 3504.080 1415.350 3504.140 ;
      LAYER via ;
        RECT 527.260 3504.080 527.520 3504.340 ;
        RECT 1415.060 3504.080 1415.320 3504.340 ;
      LAYER met2 ;
        RECT 527.110 3518.000 527.670 3524.000 ;
        RECT 527.320 3504.370 527.460 3518.000 ;
        RECT 527.260 3504.050 527.520 3504.370 ;
        RECT 1415.060 3504.050 1415.320 3504.370 ;
        RECT 1415.120 2600.050 1415.260 3504.050 ;
        RECT 1415.120 2600.000 1418.410 2600.050 ;
        RECT 1415.120 2599.910 1418.470 2600.000 ;
        RECT 1418.190 2596.000 1418.470 2599.910 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 202.470 3502.580 202.790 3502.640 ;
        RECT 1442.170 3502.580 1442.490 3502.640 ;
        RECT 202.470 3502.440 1442.490 3502.580 ;
        RECT 202.470 3502.380 202.790 3502.440 ;
        RECT 1442.170 3502.380 1442.490 3502.440 ;
      LAYER via ;
        RECT 202.500 3502.380 202.760 3502.640 ;
        RECT 1442.200 3502.380 1442.460 3502.640 ;
      LAYER met2 ;
        RECT 202.350 3518.000 202.910 3524.000 ;
        RECT 202.560 3502.670 202.700 3518.000 ;
        RECT 202.500 3502.350 202.760 3502.670 ;
        RECT 1442.200 3502.350 1442.460 3502.670 ;
        RECT 1442.260 2600.050 1442.400 3502.350 ;
        RECT 1442.260 2600.000 1444.170 2600.050 ;
        RECT 1442.260 2599.910 1444.230 2600.000 ;
        RECT 1443.950 2596.000 1444.230 2599.910 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.550 3408.740 17.870 3408.800 ;
        RECT 1462.870 3408.740 1463.190 3408.800 ;
        RECT 17.550 3408.600 1463.190 3408.740 ;
        RECT 17.550 3408.540 17.870 3408.600 ;
        RECT 1462.870 3408.540 1463.190 3408.600 ;
        RECT 1462.870 2740.300 1463.190 2740.360 ;
        RECT 1466.550 2740.300 1466.870 2740.360 ;
        RECT 1462.870 2740.160 1466.870 2740.300 ;
        RECT 1462.870 2740.100 1463.190 2740.160 ;
        RECT 1466.550 2740.100 1466.870 2740.160 ;
        RECT 1466.550 2656.660 1466.870 2656.720 ;
        RECT 1467.470 2656.660 1467.790 2656.720 ;
        RECT 1466.550 2656.520 1467.790 2656.660 ;
        RECT 1466.550 2656.460 1466.870 2656.520 ;
        RECT 1467.470 2656.460 1467.790 2656.520 ;
      LAYER via ;
        RECT 17.580 3408.540 17.840 3408.800 ;
        RECT 1462.900 3408.540 1463.160 3408.800 ;
        RECT 1462.900 2740.100 1463.160 2740.360 ;
        RECT 1466.580 2740.100 1466.840 2740.360 ;
        RECT 1466.580 2656.460 1466.840 2656.720 ;
        RECT 1467.500 2656.460 1467.760 2656.720 ;
      LAYER met2 ;
        RECT 17.570 3411.035 17.850 3411.405 ;
        RECT 17.640 3408.830 17.780 3411.035 ;
        RECT 17.580 3408.510 17.840 3408.830 ;
        RECT 1462.900 3408.510 1463.160 3408.830 ;
        RECT 1462.960 2740.390 1463.100 3408.510 ;
        RECT 1462.900 2740.070 1463.160 2740.390 ;
        RECT 1466.580 2740.070 1466.840 2740.390 ;
        RECT 1466.640 2656.750 1466.780 2740.070 ;
        RECT 1466.580 2656.605 1466.840 2656.750 ;
        RECT 1467.500 2656.605 1467.760 2656.750 ;
        RECT 1466.570 2656.235 1466.850 2656.605 ;
        RECT 1467.490 2656.235 1467.770 2656.605 ;
        RECT 1466.640 2600.050 1466.780 2656.235 ;
        RECT 1466.640 2600.000 1469.470 2600.050 ;
        RECT 1466.640 2599.910 1469.530 2600.000 ;
        RECT 1469.250 2596.000 1469.530 2599.910 ;
      LAYER via2 ;
        RECT 17.570 3411.080 17.850 3411.360 ;
        RECT 1466.570 2656.280 1466.850 2656.560 ;
        RECT 1467.490 2656.280 1467.770 2656.560 ;
      LAYER met3 ;
        RECT -4.000 3411.370 2.000 3411.820 ;
        RECT 17.545 3411.370 17.875 3411.385 ;
        RECT -4.000 3411.070 17.875 3411.370 ;
        RECT -4.000 3410.620 2.000 3411.070 ;
        RECT 17.545 3411.055 17.875 3411.070 ;
        RECT 1466.545 2656.570 1466.875 2656.585 ;
        RECT 1467.465 2656.570 1467.795 2656.585 ;
        RECT 1466.545 2656.270 1467.795 2656.570 ;
        RECT 1466.545 2656.255 1466.875 2656.270 ;
        RECT 1467.465 2656.255 1467.795 2656.270 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 3119.060 17.410 3119.120 ;
        RECT 1490.470 3119.060 1490.790 3119.120 ;
        RECT 17.090 3118.920 1490.790 3119.060 ;
        RECT 17.090 3118.860 17.410 3118.920 ;
        RECT 1490.470 3118.860 1490.790 3118.920 ;
      LAYER via ;
        RECT 17.120 3118.860 17.380 3119.120 ;
        RECT 1490.500 3118.860 1490.760 3119.120 ;
      LAYER met2 ;
        RECT 17.110 3124.075 17.390 3124.445 ;
        RECT 17.180 3119.150 17.320 3124.075 ;
        RECT 17.120 3118.830 17.380 3119.150 ;
        RECT 1490.500 3118.830 1490.760 3119.150 ;
        RECT 1490.560 2600.730 1490.700 3118.830 ;
        RECT 1490.560 2600.590 1493.000 2600.730 ;
        RECT 1492.860 2600.050 1493.000 2600.590 ;
        RECT 1492.860 2600.000 1495.230 2600.050 ;
        RECT 1492.860 2599.910 1495.290 2600.000 ;
        RECT 1495.010 2596.000 1495.290 2599.910 ;
      LAYER via2 ;
        RECT 17.110 3124.120 17.390 3124.400 ;
      LAYER met3 ;
        RECT -4.000 3124.410 2.000 3124.860 ;
        RECT 17.085 3124.410 17.415 3124.425 ;
        RECT -4.000 3124.110 17.415 3124.410 ;
        RECT -4.000 3123.660 2.000 3124.110 ;
        RECT 17.085 3124.095 17.415 3124.110 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 2836.180 17.410 2836.240 ;
        RECT 1518.070 2836.180 1518.390 2836.240 ;
        RECT 17.090 2836.040 1518.390 2836.180 ;
        RECT 17.090 2835.980 17.410 2836.040 ;
        RECT 1518.070 2835.980 1518.390 2836.040 ;
      LAYER via ;
        RECT 17.120 2835.980 17.380 2836.240 ;
        RECT 1518.100 2835.980 1518.360 2836.240 ;
      LAYER met2 ;
        RECT 17.110 2836.435 17.390 2836.805 ;
        RECT 17.180 2836.270 17.320 2836.435 ;
        RECT 17.120 2835.950 17.380 2836.270 ;
        RECT 1518.100 2835.950 1518.360 2836.270 ;
        RECT 1518.160 2600.050 1518.300 2835.950 ;
        RECT 1518.160 2600.000 1520.990 2600.050 ;
        RECT 1518.160 2599.910 1521.050 2600.000 ;
        RECT 1520.770 2596.000 1521.050 2599.910 ;
      LAYER via2 ;
        RECT 17.110 2836.480 17.390 2836.760 ;
      LAYER met3 ;
        RECT -4.000 2836.770 2.000 2837.220 ;
        RECT 17.085 2836.770 17.415 2836.785 ;
        RECT -4.000 2836.470 17.415 2836.770 ;
        RECT -4.000 2836.020 2.000 2836.470 ;
        RECT 17.085 2836.455 17.415 2836.470 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 14.790 2613.820 15.110 2613.880 ;
        RECT 1545.670 2613.820 1545.990 2613.880 ;
        RECT 14.790 2613.680 1545.990 2613.820 ;
        RECT 14.790 2613.620 15.110 2613.680 ;
        RECT 1545.670 2613.620 1545.990 2613.680 ;
      LAYER via ;
        RECT 14.820 2613.620 15.080 2613.880 ;
        RECT 1545.700 2613.620 1545.960 2613.880 ;
      LAYER met2 ;
        RECT 14.820 2613.590 15.080 2613.910 ;
        RECT 1545.700 2613.590 1545.960 2613.910 ;
        RECT 14.880 2549.845 15.020 2613.590 ;
        RECT 1545.760 2600.050 1545.900 2613.590 ;
        RECT 1545.760 2600.000 1546.750 2600.050 ;
        RECT 1545.760 2599.910 1546.810 2600.000 ;
        RECT 1546.530 2596.000 1546.810 2599.910 ;
        RECT 14.810 2549.475 15.090 2549.845 ;
      LAYER via2 ;
        RECT 14.810 2549.520 15.090 2549.800 ;
      LAYER met3 ;
        RECT -4.000 2549.810 2.000 2550.260 ;
        RECT 14.785 2549.810 15.115 2549.825 ;
        RECT -4.000 2549.510 15.115 2549.810 ;
        RECT -4.000 2549.060 2.000 2549.510 ;
        RECT 14.785 2549.495 15.115 2549.510 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 31.810 2597.500 32.130 2597.560 ;
        RECT 1570.510 2597.500 1570.830 2597.560 ;
        RECT 31.810 2597.360 1570.830 2597.500 ;
        RECT 31.810 2597.300 32.130 2597.360 ;
        RECT 1570.510 2597.300 1570.830 2597.360 ;
        RECT 15.250 2262.260 15.570 2262.320 ;
        RECT 31.810 2262.260 32.130 2262.320 ;
        RECT 15.250 2262.120 32.130 2262.260 ;
        RECT 15.250 2262.060 15.570 2262.120 ;
        RECT 31.810 2262.060 32.130 2262.120 ;
      LAYER via ;
        RECT 31.840 2597.300 32.100 2597.560 ;
        RECT 1570.540 2597.300 1570.800 2597.560 ;
        RECT 15.280 2262.060 15.540 2262.320 ;
        RECT 31.840 2262.060 32.100 2262.320 ;
      LAYER met2 ;
        RECT 31.840 2597.270 32.100 2597.590 ;
        RECT 1570.540 2597.330 1570.800 2597.590 ;
        RECT 1571.830 2597.330 1572.110 2600.000 ;
        RECT 1570.540 2597.270 1572.110 2597.330 ;
        RECT 31.900 2262.350 32.040 2597.270 ;
        RECT 1570.600 2597.190 1572.110 2597.270 ;
        RECT 1571.830 2596.000 1572.110 2597.190 ;
        RECT 15.280 2262.205 15.540 2262.350 ;
        RECT 15.270 2261.835 15.550 2262.205 ;
        RECT 31.840 2262.030 32.100 2262.350 ;
      LAYER via2 ;
        RECT 15.270 2261.880 15.550 2262.160 ;
      LAYER met3 ;
        RECT -4.000 2262.170 2.000 2262.620 ;
        RECT 15.245 2262.170 15.575 2262.185 ;
        RECT -4.000 2261.870 15.575 2262.170 ;
        RECT -4.000 2261.420 2.000 2261.870 ;
        RECT 15.245 2261.855 15.575 2261.870 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 16.170 2612.460 16.490 2612.520 ;
        RECT 1596.270 2612.460 1596.590 2612.520 ;
        RECT 16.170 2612.320 1596.590 2612.460 ;
        RECT 16.170 2612.260 16.490 2612.320 ;
        RECT 1596.270 2612.260 1596.590 2612.320 ;
      LAYER via ;
        RECT 16.200 2612.260 16.460 2612.520 ;
        RECT 1596.300 2612.260 1596.560 2612.520 ;
      LAYER met2 ;
        RECT 16.200 2612.230 16.460 2612.550 ;
        RECT 1596.300 2612.230 1596.560 2612.550 ;
        RECT 16.260 1975.245 16.400 2612.230 ;
        RECT 1596.360 2600.050 1596.500 2612.230 ;
        RECT 1596.360 2600.000 1597.810 2600.050 ;
        RECT 1596.360 2599.910 1597.870 2600.000 ;
        RECT 1597.590 2596.000 1597.870 2599.910 ;
        RECT 16.190 1974.875 16.470 1975.245 ;
      LAYER via2 ;
        RECT 16.190 1974.920 16.470 1975.200 ;
      LAYER met3 ;
        RECT -4.000 1975.210 2.000 1975.660 ;
        RECT 16.165 1975.210 16.495 1975.225 ;
        RECT -4.000 1974.910 16.495 1975.210 ;
        RECT -4.000 1974.460 2.000 1974.910 ;
        RECT 16.165 1974.895 16.495 1974.910 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 906.750 2609.995 907.030 2610.365 ;
        RECT 2903.150 2609.995 2903.430 2610.365 ;
        RECT 905.290 2599.370 905.570 2600.000 ;
        RECT 906.820 2599.370 906.960 2609.995 ;
        RECT 905.290 2599.230 906.960 2599.370 ;
        RECT 905.290 2596.000 905.570 2599.230 ;
        RECT 2903.220 557.445 2903.360 2609.995 ;
        RECT 2903.150 557.075 2903.430 557.445 ;
      LAYER via2 ;
        RECT 906.750 2610.040 907.030 2610.320 ;
        RECT 2903.150 2610.040 2903.430 2610.320 ;
        RECT 2903.150 557.120 2903.430 557.400 ;
      LAYER met3 ;
        RECT 906.725 2610.330 907.055 2610.345 ;
        RECT 2903.125 2610.330 2903.455 2610.345 ;
        RECT 906.725 2610.030 2903.455 2610.330 ;
        RECT 906.725 2610.015 907.055 2610.030 ;
        RECT 2903.125 2610.015 2903.455 2610.030 ;
        RECT 2903.125 557.410 2903.455 557.425 ;
        RECT 2918.000 557.410 2924.000 557.860 ;
        RECT 2903.125 557.110 2924.000 557.410 ;
        RECT 2903.125 557.095 2903.455 557.110 ;
        RECT 2918.000 556.660 2924.000 557.110 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 16.630 2596.820 16.950 2596.880 ;
        RECT 1622.030 2596.820 1622.350 2596.880 ;
        RECT 16.630 2596.680 1622.350 2596.820 ;
        RECT 16.630 2596.620 16.950 2596.680 ;
        RECT 1622.030 2596.620 1622.350 2596.680 ;
      LAYER via ;
        RECT 16.660 2596.620 16.920 2596.880 ;
        RECT 1622.060 2596.620 1622.320 2596.880 ;
      LAYER met2 ;
        RECT 16.660 2596.590 16.920 2596.910 ;
        RECT 1622.060 2596.650 1622.320 2596.910 ;
        RECT 1623.350 2596.650 1623.630 2600.000 ;
        RECT 1622.060 2596.590 1623.630 2596.650 ;
        RECT 16.720 1687.605 16.860 2596.590 ;
        RECT 1622.120 2596.510 1623.630 2596.590 ;
        RECT 1623.350 2596.000 1623.630 2596.510 ;
        RECT 16.650 1687.235 16.930 1687.605 ;
      LAYER via2 ;
        RECT 16.650 1687.280 16.930 1687.560 ;
      LAYER met3 ;
        RECT -4.000 1687.570 2.000 1688.020 ;
        RECT 16.625 1687.570 16.955 1687.585 ;
        RECT -4.000 1687.270 16.955 1687.570 ;
        RECT -4.000 1686.820 2.000 1687.270 ;
        RECT 16.625 1687.255 16.955 1687.270 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 19.850 2596.480 20.170 2596.540 ;
        RECT 1648.250 2596.480 1648.570 2596.540 ;
        RECT 19.850 2596.340 1648.570 2596.480 ;
        RECT 19.850 2596.280 20.170 2596.340 ;
        RECT 1648.250 2596.280 1648.570 2596.340 ;
      LAYER via ;
        RECT 19.880 2596.280 20.140 2596.540 ;
        RECT 1648.280 2596.280 1648.540 2596.540 ;
      LAYER met2 ;
        RECT 1649.110 2596.650 1649.390 2600.000 ;
        RECT 1648.340 2596.570 1649.390 2596.650 ;
        RECT 19.880 2596.250 20.140 2596.570 ;
        RECT 1648.280 2596.510 1649.390 2596.570 ;
        RECT 1648.280 2596.250 1648.540 2596.510 ;
        RECT 19.940 1472.045 20.080 2596.250 ;
        RECT 1649.110 2596.000 1649.390 2596.510 ;
        RECT 19.870 1471.675 20.150 1472.045 ;
      LAYER via2 ;
        RECT 19.870 1471.720 20.150 1472.000 ;
      LAYER met3 ;
        RECT -4.000 1472.010 2.000 1472.460 ;
        RECT 19.845 1472.010 20.175 1472.025 ;
        RECT -4.000 1471.710 20.175 1472.010 ;
        RECT -4.000 1471.260 2.000 1471.710 ;
        RECT 19.845 1471.695 20.175 1471.710 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 19.390 2609.400 19.710 2609.460 ;
        RECT 1672.630 2609.400 1672.950 2609.460 ;
        RECT 19.390 2609.260 1672.950 2609.400 ;
        RECT 19.390 2609.200 19.710 2609.260 ;
        RECT 1672.630 2609.200 1672.950 2609.260 ;
      LAYER via ;
        RECT 19.420 2609.200 19.680 2609.460 ;
        RECT 1672.660 2609.200 1672.920 2609.460 ;
      LAYER met2 ;
        RECT 19.420 2609.170 19.680 2609.490 ;
        RECT 1672.660 2609.170 1672.920 2609.490 ;
        RECT 19.480 1256.485 19.620 2609.170 ;
        RECT 1672.720 2600.050 1672.860 2609.170 ;
        RECT 1672.720 2600.000 1674.630 2600.050 ;
        RECT 1672.720 2599.910 1674.690 2600.000 ;
        RECT 1674.410 2596.000 1674.690 2599.910 ;
        RECT 19.410 1256.115 19.690 1256.485 ;
      LAYER via2 ;
        RECT 19.410 1256.160 19.690 1256.440 ;
      LAYER met3 ;
        RECT -4.000 1256.450 2.000 1256.900 ;
        RECT 19.385 1256.450 19.715 1256.465 ;
        RECT -4.000 1256.150 19.715 1256.450 ;
        RECT -4.000 1255.700 2.000 1256.150 ;
        RECT 19.385 1256.135 19.715 1256.150 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 86.165 2595.985 86.335 2597.855 ;
        RECT 113.765 2595.985 113.935 2597.855 ;
        RECT 182.765 2595.985 182.935 2597.855 ;
        RECT 210.365 2595.985 210.535 2597.855 ;
        RECT 279.365 2595.985 279.535 2597.855 ;
        RECT 306.965 2595.985 307.135 2597.855 ;
        RECT 375.965 2595.985 376.135 2597.855 ;
        RECT 403.565 2595.985 403.735 2597.855 ;
        RECT 472.565 2595.985 472.735 2597.855 ;
        RECT 500.165 2595.985 500.335 2597.855 ;
        RECT 569.165 2595.985 569.335 2597.855 ;
        RECT 596.765 2595.985 596.935 2597.855 ;
        RECT 665.765 2595.985 665.935 2597.855 ;
        RECT 693.365 2595.985 693.535 2597.855 ;
        RECT 762.365 2595.985 762.535 2597.855 ;
        RECT 789.965 2595.985 790.135 2597.855 ;
        RECT 858.965 2595.985 859.135 2598.195 ;
        RECT 907.265 2595.985 907.435 2598.195 ;
        RECT 950.045 2595.985 950.215 2597.855 ;
        RECT 979.945 2595.985 980.115 2597.855 ;
        RECT 1048.945 2595.985 1049.115 2598.195 ;
        RECT 1096.785 2595.985 1096.955 2598.195 ;
        RECT 1526.885 2595.985 1527.055 2598.195 ;
        RECT 1584.385 2595.985 1584.555 2598.195 ;
        RECT 1628.545 2595.985 1628.715 2596.835 ;
      LAYER mcon ;
        RECT 858.965 2598.025 859.135 2598.195 ;
        RECT 86.165 2597.685 86.335 2597.855 ;
        RECT 113.765 2597.685 113.935 2597.855 ;
        RECT 182.765 2597.685 182.935 2597.855 ;
        RECT 210.365 2597.685 210.535 2597.855 ;
        RECT 279.365 2597.685 279.535 2597.855 ;
        RECT 306.965 2597.685 307.135 2597.855 ;
        RECT 375.965 2597.685 376.135 2597.855 ;
        RECT 403.565 2597.685 403.735 2597.855 ;
        RECT 472.565 2597.685 472.735 2597.855 ;
        RECT 500.165 2597.685 500.335 2597.855 ;
        RECT 569.165 2597.685 569.335 2597.855 ;
        RECT 596.765 2597.685 596.935 2597.855 ;
        RECT 665.765 2597.685 665.935 2597.855 ;
        RECT 693.365 2597.685 693.535 2597.855 ;
        RECT 762.365 2597.685 762.535 2597.855 ;
        RECT 789.965 2597.685 790.135 2597.855 ;
        RECT 907.265 2598.025 907.435 2598.195 ;
        RECT 1048.945 2598.025 1049.115 2598.195 ;
        RECT 950.045 2597.685 950.215 2597.855 ;
        RECT 979.945 2597.685 980.115 2597.855 ;
        RECT 1096.785 2598.025 1096.955 2598.195 ;
        RECT 1526.885 2598.025 1527.055 2598.195 ;
        RECT 1584.385 2598.025 1584.555 2598.195 ;
        RECT 1628.545 2596.665 1628.715 2596.835 ;
      LAYER met1 ;
        RECT 858.905 2598.180 859.195 2598.225 ;
        RECT 907.205 2598.180 907.495 2598.225 ;
        RECT 858.905 2598.040 907.495 2598.180 ;
        RECT 858.905 2597.995 859.195 2598.040 ;
        RECT 907.205 2597.995 907.495 2598.040 ;
        RECT 1048.885 2598.180 1049.175 2598.225 ;
        RECT 1096.725 2598.180 1097.015 2598.225 ;
        RECT 1048.885 2598.040 1097.015 2598.180 ;
        RECT 1048.885 2597.995 1049.175 2598.040 ;
        RECT 1096.725 2597.995 1097.015 2598.040 ;
        RECT 1526.825 2598.180 1527.115 2598.225 ;
        RECT 1584.325 2598.180 1584.615 2598.225 ;
        RECT 1526.825 2598.040 1584.615 2598.180 ;
        RECT 1526.825 2597.995 1527.115 2598.040 ;
        RECT 1584.325 2597.995 1584.615 2598.040 ;
        RECT 86.105 2597.840 86.395 2597.885 ;
        RECT 113.705 2597.840 113.995 2597.885 ;
        RECT 86.105 2597.700 113.995 2597.840 ;
        RECT 86.105 2597.655 86.395 2597.700 ;
        RECT 113.705 2597.655 113.995 2597.700 ;
        RECT 182.705 2597.840 182.995 2597.885 ;
        RECT 210.305 2597.840 210.595 2597.885 ;
        RECT 182.705 2597.700 210.595 2597.840 ;
        RECT 182.705 2597.655 182.995 2597.700 ;
        RECT 210.305 2597.655 210.595 2597.700 ;
        RECT 279.305 2597.840 279.595 2597.885 ;
        RECT 306.905 2597.840 307.195 2597.885 ;
        RECT 279.305 2597.700 307.195 2597.840 ;
        RECT 279.305 2597.655 279.595 2597.700 ;
        RECT 306.905 2597.655 307.195 2597.700 ;
        RECT 375.905 2597.840 376.195 2597.885 ;
        RECT 403.505 2597.840 403.795 2597.885 ;
        RECT 375.905 2597.700 403.795 2597.840 ;
        RECT 375.905 2597.655 376.195 2597.700 ;
        RECT 403.505 2597.655 403.795 2597.700 ;
        RECT 472.505 2597.840 472.795 2597.885 ;
        RECT 500.105 2597.840 500.395 2597.885 ;
        RECT 472.505 2597.700 500.395 2597.840 ;
        RECT 472.505 2597.655 472.795 2597.700 ;
        RECT 500.105 2597.655 500.395 2597.700 ;
        RECT 569.105 2597.840 569.395 2597.885 ;
        RECT 596.705 2597.840 596.995 2597.885 ;
        RECT 569.105 2597.700 596.995 2597.840 ;
        RECT 569.105 2597.655 569.395 2597.700 ;
        RECT 596.705 2597.655 596.995 2597.700 ;
        RECT 665.705 2597.840 665.995 2597.885 ;
        RECT 693.305 2597.840 693.595 2597.885 ;
        RECT 665.705 2597.700 693.595 2597.840 ;
        RECT 665.705 2597.655 665.995 2597.700 ;
        RECT 693.305 2597.655 693.595 2597.700 ;
        RECT 762.305 2597.840 762.595 2597.885 ;
        RECT 789.905 2597.840 790.195 2597.885 ;
        RECT 762.305 2597.700 790.195 2597.840 ;
        RECT 762.305 2597.655 762.595 2597.700 ;
        RECT 789.905 2597.655 790.195 2597.700 ;
        RECT 949.985 2597.840 950.275 2597.885 ;
        RECT 979.885 2597.840 980.175 2597.885 ;
        RECT 949.985 2597.700 980.175 2597.840 ;
        RECT 949.985 2597.655 950.275 2597.700 ;
        RECT 979.885 2597.655 980.175 2597.700 ;
        RECT 1628.485 2596.820 1628.775 2596.865 ;
        RECT 1698.390 2596.820 1698.710 2596.880 ;
        RECT 1628.485 2596.680 1698.710 2596.820 ;
        RECT 1628.485 2596.635 1628.775 2596.680 ;
        RECT 1698.390 2596.620 1698.710 2596.680 ;
        RECT 18.470 2596.140 18.790 2596.200 ;
        RECT 86.105 2596.140 86.395 2596.185 ;
        RECT 18.470 2596.000 86.395 2596.140 ;
        RECT 18.470 2595.940 18.790 2596.000 ;
        RECT 86.105 2595.955 86.395 2596.000 ;
        RECT 113.705 2596.140 113.995 2596.185 ;
        RECT 182.705 2596.140 182.995 2596.185 ;
        RECT 113.705 2596.000 182.995 2596.140 ;
        RECT 113.705 2595.955 113.995 2596.000 ;
        RECT 182.705 2595.955 182.995 2596.000 ;
        RECT 210.305 2596.140 210.595 2596.185 ;
        RECT 279.305 2596.140 279.595 2596.185 ;
        RECT 210.305 2596.000 279.595 2596.140 ;
        RECT 210.305 2595.955 210.595 2596.000 ;
        RECT 279.305 2595.955 279.595 2596.000 ;
        RECT 306.905 2596.140 307.195 2596.185 ;
        RECT 375.905 2596.140 376.195 2596.185 ;
        RECT 306.905 2596.000 376.195 2596.140 ;
        RECT 306.905 2595.955 307.195 2596.000 ;
        RECT 375.905 2595.955 376.195 2596.000 ;
        RECT 403.505 2596.140 403.795 2596.185 ;
        RECT 472.505 2596.140 472.795 2596.185 ;
        RECT 403.505 2596.000 472.795 2596.140 ;
        RECT 403.505 2595.955 403.795 2596.000 ;
        RECT 472.505 2595.955 472.795 2596.000 ;
        RECT 500.105 2596.140 500.395 2596.185 ;
        RECT 569.105 2596.140 569.395 2596.185 ;
        RECT 500.105 2596.000 569.395 2596.140 ;
        RECT 500.105 2595.955 500.395 2596.000 ;
        RECT 569.105 2595.955 569.395 2596.000 ;
        RECT 596.705 2596.140 596.995 2596.185 ;
        RECT 665.705 2596.140 665.995 2596.185 ;
        RECT 596.705 2596.000 665.995 2596.140 ;
        RECT 596.705 2595.955 596.995 2596.000 ;
        RECT 665.705 2595.955 665.995 2596.000 ;
        RECT 693.305 2596.140 693.595 2596.185 ;
        RECT 762.305 2596.140 762.595 2596.185 ;
        RECT 693.305 2596.000 762.595 2596.140 ;
        RECT 693.305 2595.955 693.595 2596.000 ;
        RECT 762.305 2595.955 762.595 2596.000 ;
        RECT 789.905 2596.140 790.195 2596.185 ;
        RECT 858.905 2596.140 859.195 2596.185 ;
        RECT 789.905 2596.000 859.195 2596.140 ;
        RECT 789.905 2595.955 790.195 2596.000 ;
        RECT 858.905 2595.955 859.195 2596.000 ;
        RECT 907.205 2596.140 907.495 2596.185 ;
        RECT 949.985 2596.140 950.275 2596.185 ;
        RECT 907.205 2596.000 950.275 2596.140 ;
        RECT 907.205 2595.955 907.495 2596.000 ;
        RECT 949.985 2595.955 950.275 2596.000 ;
        RECT 979.885 2596.140 980.175 2596.185 ;
        RECT 1048.885 2596.140 1049.175 2596.185 ;
        RECT 979.885 2596.000 1049.175 2596.140 ;
        RECT 979.885 2595.955 980.175 2596.000 ;
        RECT 1048.885 2595.955 1049.175 2596.000 ;
        RECT 1096.725 2596.140 1097.015 2596.185 ;
        RECT 1526.825 2596.140 1527.115 2596.185 ;
        RECT 1096.725 2596.000 1527.115 2596.140 ;
        RECT 1096.725 2595.955 1097.015 2596.000 ;
        RECT 1526.825 2595.955 1527.115 2596.000 ;
        RECT 1584.325 2596.140 1584.615 2596.185 ;
        RECT 1628.485 2596.140 1628.775 2596.185 ;
        RECT 1584.325 2596.000 1628.775 2596.140 ;
        RECT 1584.325 2595.955 1584.615 2596.000 ;
        RECT 1628.485 2595.955 1628.775 2596.000 ;
      LAYER via ;
        RECT 1698.420 2596.620 1698.680 2596.880 ;
        RECT 18.500 2595.940 18.760 2596.200 ;
      LAYER met2 ;
        RECT 1698.420 2596.650 1698.680 2596.910 ;
        RECT 1700.170 2596.650 1700.450 2600.000 ;
        RECT 1698.420 2596.590 1700.450 2596.650 ;
        RECT 1698.480 2596.510 1700.450 2596.590 ;
        RECT 18.500 2595.910 18.760 2596.230 ;
        RECT 1700.170 2596.000 1700.450 2596.510 ;
        RECT 18.560 1040.925 18.700 2595.910 ;
        RECT 18.490 1040.555 18.770 1040.925 ;
      LAYER via2 ;
        RECT 18.490 1040.600 18.770 1040.880 ;
      LAYER met3 ;
        RECT -4.000 1040.890 2.000 1041.340 ;
        RECT 18.465 1040.890 18.795 1040.905 ;
        RECT -4.000 1040.590 18.795 1040.890 ;
        RECT -4.000 1040.140 2.000 1040.590 ;
        RECT 18.465 1040.575 18.795 1040.590 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1534.245 2595.645 1535.335 2595.815 ;
      LAYER mcon ;
        RECT 1535.165 2595.645 1535.335 2595.815 ;
      LAYER met1 ;
        RECT 1725.070 2596.280 1725.390 2596.540 ;
        RECT 25.830 2595.800 26.150 2595.860 ;
        RECT 1534.185 2595.800 1534.475 2595.845 ;
        RECT 25.830 2595.660 1534.475 2595.800 ;
        RECT 25.830 2595.600 26.150 2595.660 ;
        RECT 1534.185 2595.615 1534.475 2595.660 ;
        RECT 1535.105 2595.800 1535.395 2595.845 ;
        RECT 1725.160 2595.800 1725.300 2596.280 ;
        RECT 1535.105 2595.660 1725.300 2595.800 ;
        RECT 1535.105 2595.615 1535.395 2595.660 ;
        RECT 13.870 827.460 14.190 827.520 ;
        RECT 25.830 827.460 26.150 827.520 ;
        RECT 13.870 827.320 26.150 827.460 ;
        RECT 13.870 827.260 14.190 827.320 ;
        RECT 25.830 827.260 26.150 827.320 ;
      LAYER via ;
        RECT 1725.100 2596.280 1725.360 2596.540 ;
        RECT 25.860 2595.600 26.120 2595.860 ;
        RECT 13.900 827.260 14.160 827.520 ;
        RECT 25.860 827.260 26.120 827.520 ;
      LAYER met2 ;
        RECT 1725.930 2596.650 1726.210 2600.000 ;
        RECT 1725.160 2596.570 1726.210 2596.650 ;
        RECT 1725.100 2596.510 1726.210 2596.570 ;
        RECT 1725.100 2596.250 1725.360 2596.510 ;
        RECT 1725.930 2596.000 1726.210 2596.510 ;
        RECT 25.860 2595.570 26.120 2595.890 ;
        RECT 25.920 827.550 26.060 2595.570 ;
        RECT 13.900 827.230 14.160 827.550 ;
        RECT 25.860 827.230 26.120 827.550 ;
        RECT 13.960 825.365 14.100 827.230 ;
        RECT 13.890 824.995 14.170 825.365 ;
      LAYER via2 ;
        RECT 13.890 825.040 14.170 825.320 ;
      LAYER met3 ;
        RECT -4.000 825.330 2.000 825.780 ;
        RECT 13.865 825.330 14.195 825.345 ;
        RECT -4.000 825.030 14.195 825.330 ;
        RECT -4.000 824.580 2.000 825.030 ;
        RECT 13.865 825.015 14.195 825.030 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 85.705 2595.305 85.875 2598.195 ;
        RECT 134.465 2595.305 134.635 2598.195 ;
        RECT 182.305 2595.305 182.475 2598.195 ;
        RECT 231.065 2595.305 231.235 2598.195 ;
        RECT 278.905 2595.305 279.075 2598.195 ;
        RECT 327.665 2595.305 327.835 2598.195 ;
        RECT 375.505 2595.305 375.675 2598.195 ;
        RECT 424.265 2595.305 424.435 2598.195 ;
        RECT 472.105 2595.305 472.275 2598.195 ;
        RECT 520.865 2595.305 521.035 2598.195 ;
        RECT 568.705 2595.305 568.875 2598.195 ;
        RECT 617.465 2595.305 617.635 2598.195 ;
        RECT 665.305 2595.305 665.475 2598.195 ;
        RECT 714.065 2595.305 714.235 2598.195 ;
        RECT 761.905 2595.305 762.075 2598.195 ;
        RECT 810.665 2595.305 810.835 2598.195 ;
        RECT 858.505 2595.305 858.675 2598.535 ;
        RECT 906.805 2595.305 906.975 2598.535 ;
        RECT 955.565 2595.305 955.735 2598.195 ;
        RECT 1003.865 2595.305 1004.035 2598.195 ;
        RECT 1049.405 2595.475 1049.575 2598.535 ;
        RECT 1048.945 2595.305 1049.575 2595.475 ;
        RECT 1096.325 2595.475 1096.495 2598.535 ;
        RECT 1096.325 2595.305 1096.955 2595.475 ;
        RECT 1583.925 2595.305 1584.095 2596.155 ;
        RECT 1629.005 2595.475 1629.175 2597.175 ;
        RECT 1628.545 2595.305 1629.175 2595.475 ;
        RECT 1676.385 2595.305 1676.555 2597.175 ;
        RECT 1749.985 2595.305 1750.155 2596.495 ;
      LAYER mcon ;
        RECT 858.505 2598.365 858.675 2598.535 ;
        RECT 85.705 2598.025 85.875 2598.195 ;
        RECT 134.465 2598.025 134.635 2598.195 ;
        RECT 182.305 2598.025 182.475 2598.195 ;
        RECT 231.065 2598.025 231.235 2598.195 ;
        RECT 278.905 2598.025 279.075 2598.195 ;
        RECT 327.665 2598.025 327.835 2598.195 ;
        RECT 375.505 2598.025 375.675 2598.195 ;
        RECT 424.265 2598.025 424.435 2598.195 ;
        RECT 472.105 2598.025 472.275 2598.195 ;
        RECT 520.865 2598.025 521.035 2598.195 ;
        RECT 568.705 2598.025 568.875 2598.195 ;
        RECT 617.465 2598.025 617.635 2598.195 ;
        RECT 665.305 2598.025 665.475 2598.195 ;
        RECT 714.065 2598.025 714.235 2598.195 ;
        RECT 761.905 2598.025 762.075 2598.195 ;
        RECT 810.665 2598.025 810.835 2598.195 ;
        RECT 906.805 2598.365 906.975 2598.535 ;
        RECT 1049.405 2598.365 1049.575 2598.535 ;
        RECT 955.565 2598.025 955.735 2598.195 ;
        RECT 1003.865 2598.025 1004.035 2598.195 ;
        RECT 1096.325 2598.365 1096.495 2598.535 ;
        RECT 1629.005 2597.005 1629.175 2597.175 ;
        RECT 1583.925 2595.985 1584.095 2596.155 ;
        RECT 1096.785 2595.305 1096.955 2595.475 ;
        RECT 1676.385 2597.005 1676.555 2597.175 ;
        RECT 1749.985 2596.325 1750.155 2596.495 ;
      LAYER met1 ;
        RECT 858.445 2598.520 858.735 2598.565 ;
        RECT 906.745 2598.520 907.035 2598.565 ;
        RECT 858.445 2598.380 907.035 2598.520 ;
        RECT 858.445 2598.335 858.735 2598.380 ;
        RECT 906.745 2598.335 907.035 2598.380 ;
        RECT 1049.345 2598.520 1049.635 2598.565 ;
        RECT 1096.265 2598.520 1096.555 2598.565 ;
        RECT 1049.345 2598.380 1096.555 2598.520 ;
        RECT 1049.345 2598.335 1049.635 2598.380 ;
        RECT 1096.265 2598.335 1096.555 2598.380 ;
        RECT 85.645 2598.180 85.935 2598.225 ;
        RECT 134.405 2598.180 134.695 2598.225 ;
        RECT 85.645 2598.040 134.695 2598.180 ;
        RECT 85.645 2597.995 85.935 2598.040 ;
        RECT 134.405 2597.995 134.695 2598.040 ;
        RECT 182.245 2598.180 182.535 2598.225 ;
        RECT 231.005 2598.180 231.295 2598.225 ;
        RECT 182.245 2598.040 231.295 2598.180 ;
        RECT 182.245 2597.995 182.535 2598.040 ;
        RECT 231.005 2597.995 231.295 2598.040 ;
        RECT 278.845 2598.180 279.135 2598.225 ;
        RECT 327.605 2598.180 327.895 2598.225 ;
        RECT 278.845 2598.040 327.895 2598.180 ;
        RECT 278.845 2597.995 279.135 2598.040 ;
        RECT 327.605 2597.995 327.895 2598.040 ;
        RECT 375.445 2598.180 375.735 2598.225 ;
        RECT 424.205 2598.180 424.495 2598.225 ;
        RECT 375.445 2598.040 424.495 2598.180 ;
        RECT 375.445 2597.995 375.735 2598.040 ;
        RECT 424.205 2597.995 424.495 2598.040 ;
        RECT 472.045 2598.180 472.335 2598.225 ;
        RECT 520.805 2598.180 521.095 2598.225 ;
        RECT 472.045 2598.040 521.095 2598.180 ;
        RECT 472.045 2597.995 472.335 2598.040 ;
        RECT 520.805 2597.995 521.095 2598.040 ;
        RECT 568.645 2598.180 568.935 2598.225 ;
        RECT 617.405 2598.180 617.695 2598.225 ;
        RECT 568.645 2598.040 617.695 2598.180 ;
        RECT 568.645 2597.995 568.935 2598.040 ;
        RECT 617.405 2597.995 617.695 2598.040 ;
        RECT 665.245 2598.180 665.535 2598.225 ;
        RECT 714.005 2598.180 714.295 2598.225 ;
        RECT 665.245 2598.040 714.295 2598.180 ;
        RECT 665.245 2597.995 665.535 2598.040 ;
        RECT 714.005 2597.995 714.295 2598.040 ;
        RECT 761.845 2598.180 762.135 2598.225 ;
        RECT 810.605 2598.180 810.895 2598.225 ;
        RECT 761.845 2598.040 810.895 2598.180 ;
        RECT 761.845 2597.995 762.135 2598.040 ;
        RECT 810.605 2597.995 810.895 2598.040 ;
        RECT 955.505 2598.180 955.795 2598.225 ;
        RECT 1003.805 2598.180 1004.095 2598.225 ;
        RECT 955.505 2598.040 1004.095 2598.180 ;
        RECT 955.505 2597.995 955.795 2598.040 ;
        RECT 1003.805 2597.995 1004.095 2598.040 ;
        RECT 1628.945 2597.160 1629.235 2597.205 ;
        RECT 1676.325 2597.160 1676.615 2597.205 ;
        RECT 1628.945 2597.020 1676.615 2597.160 ;
        RECT 1628.945 2596.975 1629.235 2597.020 ;
        RECT 1676.325 2596.975 1676.615 2597.020 ;
        RECT 1749.910 2596.480 1750.230 2596.540 ;
        RECT 1749.715 2596.340 1750.230 2596.480 ;
        RECT 1749.910 2596.280 1750.230 2596.340 ;
        RECT 1583.865 2596.140 1584.155 2596.185 ;
        RECT 1534.720 2596.000 1584.155 2596.140 ;
        RECT 24.910 2595.460 25.230 2595.520 ;
        RECT 85.645 2595.460 85.935 2595.505 ;
        RECT 24.910 2595.320 85.935 2595.460 ;
        RECT 24.910 2595.260 25.230 2595.320 ;
        RECT 85.645 2595.275 85.935 2595.320 ;
        RECT 134.405 2595.460 134.695 2595.505 ;
        RECT 182.245 2595.460 182.535 2595.505 ;
        RECT 134.405 2595.320 182.535 2595.460 ;
        RECT 134.405 2595.275 134.695 2595.320 ;
        RECT 182.245 2595.275 182.535 2595.320 ;
        RECT 231.005 2595.460 231.295 2595.505 ;
        RECT 278.845 2595.460 279.135 2595.505 ;
        RECT 231.005 2595.320 279.135 2595.460 ;
        RECT 231.005 2595.275 231.295 2595.320 ;
        RECT 278.845 2595.275 279.135 2595.320 ;
        RECT 327.605 2595.460 327.895 2595.505 ;
        RECT 375.445 2595.460 375.735 2595.505 ;
        RECT 327.605 2595.320 375.735 2595.460 ;
        RECT 327.605 2595.275 327.895 2595.320 ;
        RECT 375.445 2595.275 375.735 2595.320 ;
        RECT 424.205 2595.460 424.495 2595.505 ;
        RECT 472.045 2595.460 472.335 2595.505 ;
        RECT 424.205 2595.320 472.335 2595.460 ;
        RECT 424.205 2595.275 424.495 2595.320 ;
        RECT 472.045 2595.275 472.335 2595.320 ;
        RECT 520.805 2595.460 521.095 2595.505 ;
        RECT 568.645 2595.460 568.935 2595.505 ;
        RECT 520.805 2595.320 568.935 2595.460 ;
        RECT 520.805 2595.275 521.095 2595.320 ;
        RECT 568.645 2595.275 568.935 2595.320 ;
        RECT 617.405 2595.460 617.695 2595.505 ;
        RECT 665.245 2595.460 665.535 2595.505 ;
        RECT 617.405 2595.320 665.535 2595.460 ;
        RECT 617.405 2595.275 617.695 2595.320 ;
        RECT 665.245 2595.275 665.535 2595.320 ;
        RECT 714.005 2595.460 714.295 2595.505 ;
        RECT 761.845 2595.460 762.135 2595.505 ;
        RECT 714.005 2595.320 762.135 2595.460 ;
        RECT 714.005 2595.275 714.295 2595.320 ;
        RECT 761.845 2595.275 762.135 2595.320 ;
        RECT 810.605 2595.460 810.895 2595.505 ;
        RECT 858.445 2595.460 858.735 2595.505 ;
        RECT 810.605 2595.320 858.735 2595.460 ;
        RECT 810.605 2595.275 810.895 2595.320 ;
        RECT 858.445 2595.275 858.735 2595.320 ;
        RECT 906.745 2595.460 907.035 2595.505 ;
        RECT 955.505 2595.460 955.795 2595.505 ;
        RECT 906.745 2595.320 955.795 2595.460 ;
        RECT 906.745 2595.275 907.035 2595.320 ;
        RECT 955.505 2595.275 955.795 2595.320 ;
        RECT 1003.805 2595.460 1004.095 2595.505 ;
        RECT 1048.885 2595.460 1049.175 2595.505 ;
        RECT 1003.805 2595.320 1049.175 2595.460 ;
        RECT 1003.805 2595.275 1004.095 2595.320 ;
        RECT 1048.885 2595.275 1049.175 2595.320 ;
        RECT 1096.725 2595.460 1097.015 2595.505 ;
        RECT 1534.720 2595.460 1534.860 2596.000 ;
        RECT 1583.865 2595.955 1584.155 2596.000 ;
        RECT 1096.725 2595.320 1534.860 2595.460 ;
        RECT 1583.865 2595.460 1584.155 2595.505 ;
        RECT 1628.485 2595.460 1628.775 2595.505 ;
        RECT 1583.865 2595.320 1628.775 2595.460 ;
        RECT 1096.725 2595.275 1097.015 2595.320 ;
        RECT 1583.865 2595.275 1584.155 2595.320 ;
        RECT 1628.485 2595.275 1628.775 2595.320 ;
        RECT 1676.325 2595.460 1676.615 2595.505 ;
        RECT 1749.925 2595.460 1750.215 2595.505 ;
        RECT 1676.325 2595.320 1750.215 2595.460 ;
        RECT 1676.325 2595.275 1676.615 2595.320 ;
        RECT 1749.925 2595.275 1750.215 2595.320 ;
        RECT 13.870 611.560 14.190 611.620 ;
        RECT 24.910 611.560 25.230 611.620 ;
        RECT 13.870 611.420 25.230 611.560 ;
        RECT 13.870 611.360 14.190 611.420 ;
        RECT 24.910 611.360 25.230 611.420 ;
      LAYER via ;
        RECT 1749.940 2596.280 1750.200 2596.540 ;
        RECT 24.940 2595.260 25.200 2595.520 ;
        RECT 13.900 611.360 14.160 611.620 ;
        RECT 24.940 611.360 25.200 611.620 ;
      LAYER met2 ;
        RECT 1751.690 2596.650 1751.970 2600.000 ;
        RECT 1750.000 2596.570 1751.970 2596.650 ;
        RECT 1749.940 2596.510 1751.970 2596.570 ;
        RECT 1749.940 2596.250 1750.200 2596.510 ;
        RECT 1751.690 2596.000 1751.970 2596.510 ;
        RECT 24.940 2595.230 25.200 2595.550 ;
        RECT 25.000 611.650 25.140 2595.230 ;
        RECT 13.900 611.330 14.160 611.650 ;
        RECT 24.940 611.330 25.200 611.650 ;
        RECT 13.960 610.485 14.100 611.330 ;
        RECT 13.890 610.115 14.170 610.485 ;
      LAYER via2 ;
        RECT 13.890 610.160 14.170 610.440 ;
      LAYER met3 ;
        RECT -4.000 610.450 2.000 610.900 ;
        RECT 13.865 610.450 14.195 610.465 ;
        RECT -4.000 610.150 14.195 610.450 ;
        RECT -4.000 609.700 2.000 610.150 ;
        RECT 13.865 610.135 14.195 610.150 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1775.745 2594.965 1775.915 2596.495 ;
      LAYER mcon ;
        RECT 1775.745 2596.325 1775.915 2596.495 ;
      LAYER met1 ;
        RECT 1775.670 2596.480 1775.990 2596.540 ;
        RECT 1775.475 2596.340 1775.990 2596.480 ;
        RECT 1775.670 2596.280 1775.990 2596.340 ;
        RECT 17.090 2595.120 17.410 2595.180 ;
        RECT 1775.685 2595.120 1775.975 2595.165 ;
        RECT 17.090 2594.980 1534.860 2595.120 ;
        RECT 17.090 2594.920 17.410 2594.980 ;
        RECT 1534.720 2594.440 1534.860 2594.980 ;
        RECT 1559.560 2594.980 1775.975 2595.120 ;
        RECT 1559.560 2594.780 1559.700 2594.980 ;
        RECT 1775.685 2594.935 1775.975 2594.980 ;
        RECT 1535.640 2594.640 1559.700 2594.780 ;
        RECT 1535.640 2594.440 1535.780 2594.640 ;
        RECT 1534.720 2594.300 1535.780 2594.440 ;
      LAYER via ;
        RECT 1775.700 2596.280 1775.960 2596.540 ;
        RECT 17.120 2594.920 17.380 2595.180 ;
      LAYER met2 ;
        RECT 1776.990 2596.650 1777.270 2600.000 ;
        RECT 1775.760 2596.570 1777.270 2596.650 ;
        RECT 1775.700 2596.510 1777.270 2596.570 ;
        RECT 1775.700 2596.250 1775.960 2596.510 ;
        RECT 1776.990 2596.000 1777.270 2596.510 ;
        RECT 17.120 2594.890 17.380 2595.210 ;
        RECT 17.180 394.925 17.320 2594.890 ;
        RECT 17.110 394.555 17.390 394.925 ;
      LAYER via2 ;
        RECT 17.110 394.600 17.390 394.880 ;
      LAYER met3 ;
        RECT -4.000 394.890 2.000 395.340 ;
        RECT 17.085 394.890 17.415 394.905 ;
        RECT -4.000 394.590 17.415 394.890 ;
        RECT -4.000 394.140 2.000 394.590 ;
        RECT 17.085 394.575 17.415 394.590 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 86.625 2594.625 86.795 2598.535 ;
        RECT 134.005 2594.625 134.175 2598.535 ;
        RECT 183.225 2594.625 183.395 2598.535 ;
        RECT 230.605 2594.625 230.775 2598.535 ;
        RECT 279.825 2594.625 279.995 2598.535 ;
        RECT 327.205 2594.625 327.375 2598.535 ;
        RECT 376.425 2594.625 376.595 2598.535 ;
        RECT 423.805 2594.625 423.975 2598.535 ;
        RECT 473.025 2594.625 473.195 2598.535 ;
        RECT 520.405 2594.625 520.575 2598.535 ;
        RECT 569.625 2594.625 569.795 2598.535 ;
        RECT 617.005 2594.625 617.175 2598.535 ;
        RECT 666.225 2594.625 666.395 2598.535 ;
        RECT 713.605 2594.625 713.775 2598.535 ;
        RECT 762.825 2594.625 762.995 2598.535 ;
        RECT 810.205 2594.625 810.375 2598.535 ;
        RECT 859.425 2594.625 859.595 2598.875 ;
        RECT 907.725 2594.625 907.895 2598.875 ;
        RECT 941.765 2594.625 941.935 2598.535 ;
        RECT 1003.405 2594.625 1003.575 2598.535 ;
        RECT 1049.865 2594.795 1050.035 2598.875 ;
        RECT 1048.945 2594.625 1050.035 2594.795 ;
        RECT 1095.865 2594.795 1096.035 2598.875 ;
        RECT 1534.245 2595.305 1535.795 2595.475 ;
        RECT 1095.865 2594.625 1096.955 2594.795 ;
        RECT 1534.245 2594.625 1534.415 2595.305 ;
        RECT 1583.465 2594.625 1583.635 2595.475 ;
        RECT 1629.465 2594.795 1629.635 2597.515 ;
        RECT 1628.545 2594.625 1629.635 2594.795 ;
        RECT 1675.925 2594.795 1676.095 2597.515 ;
        RECT 1725.605 2594.795 1725.775 2595.815 ;
        RECT 1675.925 2594.625 1676.555 2594.795 ;
        RECT 1725.145 2594.625 1725.775 2594.795 ;
      LAYER mcon ;
        RECT 859.425 2598.705 859.595 2598.875 ;
        RECT 86.625 2598.365 86.795 2598.535 ;
        RECT 134.005 2598.365 134.175 2598.535 ;
        RECT 183.225 2598.365 183.395 2598.535 ;
        RECT 230.605 2598.365 230.775 2598.535 ;
        RECT 279.825 2598.365 279.995 2598.535 ;
        RECT 327.205 2598.365 327.375 2598.535 ;
        RECT 376.425 2598.365 376.595 2598.535 ;
        RECT 423.805 2598.365 423.975 2598.535 ;
        RECT 473.025 2598.365 473.195 2598.535 ;
        RECT 520.405 2598.365 520.575 2598.535 ;
        RECT 569.625 2598.365 569.795 2598.535 ;
        RECT 617.005 2598.365 617.175 2598.535 ;
        RECT 666.225 2598.365 666.395 2598.535 ;
        RECT 713.605 2598.365 713.775 2598.535 ;
        RECT 762.825 2598.365 762.995 2598.535 ;
        RECT 810.205 2598.365 810.375 2598.535 ;
        RECT 907.725 2598.705 907.895 2598.875 ;
        RECT 1049.865 2598.705 1050.035 2598.875 ;
        RECT 941.765 2598.365 941.935 2598.535 ;
        RECT 1003.405 2598.365 1003.575 2598.535 ;
        RECT 1095.865 2598.705 1096.035 2598.875 ;
        RECT 1629.465 2597.345 1629.635 2597.515 ;
        RECT 1535.625 2595.305 1535.795 2595.475 ;
        RECT 1583.465 2595.305 1583.635 2595.475 ;
        RECT 1096.785 2594.625 1096.955 2594.795 ;
        RECT 1675.925 2597.345 1676.095 2597.515 ;
        RECT 1725.605 2595.645 1725.775 2595.815 ;
        RECT 1676.385 2594.625 1676.555 2594.795 ;
      LAYER met1 ;
        RECT 859.365 2598.860 859.655 2598.905 ;
        RECT 907.665 2598.860 907.955 2598.905 ;
        RECT 859.365 2598.720 907.955 2598.860 ;
        RECT 859.365 2598.675 859.655 2598.720 ;
        RECT 907.665 2598.675 907.955 2598.720 ;
        RECT 1049.805 2598.860 1050.095 2598.905 ;
        RECT 1095.805 2598.860 1096.095 2598.905 ;
        RECT 1049.805 2598.720 1096.095 2598.860 ;
        RECT 1049.805 2598.675 1050.095 2598.720 ;
        RECT 1095.805 2598.675 1096.095 2598.720 ;
        RECT 86.565 2598.520 86.855 2598.565 ;
        RECT 133.945 2598.520 134.235 2598.565 ;
        RECT 86.565 2598.380 134.235 2598.520 ;
        RECT 86.565 2598.335 86.855 2598.380 ;
        RECT 133.945 2598.335 134.235 2598.380 ;
        RECT 183.165 2598.520 183.455 2598.565 ;
        RECT 230.545 2598.520 230.835 2598.565 ;
        RECT 183.165 2598.380 230.835 2598.520 ;
        RECT 183.165 2598.335 183.455 2598.380 ;
        RECT 230.545 2598.335 230.835 2598.380 ;
        RECT 279.765 2598.520 280.055 2598.565 ;
        RECT 327.145 2598.520 327.435 2598.565 ;
        RECT 279.765 2598.380 327.435 2598.520 ;
        RECT 279.765 2598.335 280.055 2598.380 ;
        RECT 327.145 2598.335 327.435 2598.380 ;
        RECT 376.365 2598.520 376.655 2598.565 ;
        RECT 423.745 2598.520 424.035 2598.565 ;
        RECT 376.365 2598.380 424.035 2598.520 ;
        RECT 376.365 2598.335 376.655 2598.380 ;
        RECT 423.745 2598.335 424.035 2598.380 ;
        RECT 472.965 2598.520 473.255 2598.565 ;
        RECT 520.345 2598.520 520.635 2598.565 ;
        RECT 472.965 2598.380 520.635 2598.520 ;
        RECT 472.965 2598.335 473.255 2598.380 ;
        RECT 520.345 2598.335 520.635 2598.380 ;
        RECT 569.565 2598.520 569.855 2598.565 ;
        RECT 616.945 2598.520 617.235 2598.565 ;
        RECT 569.565 2598.380 617.235 2598.520 ;
        RECT 569.565 2598.335 569.855 2598.380 ;
        RECT 616.945 2598.335 617.235 2598.380 ;
        RECT 666.165 2598.520 666.455 2598.565 ;
        RECT 713.545 2598.520 713.835 2598.565 ;
        RECT 666.165 2598.380 713.835 2598.520 ;
        RECT 666.165 2598.335 666.455 2598.380 ;
        RECT 713.545 2598.335 713.835 2598.380 ;
        RECT 762.765 2598.520 763.055 2598.565 ;
        RECT 810.145 2598.520 810.435 2598.565 ;
        RECT 762.765 2598.380 810.435 2598.520 ;
        RECT 762.765 2598.335 763.055 2598.380 ;
        RECT 810.145 2598.335 810.435 2598.380 ;
        RECT 941.705 2598.520 941.995 2598.565 ;
        RECT 1003.345 2598.520 1003.635 2598.565 ;
        RECT 941.705 2598.380 1003.635 2598.520 ;
        RECT 941.705 2598.335 941.995 2598.380 ;
        RECT 1003.345 2598.335 1003.635 2598.380 ;
        RECT 1629.405 2597.500 1629.695 2597.545 ;
        RECT 1675.865 2597.500 1676.155 2597.545 ;
        RECT 1629.405 2597.360 1676.155 2597.500 ;
        RECT 1629.405 2597.315 1629.695 2597.360 ;
        RECT 1675.865 2597.315 1676.155 2597.360 ;
        RECT 1801.430 2596.480 1801.750 2596.540 ;
        RECT 1776.220 2596.340 1801.750 2596.480 ;
        RECT 1725.545 2595.800 1725.835 2595.845 ;
        RECT 1776.220 2595.800 1776.360 2596.340 ;
        RECT 1801.430 2596.280 1801.750 2596.340 ;
        RECT 1725.545 2595.660 1776.360 2595.800 ;
        RECT 1725.545 2595.615 1725.835 2595.660 ;
        RECT 1535.565 2595.460 1535.855 2595.505 ;
        RECT 1583.405 2595.460 1583.695 2595.505 ;
        RECT 1535.565 2595.320 1583.695 2595.460 ;
        RECT 1535.565 2595.275 1535.855 2595.320 ;
        RECT 1583.405 2595.275 1583.695 2595.320 ;
        RECT 23.990 2594.780 24.310 2594.840 ;
        RECT 86.565 2594.780 86.855 2594.825 ;
        RECT 23.990 2594.640 86.855 2594.780 ;
        RECT 23.990 2594.580 24.310 2594.640 ;
        RECT 86.565 2594.595 86.855 2594.640 ;
        RECT 133.945 2594.780 134.235 2594.825 ;
        RECT 183.165 2594.780 183.455 2594.825 ;
        RECT 133.945 2594.640 183.455 2594.780 ;
        RECT 133.945 2594.595 134.235 2594.640 ;
        RECT 183.165 2594.595 183.455 2594.640 ;
        RECT 230.545 2594.780 230.835 2594.825 ;
        RECT 279.765 2594.780 280.055 2594.825 ;
        RECT 230.545 2594.640 280.055 2594.780 ;
        RECT 230.545 2594.595 230.835 2594.640 ;
        RECT 279.765 2594.595 280.055 2594.640 ;
        RECT 327.145 2594.780 327.435 2594.825 ;
        RECT 376.365 2594.780 376.655 2594.825 ;
        RECT 327.145 2594.640 376.655 2594.780 ;
        RECT 327.145 2594.595 327.435 2594.640 ;
        RECT 376.365 2594.595 376.655 2594.640 ;
        RECT 423.745 2594.780 424.035 2594.825 ;
        RECT 472.965 2594.780 473.255 2594.825 ;
        RECT 423.745 2594.640 473.255 2594.780 ;
        RECT 423.745 2594.595 424.035 2594.640 ;
        RECT 472.965 2594.595 473.255 2594.640 ;
        RECT 520.345 2594.780 520.635 2594.825 ;
        RECT 569.565 2594.780 569.855 2594.825 ;
        RECT 520.345 2594.640 569.855 2594.780 ;
        RECT 520.345 2594.595 520.635 2594.640 ;
        RECT 569.565 2594.595 569.855 2594.640 ;
        RECT 616.945 2594.780 617.235 2594.825 ;
        RECT 666.165 2594.780 666.455 2594.825 ;
        RECT 616.945 2594.640 666.455 2594.780 ;
        RECT 616.945 2594.595 617.235 2594.640 ;
        RECT 666.165 2594.595 666.455 2594.640 ;
        RECT 713.545 2594.780 713.835 2594.825 ;
        RECT 762.765 2594.780 763.055 2594.825 ;
        RECT 713.545 2594.640 763.055 2594.780 ;
        RECT 713.545 2594.595 713.835 2594.640 ;
        RECT 762.765 2594.595 763.055 2594.640 ;
        RECT 810.145 2594.780 810.435 2594.825 ;
        RECT 859.365 2594.780 859.655 2594.825 ;
        RECT 810.145 2594.640 859.655 2594.780 ;
        RECT 810.145 2594.595 810.435 2594.640 ;
        RECT 859.365 2594.595 859.655 2594.640 ;
        RECT 907.665 2594.780 907.955 2594.825 ;
        RECT 941.705 2594.780 941.995 2594.825 ;
        RECT 907.665 2594.640 941.995 2594.780 ;
        RECT 907.665 2594.595 907.955 2594.640 ;
        RECT 941.705 2594.595 941.995 2594.640 ;
        RECT 1003.345 2594.780 1003.635 2594.825 ;
        RECT 1048.885 2594.780 1049.175 2594.825 ;
        RECT 1003.345 2594.640 1049.175 2594.780 ;
        RECT 1003.345 2594.595 1003.635 2594.640 ;
        RECT 1048.885 2594.595 1049.175 2594.640 ;
        RECT 1096.725 2594.780 1097.015 2594.825 ;
        RECT 1534.185 2594.780 1534.475 2594.825 ;
        RECT 1096.725 2594.640 1534.475 2594.780 ;
        RECT 1096.725 2594.595 1097.015 2594.640 ;
        RECT 1534.185 2594.595 1534.475 2594.640 ;
        RECT 1583.405 2594.780 1583.695 2594.825 ;
        RECT 1628.485 2594.780 1628.775 2594.825 ;
        RECT 1583.405 2594.640 1628.775 2594.780 ;
        RECT 1583.405 2594.595 1583.695 2594.640 ;
        RECT 1628.485 2594.595 1628.775 2594.640 ;
        RECT 1676.325 2594.780 1676.615 2594.825 ;
        RECT 1725.085 2594.780 1725.375 2594.825 ;
        RECT 1676.325 2594.640 1725.375 2594.780 ;
        RECT 1676.325 2594.595 1676.615 2594.640 ;
        RECT 1725.085 2594.595 1725.375 2594.640 ;
        RECT 13.870 179.420 14.190 179.480 ;
        RECT 23.990 179.420 24.310 179.480 ;
        RECT 13.870 179.280 24.310 179.420 ;
        RECT 13.870 179.220 14.190 179.280 ;
        RECT 23.990 179.220 24.310 179.280 ;
      LAYER via ;
        RECT 1801.460 2596.280 1801.720 2596.540 ;
        RECT 24.020 2594.580 24.280 2594.840 ;
        RECT 13.900 179.220 14.160 179.480 ;
        RECT 24.020 179.220 24.280 179.480 ;
      LAYER met2 ;
        RECT 1802.750 2596.650 1803.030 2600.000 ;
        RECT 1801.520 2596.570 1803.030 2596.650 ;
        RECT 1801.460 2596.510 1803.030 2596.570 ;
        RECT 1801.460 2596.250 1801.720 2596.510 ;
        RECT 1802.750 2596.000 1803.030 2596.510 ;
        RECT 24.020 2594.550 24.280 2594.870 ;
        RECT 24.080 179.510 24.220 2594.550 ;
        RECT 13.900 179.365 14.160 179.510 ;
        RECT 13.890 178.995 14.170 179.365 ;
        RECT 24.020 179.190 24.280 179.510 ;
      LAYER via2 ;
        RECT 13.890 179.040 14.170 179.320 ;
      LAYER met3 ;
        RECT -4.000 179.330 2.000 179.780 ;
        RECT 13.865 179.330 14.195 179.345 ;
        RECT -4.000 179.030 14.195 179.330 ;
        RECT -4.000 178.580 2.000 179.030 ;
        RECT 13.865 179.015 14.195 179.030 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1381.065 2608.225 1382.615 2608.395 ;
        RECT 1435.345 2608.225 1436.895 2608.395 ;
      LAYER mcon ;
        RECT 1382.445 2608.225 1382.615 2608.395 ;
        RECT 1436.725 2608.225 1436.895 2608.395 ;
      LAYER met1 ;
        RECT 930.650 2608.380 930.970 2608.440 ;
        RECT 1381.005 2608.380 1381.295 2608.425 ;
        RECT 930.650 2608.240 1381.295 2608.380 ;
        RECT 930.650 2608.180 930.970 2608.240 ;
        RECT 1381.005 2608.195 1381.295 2608.240 ;
        RECT 1382.385 2608.380 1382.675 2608.425 ;
        RECT 1435.285 2608.380 1435.575 2608.425 ;
        RECT 1382.385 2608.240 1435.575 2608.380 ;
        RECT 1382.385 2608.195 1382.675 2608.240 ;
        RECT 1435.285 2608.195 1435.575 2608.240 ;
        RECT 1436.665 2608.380 1436.955 2608.425 ;
        RECT 2903.590 2608.380 2903.910 2608.440 ;
        RECT 1436.665 2608.240 2903.910 2608.380 ;
        RECT 1436.665 2608.195 1436.955 2608.240 ;
        RECT 2903.590 2608.180 2903.910 2608.240 ;
      LAYER via ;
        RECT 930.680 2608.180 930.940 2608.440 ;
        RECT 2903.620 2608.180 2903.880 2608.440 ;
      LAYER met2 ;
        RECT 930.680 2608.150 930.940 2608.470 ;
        RECT 2903.620 2608.150 2903.880 2608.470 ;
        RECT 930.740 2600.050 930.880 2608.150 ;
        RECT 930.740 2600.000 931.270 2600.050 ;
        RECT 930.740 2599.910 931.330 2600.000 ;
        RECT 931.050 2596.000 931.330 2599.910 ;
        RECT 2903.680 792.045 2903.820 2608.150 ;
        RECT 2903.610 791.675 2903.890 792.045 ;
      LAYER via2 ;
        RECT 2903.610 791.720 2903.890 792.000 ;
      LAYER met3 ;
        RECT 2903.585 792.010 2903.915 792.025 ;
        RECT 2918.000 792.010 2924.000 792.460 ;
        RECT 2903.585 791.710 2924.000 792.010 ;
        RECT 2903.585 791.695 2903.915 791.710 ;
        RECT 2918.000 791.260 2924.000 791.710 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 958.270 2601.155 958.550 2601.525 ;
        RECT 956.350 2599.370 956.630 2600.000 ;
        RECT 958.340 2599.370 958.480 2601.155 ;
        RECT 956.350 2599.230 958.480 2599.370 ;
        RECT 956.350 2596.000 956.630 2599.230 ;
        RECT 2884.290 1026.955 2884.570 1027.325 ;
        RECT 2916.950 1026.955 2917.230 1027.325 ;
        RECT 2884.360 1021.885 2884.500 1026.955 ;
        RECT 2917.020 1026.645 2917.160 1026.955 ;
        RECT 2916.950 1026.275 2917.230 1026.645 ;
        RECT 2884.290 1021.515 2884.570 1021.885 ;
      LAYER via2 ;
        RECT 958.270 2601.200 958.550 2601.480 ;
        RECT 2884.290 1027.000 2884.570 1027.280 ;
        RECT 2916.950 1027.000 2917.230 1027.280 ;
        RECT 2916.950 1026.320 2917.230 1026.600 ;
        RECT 2884.290 1021.560 2884.570 1021.840 ;
      LAYER met3 ;
        RECT 958.245 2601.490 958.575 2601.505 ;
        RECT 1831.070 2601.490 1831.450 2601.500 ;
        RECT 958.245 2601.190 1831.450 2601.490 ;
        RECT 958.245 2601.175 958.575 2601.190 ;
        RECT 1831.070 2601.180 1831.450 2601.190 ;
        RECT 2884.265 1027.290 2884.595 1027.305 ;
        RECT 2916.925 1027.290 2917.255 1027.305 ;
        RECT 2884.265 1026.990 2917.255 1027.290 ;
        RECT 2884.265 1026.975 2884.595 1026.990 ;
        RECT 2916.925 1026.975 2917.255 1026.990 ;
        RECT 2916.925 1026.610 2917.255 1026.625 ;
        RECT 2918.000 1026.610 2924.000 1027.060 ;
        RECT 2916.925 1026.310 2924.000 1026.610 ;
        RECT 2916.925 1026.295 2917.255 1026.310 ;
        RECT 2918.000 1025.860 2924.000 1026.310 ;
        RECT 1831.070 1023.210 1831.450 1023.220 ;
        RECT 1831.070 1022.910 1870.050 1023.210 ;
        RECT 1831.070 1022.900 1831.450 1022.910 ;
        RECT 1869.750 1022.530 1870.050 1022.910 ;
        RECT 1918.510 1022.910 1966.650 1023.210 ;
        RECT 1869.750 1022.230 1917.890 1022.530 ;
        RECT 1917.590 1021.850 1917.890 1022.230 ;
        RECT 1918.510 1021.850 1918.810 1022.910 ;
        RECT 1966.350 1022.530 1966.650 1022.910 ;
        RECT 2015.110 1022.910 2063.250 1023.210 ;
        RECT 1966.350 1022.230 2014.490 1022.530 ;
        RECT 1917.590 1021.550 1918.810 1021.850 ;
        RECT 2014.190 1021.850 2014.490 1022.230 ;
        RECT 2015.110 1021.850 2015.410 1022.910 ;
        RECT 2062.950 1022.530 2063.250 1022.910 ;
        RECT 2111.710 1022.910 2159.850 1023.210 ;
        RECT 2062.950 1022.230 2111.090 1022.530 ;
        RECT 2014.190 1021.550 2015.410 1021.850 ;
        RECT 2110.790 1021.850 2111.090 1022.230 ;
        RECT 2111.710 1021.850 2112.010 1022.910 ;
        RECT 2159.550 1022.530 2159.850 1022.910 ;
        RECT 2208.310 1022.910 2256.450 1023.210 ;
        RECT 2159.550 1022.230 2207.690 1022.530 ;
        RECT 2110.790 1021.550 2112.010 1021.850 ;
        RECT 2207.390 1021.850 2207.690 1022.230 ;
        RECT 2208.310 1021.850 2208.610 1022.910 ;
        RECT 2256.150 1022.530 2256.450 1022.910 ;
        RECT 2304.910 1022.910 2353.050 1023.210 ;
        RECT 2256.150 1022.230 2304.290 1022.530 ;
        RECT 2207.390 1021.550 2208.610 1021.850 ;
        RECT 2303.990 1021.850 2304.290 1022.230 ;
        RECT 2304.910 1021.850 2305.210 1022.910 ;
        RECT 2352.750 1022.530 2353.050 1022.910 ;
        RECT 2401.510 1022.910 2449.650 1023.210 ;
        RECT 2352.750 1022.230 2400.890 1022.530 ;
        RECT 2303.990 1021.550 2305.210 1021.850 ;
        RECT 2400.590 1021.850 2400.890 1022.230 ;
        RECT 2401.510 1021.850 2401.810 1022.910 ;
        RECT 2449.350 1022.530 2449.650 1022.910 ;
        RECT 2498.110 1022.910 2546.250 1023.210 ;
        RECT 2449.350 1022.230 2497.490 1022.530 ;
        RECT 2400.590 1021.550 2401.810 1021.850 ;
        RECT 2497.190 1021.850 2497.490 1022.230 ;
        RECT 2498.110 1021.850 2498.410 1022.910 ;
        RECT 2545.950 1022.530 2546.250 1022.910 ;
        RECT 2594.710 1022.910 2642.850 1023.210 ;
        RECT 2545.950 1022.230 2594.090 1022.530 ;
        RECT 2497.190 1021.550 2498.410 1021.850 ;
        RECT 2593.790 1021.850 2594.090 1022.230 ;
        RECT 2594.710 1021.850 2595.010 1022.910 ;
        RECT 2642.550 1022.530 2642.850 1022.910 ;
        RECT 2691.310 1022.910 2739.450 1023.210 ;
        RECT 2642.550 1022.230 2690.690 1022.530 ;
        RECT 2593.790 1021.550 2595.010 1021.850 ;
        RECT 2690.390 1021.850 2690.690 1022.230 ;
        RECT 2691.310 1021.850 2691.610 1022.910 ;
        RECT 2739.150 1022.530 2739.450 1022.910 ;
        RECT 2787.910 1022.910 2836.050 1023.210 ;
        RECT 2739.150 1022.230 2787.290 1022.530 ;
        RECT 2690.390 1021.550 2691.610 1021.850 ;
        RECT 2786.990 1021.850 2787.290 1022.230 ;
        RECT 2787.910 1021.850 2788.210 1022.910 ;
        RECT 2835.750 1022.530 2836.050 1022.910 ;
        RECT 2835.750 1022.230 2883.890 1022.530 ;
        RECT 2786.990 1021.550 2788.210 1021.850 ;
        RECT 2883.590 1021.850 2883.890 1022.230 ;
        RECT 2884.265 1021.850 2884.595 1021.865 ;
        RECT 2883.590 1021.550 2884.595 1021.850 ;
        RECT 2884.265 1021.535 2884.595 1021.550 ;
      LAYER via3 ;
        RECT 1831.100 2601.180 1831.420 2601.500 ;
        RECT 1831.100 1022.900 1831.420 1023.220 ;
      LAYER met4 ;
        RECT 1831.095 2601.175 1831.425 2601.505 ;
        RECT 1831.110 1023.225 1831.410 2601.175 ;
        RECT 1831.095 1022.895 1831.425 1023.225 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 984.030 2614.755 984.310 2615.125 ;
        RECT 1048.430 2614.755 1048.710 2615.125 ;
        RECT 982.110 2599.370 982.390 2600.000 ;
        RECT 984.100 2599.370 984.240 2614.755 ;
        RECT 1048.500 2613.765 1048.640 2614.755 ;
        RECT 1048.430 2613.395 1048.710 2613.765 ;
        RECT 982.110 2599.230 984.240 2599.370 ;
        RECT 982.110 2596.000 982.390 2599.230 ;
        RECT 2884.290 1261.555 2884.570 1261.925 ;
        RECT 2916.950 1261.555 2917.230 1261.925 ;
        RECT 2884.360 1256.485 2884.500 1261.555 ;
        RECT 2917.020 1261.245 2917.160 1261.555 ;
        RECT 2916.950 1260.875 2917.230 1261.245 ;
        RECT 2884.290 1256.115 2884.570 1256.485 ;
      LAYER via2 ;
        RECT 984.030 2614.800 984.310 2615.080 ;
        RECT 1048.430 2614.800 1048.710 2615.080 ;
        RECT 1048.430 2613.440 1048.710 2613.720 ;
        RECT 2884.290 1261.600 2884.570 1261.880 ;
        RECT 2916.950 1261.600 2917.230 1261.880 ;
        RECT 2916.950 1260.920 2917.230 1261.200 ;
        RECT 2884.290 1256.160 2884.570 1256.440 ;
      LAYER met3 ;
        RECT 984.005 2615.090 984.335 2615.105 ;
        RECT 1048.405 2615.090 1048.735 2615.105 ;
        RECT 984.005 2614.790 1048.735 2615.090 ;
        RECT 984.005 2614.775 984.335 2614.790 ;
        RECT 1048.405 2614.775 1048.735 2614.790 ;
        RECT 1048.405 2613.730 1048.735 2613.745 ;
        RECT 1797.030 2613.730 1797.410 2613.740 ;
        RECT 1048.405 2613.430 1797.410 2613.730 ;
        RECT 1048.405 2613.415 1048.735 2613.430 ;
        RECT 1797.030 2613.420 1797.410 2613.430 ;
        RECT 2884.265 1261.890 2884.595 1261.905 ;
        RECT 2916.925 1261.890 2917.255 1261.905 ;
        RECT 2884.265 1261.590 2917.255 1261.890 ;
        RECT 2884.265 1261.575 2884.595 1261.590 ;
        RECT 2916.925 1261.575 2917.255 1261.590 ;
        RECT 2916.925 1261.210 2917.255 1261.225 ;
        RECT 2918.000 1261.210 2924.000 1261.660 ;
        RECT 2916.925 1260.910 2924.000 1261.210 ;
        RECT 2916.925 1260.895 2917.255 1260.910 ;
        RECT 2918.000 1260.460 2924.000 1260.910 ;
        RECT 1821.910 1257.510 1870.050 1257.810 ;
        RECT 1797.030 1256.450 1797.410 1256.460 ;
        RECT 1821.910 1256.450 1822.210 1257.510 ;
        RECT 1869.750 1257.130 1870.050 1257.510 ;
        RECT 1918.510 1257.510 1966.650 1257.810 ;
        RECT 1869.750 1256.830 1917.890 1257.130 ;
        RECT 1797.030 1256.150 1822.210 1256.450 ;
        RECT 1917.590 1256.450 1917.890 1256.830 ;
        RECT 1918.510 1256.450 1918.810 1257.510 ;
        RECT 1966.350 1257.130 1966.650 1257.510 ;
        RECT 2015.110 1257.510 2063.250 1257.810 ;
        RECT 1966.350 1256.830 2014.490 1257.130 ;
        RECT 1917.590 1256.150 1918.810 1256.450 ;
        RECT 2014.190 1256.450 2014.490 1256.830 ;
        RECT 2015.110 1256.450 2015.410 1257.510 ;
        RECT 2062.950 1257.130 2063.250 1257.510 ;
        RECT 2111.710 1257.510 2159.850 1257.810 ;
        RECT 2062.950 1256.830 2111.090 1257.130 ;
        RECT 2014.190 1256.150 2015.410 1256.450 ;
        RECT 2110.790 1256.450 2111.090 1256.830 ;
        RECT 2111.710 1256.450 2112.010 1257.510 ;
        RECT 2159.550 1257.130 2159.850 1257.510 ;
        RECT 2208.310 1257.510 2256.450 1257.810 ;
        RECT 2159.550 1256.830 2207.690 1257.130 ;
        RECT 2110.790 1256.150 2112.010 1256.450 ;
        RECT 2207.390 1256.450 2207.690 1256.830 ;
        RECT 2208.310 1256.450 2208.610 1257.510 ;
        RECT 2256.150 1257.130 2256.450 1257.510 ;
        RECT 2304.910 1257.510 2353.050 1257.810 ;
        RECT 2256.150 1256.830 2304.290 1257.130 ;
        RECT 2207.390 1256.150 2208.610 1256.450 ;
        RECT 2303.990 1256.450 2304.290 1256.830 ;
        RECT 2304.910 1256.450 2305.210 1257.510 ;
        RECT 2352.750 1257.130 2353.050 1257.510 ;
        RECT 2401.510 1257.510 2449.650 1257.810 ;
        RECT 2352.750 1256.830 2400.890 1257.130 ;
        RECT 2303.990 1256.150 2305.210 1256.450 ;
        RECT 2400.590 1256.450 2400.890 1256.830 ;
        RECT 2401.510 1256.450 2401.810 1257.510 ;
        RECT 2449.350 1257.130 2449.650 1257.510 ;
        RECT 2498.110 1257.510 2546.250 1257.810 ;
        RECT 2449.350 1256.830 2497.490 1257.130 ;
        RECT 2400.590 1256.150 2401.810 1256.450 ;
        RECT 2497.190 1256.450 2497.490 1256.830 ;
        RECT 2498.110 1256.450 2498.410 1257.510 ;
        RECT 2545.950 1257.130 2546.250 1257.510 ;
        RECT 2594.710 1257.510 2642.850 1257.810 ;
        RECT 2545.950 1256.830 2594.090 1257.130 ;
        RECT 2497.190 1256.150 2498.410 1256.450 ;
        RECT 2593.790 1256.450 2594.090 1256.830 ;
        RECT 2594.710 1256.450 2595.010 1257.510 ;
        RECT 2642.550 1257.130 2642.850 1257.510 ;
        RECT 2691.310 1257.510 2739.450 1257.810 ;
        RECT 2642.550 1256.830 2690.690 1257.130 ;
        RECT 2593.790 1256.150 2595.010 1256.450 ;
        RECT 2690.390 1256.450 2690.690 1256.830 ;
        RECT 2691.310 1256.450 2691.610 1257.510 ;
        RECT 2739.150 1257.130 2739.450 1257.510 ;
        RECT 2787.910 1257.510 2836.050 1257.810 ;
        RECT 2739.150 1256.830 2787.290 1257.130 ;
        RECT 2690.390 1256.150 2691.610 1256.450 ;
        RECT 2786.990 1256.450 2787.290 1256.830 ;
        RECT 2787.910 1256.450 2788.210 1257.510 ;
        RECT 2835.750 1257.130 2836.050 1257.510 ;
        RECT 2835.750 1256.830 2883.890 1257.130 ;
        RECT 2786.990 1256.150 2788.210 1256.450 ;
        RECT 2883.590 1256.450 2883.890 1256.830 ;
        RECT 2884.265 1256.450 2884.595 1256.465 ;
        RECT 2883.590 1256.150 2884.595 1256.450 ;
        RECT 1797.030 1256.140 1797.410 1256.150 ;
        RECT 2884.265 1256.135 2884.595 1256.150 ;
      LAYER via3 ;
        RECT 1797.060 2613.420 1797.380 2613.740 ;
        RECT 1797.060 1256.140 1797.380 1256.460 ;
      LAYER met4 ;
        RECT 1797.055 2613.415 1797.385 2613.745 ;
        RECT 1797.070 1256.465 1797.370 2613.415 ;
        RECT 1797.055 1256.135 1797.385 1256.465 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1009.790 2614.075 1010.070 2614.445 ;
        RECT 1007.870 2599.370 1008.150 2600.000 ;
        RECT 1009.860 2599.370 1010.000 2614.075 ;
        RECT 1007.870 2599.230 1010.000 2599.370 ;
        RECT 1007.870 2596.000 1008.150 2599.230 ;
        RECT 2884.290 1496.155 2884.570 1496.525 ;
        RECT 2916.950 1496.155 2917.230 1496.525 ;
        RECT 2884.360 1491.085 2884.500 1496.155 ;
        RECT 2917.020 1495.845 2917.160 1496.155 ;
        RECT 2916.950 1495.475 2917.230 1495.845 ;
        RECT 2884.290 1490.715 2884.570 1491.085 ;
      LAYER via2 ;
        RECT 1009.790 2614.120 1010.070 2614.400 ;
        RECT 2884.290 1496.200 2884.570 1496.480 ;
        RECT 2916.950 1496.200 2917.230 1496.480 ;
        RECT 2916.950 1495.520 2917.230 1495.800 ;
        RECT 2884.290 1490.760 2884.570 1491.040 ;
      LAYER met3 ;
        RECT 1009.765 2614.410 1010.095 2614.425 ;
        RECT 1797.950 2614.410 1798.330 2614.420 ;
        RECT 1009.765 2614.110 1798.330 2614.410 ;
        RECT 1009.765 2614.095 1010.095 2614.110 ;
        RECT 1797.950 2614.100 1798.330 2614.110 ;
        RECT 2884.265 1496.490 2884.595 1496.505 ;
        RECT 2916.925 1496.490 2917.255 1496.505 ;
        RECT 2884.265 1496.190 2917.255 1496.490 ;
        RECT 2884.265 1496.175 2884.595 1496.190 ;
        RECT 2916.925 1496.175 2917.255 1496.190 ;
        RECT 2916.925 1495.810 2917.255 1495.825 ;
        RECT 2918.000 1495.810 2924.000 1496.260 ;
        RECT 2916.925 1495.510 2924.000 1495.810 ;
        RECT 2916.925 1495.495 2917.255 1495.510 ;
        RECT 2918.000 1495.060 2924.000 1495.510 ;
        RECT 1821.910 1492.110 1870.050 1492.410 ;
        RECT 1797.950 1491.050 1798.330 1491.060 ;
        RECT 1821.910 1491.050 1822.210 1492.110 ;
        RECT 1869.750 1491.730 1870.050 1492.110 ;
        RECT 1918.510 1492.110 1966.650 1492.410 ;
        RECT 1869.750 1491.430 1917.890 1491.730 ;
        RECT 1797.950 1490.750 1822.210 1491.050 ;
        RECT 1917.590 1491.050 1917.890 1491.430 ;
        RECT 1918.510 1491.050 1918.810 1492.110 ;
        RECT 1966.350 1491.730 1966.650 1492.110 ;
        RECT 2015.110 1492.110 2063.250 1492.410 ;
        RECT 1966.350 1491.430 2014.490 1491.730 ;
        RECT 1917.590 1490.750 1918.810 1491.050 ;
        RECT 2014.190 1491.050 2014.490 1491.430 ;
        RECT 2015.110 1491.050 2015.410 1492.110 ;
        RECT 2062.950 1491.730 2063.250 1492.110 ;
        RECT 2111.710 1492.110 2159.850 1492.410 ;
        RECT 2062.950 1491.430 2111.090 1491.730 ;
        RECT 2014.190 1490.750 2015.410 1491.050 ;
        RECT 2110.790 1491.050 2111.090 1491.430 ;
        RECT 2111.710 1491.050 2112.010 1492.110 ;
        RECT 2159.550 1491.730 2159.850 1492.110 ;
        RECT 2208.310 1492.110 2256.450 1492.410 ;
        RECT 2159.550 1491.430 2207.690 1491.730 ;
        RECT 2110.790 1490.750 2112.010 1491.050 ;
        RECT 2207.390 1491.050 2207.690 1491.430 ;
        RECT 2208.310 1491.050 2208.610 1492.110 ;
        RECT 2256.150 1491.730 2256.450 1492.110 ;
        RECT 2304.910 1492.110 2353.050 1492.410 ;
        RECT 2256.150 1491.430 2304.290 1491.730 ;
        RECT 2207.390 1490.750 2208.610 1491.050 ;
        RECT 2303.990 1491.050 2304.290 1491.430 ;
        RECT 2304.910 1491.050 2305.210 1492.110 ;
        RECT 2352.750 1491.730 2353.050 1492.110 ;
        RECT 2401.510 1492.110 2449.650 1492.410 ;
        RECT 2352.750 1491.430 2400.890 1491.730 ;
        RECT 2303.990 1490.750 2305.210 1491.050 ;
        RECT 2400.590 1491.050 2400.890 1491.430 ;
        RECT 2401.510 1491.050 2401.810 1492.110 ;
        RECT 2449.350 1491.730 2449.650 1492.110 ;
        RECT 2498.110 1492.110 2546.250 1492.410 ;
        RECT 2449.350 1491.430 2497.490 1491.730 ;
        RECT 2400.590 1490.750 2401.810 1491.050 ;
        RECT 2497.190 1491.050 2497.490 1491.430 ;
        RECT 2498.110 1491.050 2498.410 1492.110 ;
        RECT 2545.950 1491.730 2546.250 1492.110 ;
        RECT 2594.710 1492.110 2642.850 1492.410 ;
        RECT 2545.950 1491.430 2594.090 1491.730 ;
        RECT 2497.190 1490.750 2498.410 1491.050 ;
        RECT 2593.790 1491.050 2594.090 1491.430 ;
        RECT 2594.710 1491.050 2595.010 1492.110 ;
        RECT 2642.550 1491.730 2642.850 1492.110 ;
        RECT 2691.310 1492.110 2739.450 1492.410 ;
        RECT 2642.550 1491.430 2690.690 1491.730 ;
        RECT 2593.790 1490.750 2595.010 1491.050 ;
        RECT 2690.390 1491.050 2690.690 1491.430 ;
        RECT 2691.310 1491.050 2691.610 1492.110 ;
        RECT 2739.150 1491.730 2739.450 1492.110 ;
        RECT 2787.910 1492.110 2836.050 1492.410 ;
        RECT 2739.150 1491.430 2787.290 1491.730 ;
        RECT 2690.390 1490.750 2691.610 1491.050 ;
        RECT 2786.990 1491.050 2787.290 1491.430 ;
        RECT 2787.910 1491.050 2788.210 1492.110 ;
        RECT 2835.750 1491.730 2836.050 1492.110 ;
        RECT 2835.750 1491.430 2883.890 1491.730 ;
        RECT 2786.990 1490.750 2788.210 1491.050 ;
        RECT 2883.590 1491.050 2883.890 1491.430 ;
        RECT 2884.265 1491.050 2884.595 1491.065 ;
        RECT 2883.590 1490.750 2884.595 1491.050 ;
        RECT 1797.950 1490.740 1798.330 1490.750 ;
        RECT 2884.265 1490.735 2884.595 1490.750 ;
      LAYER via3 ;
        RECT 1797.980 2614.100 1798.300 2614.420 ;
        RECT 1797.980 1490.740 1798.300 1491.060 ;
      LAYER met4 ;
        RECT 1797.975 2614.095 1798.305 2614.425 ;
        RECT 1797.990 1491.065 1798.290 2614.095 ;
        RECT 1797.975 1490.735 1798.305 1491.065 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1034.610 2602.600 1034.930 2602.660 ;
        RECT 1847.890 2602.600 1848.210 2602.660 ;
        RECT 1034.610 2602.460 1848.210 2602.600 ;
        RECT 1034.610 2602.400 1034.930 2602.460 ;
        RECT 1847.890 2602.400 1848.210 2602.460 ;
        RECT 1847.890 1731.860 1848.210 1731.920 ;
        RECT 2900.370 1731.860 2900.690 1731.920 ;
        RECT 1847.890 1731.720 2900.690 1731.860 ;
        RECT 1847.890 1731.660 1848.210 1731.720 ;
        RECT 2900.370 1731.660 2900.690 1731.720 ;
      LAYER via ;
        RECT 1034.640 2602.400 1034.900 2602.660 ;
        RECT 1847.920 2602.400 1848.180 2602.660 ;
        RECT 1847.920 1731.660 1848.180 1731.920 ;
        RECT 2900.400 1731.660 2900.660 1731.920 ;
      LAYER met2 ;
        RECT 1034.640 2602.370 1034.900 2602.690 ;
        RECT 1847.920 2602.370 1848.180 2602.690 ;
        RECT 1033.630 2599.370 1033.910 2600.000 ;
        RECT 1034.700 2599.370 1034.840 2602.370 ;
        RECT 1033.630 2599.230 1034.840 2599.370 ;
        RECT 1033.630 2596.000 1033.910 2599.230 ;
        RECT 1847.980 1731.950 1848.120 2602.370 ;
        RECT 1847.920 1731.630 1848.180 1731.950 ;
        RECT 2900.400 1731.630 2900.660 1731.950 ;
        RECT 2900.460 1730.445 2900.600 1731.630 ;
        RECT 2900.390 1730.075 2900.670 1730.445 ;
      LAYER via2 ;
        RECT 2900.390 1730.120 2900.670 1730.400 ;
      LAYER met3 ;
        RECT 2900.365 1730.410 2900.695 1730.425 ;
        RECT 2918.000 1730.410 2924.000 1730.860 ;
        RECT 2900.365 1730.110 2924.000 1730.410 ;
        RECT 2900.365 1730.095 2900.695 1730.110 ;
        RECT 2918.000 1729.660 2924.000 1730.110 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1060.370 2603.280 1060.690 2603.340 ;
        RECT 1852.950 2603.280 1853.270 2603.340 ;
        RECT 1060.370 2603.140 1853.270 2603.280 ;
        RECT 1060.370 2603.080 1060.690 2603.140 ;
        RECT 1852.950 2603.080 1853.270 2603.140 ;
        RECT 1852.950 1966.460 1853.270 1966.520 ;
        RECT 2899.450 1966.460 2899.770 1966.520 ;
        RECT 1852.950 1966.320 2899.770 1966.460 ;
        RECT 1852.950 1966.260 1853.270 1966.320 ;
        RECT 2899.450 1966.260 2899.770 1966.320 ;
      LAYER via ;
        RECT 1060.400 2603.080 1060.660 2603.340 ;
        RECT 1852.980 2603.080 1853.240 2603.340 ;
        RECT 1852.980 1966.260 1853.240 1966.520 ;
        RECT 2899.480 1966.260 2899.740 1966.520 ;
      LAYER met2 ;
        RECT 1060.400 2603.050 1060.660 2603.370 ;
        RECT 1852.980 2603.050 1853.240 2603.370 ;
        RECT 1058.930 2599.370 1059.210 2600.000 ;
        RECT 1060.460 2599.370 1060.600 2603.050 ;
        RECT 1058.930 2599.230 1060.600 2599.370 ;
        RECT 1058.930 2596.000 1059.210 2599.230 ;
        RECT 1853.040 1966.550 1853.180 2603.050 ;
        RECT 1852.980 1966.230 1853.240 1966.550 ;
        RECT 2899.480 1966.230 2899.740 1966.550 ;
        RECT 2899.540 1965.045 2899.680 1966.230 ;
        RECT 2899.470 1964.675 2899.750 1965.045 ;
      LAYER via2 ;
        RECT 2899.470 1964.720 2899.750 1965.000 ;
      LAYER met3 ;
        RECT 2899.445 1965.010 2899.775 1965.025 ;
        RECT 2918.000 1965.010 2924.000 1965.460 ;
        RECT 2899.445 1964.710 2924.000 1965.010 ;
        RECT 2899.445 1964.695 2899.775 1964.710 ;
        RECT 2918.000 1964.260 2924.000 1964.710 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1086.130 2603.620 1086.450 2603.680 ;
        RECT 1854.330 2603.620 1854.650 2603.680 ;
        RECT 1086.130 2603.480 1854.650 2603.620 ;
        RECT 1086.130 2603.420 1086.450 2603.480 ;
        RECT 1854.330 2603.420 1854.650 2603.480 ;
        RECT 1854.330 2201.060 1854.650 2201.120 ;
        RECT 2899.450 2201.060 2899.770 2201.120 ;
        RECT 1854.330 2200.920 2899.770 2201.060 ;
        RECT 1854.330 2200.860 1854.650 2200.920 ;
        RECT 2899.450 2200.860 2899.770 2200.920 ;
      LAYER via ;
        RECT 1086.160 2603.420 1086.420 2603.680 ;
        RECT 1854.360 2603.420 1854.620 2603.680 ;
        RECT 1854.360 2200.860 1854.620 2201.120 ;
        RECT 2899.480 2200.860 2899.740 2201.120 ;
      LAYER met2 ;
        RECT 1086.160 2603.390 1086.420 2603.710 ;
        RECT 1854.360 2603.390 1854.620 2603.710 ;
        RECT 1084.690 2599.370 1084.970 2600.000 ;
        RECT 1086.220 2599.370 1086.360 2603.390 ;
        RECT 1084.690 2599.230 1086.360 2599.370 ;
        RECT 1084.690 2596.000 1084.970 2599.230 ;
        RECT 1854.420 2201.150 1854.560 2603.390 ;
        RECT 1854.360 2200.830 1854.620 2201.150 ;
        RECT 2899.480 2200.830 2899.740 2201.150 ;
        RECT 2899.540 2199.645 2899.680 2200.830 ;
        RECT 2899.470 2199.275 2899.750 2199.645 ;
      LAYER via2 ;
        RECT 2899.470 2199.320 2899.750 2199.600 ;
      LAYER met3 ;
        RECT 2899.445 2199.610 2899.775 2199.625 ;
        RECT 2918.000 2199.610 2924.000 2200.060 ;
        RECT 2899.445 2199.310 2924.000 2199.610 ;
        RECT 2899.445 2199.295 2899.775 2199.310 ;
        RECT 2918.000 2198.860 2924.000 2199.310 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1835.470 201.520 1835.790 201.580 ;
        RECT 1849.730 201.520 1850.050 201.580 ;
        RECT 1835.470 201.380 1850.050 201.520 ;
        RECT 1835.470 201.320 1835.790 201.380 ;
        RECT 1849.730 201.320 1850.050 201.380 ;
        RECT 1352.470 201.180 1352.790 201.240 ;
        RECT 1378.690 201.180 1379.010 201.240 ;
        RECT 1352.470 201.040 1379.010 201.180 ;
        RECT 1352.470 200.980 1352.790 201.040 ;
        RECT 1378.690 200.980 1379.010 201.040 ;
        RECT 1993.710 201.180 1994.030 201.240 ;
        RECT 2028.210 201.180 2028.530 201.240 ;
        RECT 1993.710 201.040 2028.530 201.180 ;
        RECT 1993.710 200.980 1994.030 201.040 ;
        RECT 2028.210 200.980 2028.530 201.040 ;
        RECT 1062.210 200.500 1062.530 200.560 ;
        RECT 1103.610 200.500 1103.930 200.560 ;
        RECT 1062.210 200.360 1103.930 200.500 ;
        RECT 1062.210 200.300 1062.530 200.360 ;
        RECT 1103.610 200.300 1103.930 200.360 ;
        RECT 1007.470 199.820 1007.790 199.880 ;
        RECT 1009.310 199.820 1009.630 199.880 ;
        RECT 1007.470 199.680 1009.630 199.820 ;
        RECT 1007.470 199.620 1007.790 199.680 ;
        RECT 1009.310 199.620 1009.630 199.680 ;
      LAYER via ;
        RECT 1835.500 201.320 1835.760 201.580 ;
        RECT 1849.760 201.320 1850.020 201.580 ;
        RECT 1352.500 200.980 1352.760 201.240 ;
        RECT 1378.720 200.980 1378.980 201.240 ;
        RECT 1993.740 200.980 1994.000 201.240 ;
        RECT 2028.240 200.980 2028.500 201.240 ;
        RECT 1062.240 200.300 1062.500 200.560 ;
        RECT 1103.640 200.300 1103.900 200.560 ;
        RECT 1007.500 199.620 1007.760 199.880 ;
        RECT 1009.340 199.620 1009.600 199.880 ;
      LAYER met2 ;
        RECT 862.510 2596.650 862.790 2600.000 ;
        RECT 864.430 2596.650 864.710 2596.765 ;
        RECT 862.510 2596.510 864.710 2596.650 ;
        RECT 862.510 2596.000 862.790 2596.510 ;
        RECT 864.430 2596.395 864.710 2596.510 ;
        RECT 2884.290 205.515 2884.570 205.885 ;
        RECT 2916.950 205.515 2917.230 205.885 ;
        RECT 1691.050 202.795 1691.330 203.165 ;
        RECT 1449.550 201.435 1449.830 201.805 ;
        RECT 1352.500 201.125 1352.760 201.270 ;
        RECT 1378.720 201.125 1378.980 201.270 ;
        RECT 1103.630 200.755 1103.910 201.125 ;
        RECT 1352.490 200.755 1352.770 201.125 ;
        RECT 1378.710 200.755 1378.990 201.125 ;
        RECT 1449.090 201.010 1449.370 201.125 ;
        RECT 1449.620 201.010 1449.760 201.435 ;
        RECT 1691.120 201.125 1691.260 202.795 ;
        RECT 1973.030 202.115 1973.310 202.485 ;
        RECT 1835.490 201.435 1835.770 201.805 ;
        RECT 1835.500 201.290 1835.760 201.435 ;
        RECT 1849.760 201.290 1850.020 201.610 ;
        RECT 1449.090 200.870 1449.760 201.010 ;
        RECT 1449.090 200.755 1449.370 200.870 ;
        RECT 1691.050 200.755 1691.330 201.125 ;
        RECT 1103.700 200.590 1103.840 200.755 ;
        RECT 1062.240 200.445 1062.500 200.590 ;
        RECT 1009.330 200.075 1009.610 200.445 ;
        RECT 1062.230 200.075 1062.510 200.445 ;
        RECT 1103.640 200.270 1103.900 200.590 ;
        RECT 1849.820 200.445 1849.960 201.290 ;
        RECT 1898.050 201.010 1898.330 201.125 ;
        RECT 1897.200 200.870 1898.330 201.010 ;
        RECT 1897.200 200.445 1897.340 200.870 ;
        RECT 1898.050 200.755 1898.330 200.870 ;
        RECT 1973.100 200.445 1973.240 202.115 ;
        RECT 2028.230 201.435 2028.510 201.805 ;
        RECT 2028.300 201.270 2028.440 201.435 ;
        RECT 1993.740 201.125 1994.000 201.270 ;
        RECT 1993.730 200.755 1994.010 201.125 ;
        RECT 2028.240 200.950 2028.500 201.270 ;
        RECT 2884.360 200.445 2884.500 205.515 ;
        RECT 2917.020 205.205 2917.160 205.515 ;
        RECT 2916.950 204.835 2917.230 205.205 ;
        RECT 1849.750 200.075 1850.030 200.445 ;
        RECT 1897.130 200.075 1897.410 200.445 ;
        RECT 1973.030 200.075 1973.310 200.445 ;
        RECT 2884.290 200.075 2884.570 200.445 ;
        RECT 1009.400 199.910 1009.540 200.075 ;
        RECT 1007.500 199.765 1007.760 199.910 ;
        RECT 1007.490 199.395 1007.770 199.765 ;
        RECT 1009.340 199.590 1009.600 199.910 ;
      LAYER via2 ;
        RECT 864.430 2596.440 864.710 2596.720 ;
        RECT 2884.290 205.560 2884.570 205.840 ;
        RECT 2916.950 205.560 2917.230 205.840 ;
        RECT 1691.050 202.840 1691.330 203.120 ;
        RECT 1449.550 201.480 1449.830 201.760 ;
        RECT 1103.630 200.800 1103.910 201.080 ;
        RECT 1352.490 200.800 1352.770 201.080 ;
        RECT 1378.710 200.800 1378.990 201.080 ;
        RECT 1449.090 200.800 1449.370 201.080 ;
        RECT 1973.030 202.160 1973.310 202.440 ;
        RECT 1835.490 201.480 1835.770 201.760 ;
        RECT 1691.050 200.800 1691.330 201.080 ;
        RECT 1009.330 200.120 1009.610 200.400 ;
        RECT 1062.230 200.120 1062.510 200.400 ;
        RECT 1898.050 200.800 1898.330 201.080 ;
        RECT 2028.230 201.480 2028.510 201.760 ;
        RECT 1993.730 200.800 1994.010 201.080 ;
        RECT 2916.950 204.880 2917.230 205.160 ;
        RECT 1849.750 200.120 1850.030 200.400 ;
        RECT 1897.130 200.120 1897.410 200.400 ;
        RECT 1973.030 200.120 1973.310 200.400 ;
        RECT 2884.290 200.120 2884.570 200.400 ;
        RECT 1007.490 199.440 1007.770 199.720 ;
      LAYER met3 ;
        RECT 864.405 2596.730 864.735 2596.745 ;
        RECT 866.910 2596.730 867.290 2596.740 ;
        RECT 864.405 2596.430 867.290 2596.730 ;
        RECT 864.405 2596.415 864.735 2596.430 ;
        RECT 866.910 2596.420 867.290 2596.430 ;
        RECT 2884.265 205.850 2884.595 205.865 ;
        RECT 2916.925 205.850 2917.255 205.865 ;
        RECT 2884.265 205.550 2917.255 205.850 ;
        RECT 2884.265 205.535 2884.595 205.550 ;
        RECT 2916.925 205.535 2917.255 205.550 ;
        RECT 2916.925 205.170 2917.255 205.185 ;
        RECT 2918.000 205.170 2924.000 205.620 ;
        RECT 2916.925 204.870 2924.000 205.170 ;
        RECT 2916.925 204.855 2917.255 204.870 ;
        RECT 2918.000 204.420 2924.000 204.870 ;
        RECT 1635.110 203.130 1635.490 203.140 ;
        RECT 1683.870 203.130 1684.250 203.140 ;
        RECT 1691.025 203.130 1691.355 203.145 ;
        RECT 1635.110 202.830 1683.290 203.130 ;
        RECT 1635.110 202.820 1635.490 202.830 ;
        RECT 1682.990 202.460 1683.290 202.830 ;
        RECT 1683.870 202.830 1691.355 203.130 ;
        RECT 1683.870 202.820 1684.250 202.830 ;
        RECT 1691.025 202.815 1691.355 202.830 ;
        RECT 1538.510 202.450 1538.890 202.460 ;
        RECT 1538.510 202.150 1586.690 202.450 ;
        RECT 1538.510 202.140 1538.890 202.150 ;
        RECT 866.910 201.770 867.290 201.780 ;
        RECT 1449.525 201.770 1449.855 201.785 ;
        RECT 1586.390 201.770 1586.690 202.150 ;
        RECT 1606.630 202.150 1611.530 202.450 ;
        RECT 1606.630 201.770 1606.930 202.150 ;
        RECT 866.910 201.470 883.810 201.770 ;
        RECT 866.910 201.460 867.290 201.470 ;
        RECT 883.510 201.090 883.810 201.470 ;
        RECT 1161.350 201.470 1321.730 201.770 ;
        RECT 1103.605 201.090 1103.935 201.105 ;
        RECT 883.510 200.790 959.250 201.090 ;
        RECT 958.950 200.410 959.250 200.790 ;
        RECT 1103.605 200.790 1110.130 201.090 ;
        RECT 1103.605 200.775 1103.935 200.790 ;
        RECT 1109.830 200.580 1110.130 200.790 ;
        RECT 1009.305 200.410 1009.635 200.425 ;
        RECT 1062.205 200.410 1062.535 200.425 ;
        RECT 958.950 200.110 960.170 200.410 ;
        RECT 959.870 199.730 960.170 200.110 ;
        RECT 1009.305 200.110 1062.535 200.410 ;
        RECT 1109.830 200.410 1111.970 200.580 ;
        RECT 1161.350 200.410 1161.650 201.470 ;
        RECT 1321.430 201.090 1321.730 201.470 ;
        RECT 1449.525 201.470 1521.370 201.770 ;
        RECT 1586.390 201.470 1606.930 201.770 ;
        RECT 1449.525 201.455 1449.855 201.470 ;
        RECT 1352.465 201.090 1352.795 201.105 ;
        RECT 1321.430 200.790 1352.795 201.090 ;
        RECT 1352.465 200.775 1352.795 200.790 ;
        RECT 1378.685 201.090 1379.015 201.105 ;
        RECT 1449.065 201.090 1449.395 201.105 ;
        RECT 1378.685 200.790 1449.395 201.090 ;
        RECT 1521.070 201.090 1521.370 201.470 ;
        RECT 1538.510 201.090 1538.890 201.100 ;
        RECT 1521.070 200.790 1538.890 201.090 ;
        RECT 1611.230 201.090 1611.530 202.150 ;
        RECT 1682.950 202.140 1683.330 202.460 ;
        RECT 1924.910 202.450 1925.290 202.460 ;
        RECT 1973.005 202.450 1973.335 202.465 ;
        RECT 1924.910 202.150 1973.335 202.450 ;
        RECT 1924.910 202.140 1925.290 202.150 ;
        RECT 1973.005 202.135 1973.335 202.150 ;
        RECT 1635.110 201.460 1635.490 201.780 ;
        RECT 1835.465 201.770 1835.795 201.785 ;
        RECT 1800.750 201.470 1835.795 201.770 ;
        RECT 1635.150 201.090 1635.450 201.460 ;
        RECT 1611.230 200.790 1635.450 201.090 ;
        RECT 1691.025 201.090 1691.355 201.105 ;
        RECT 1691.025 200.790 1739.410 201.090 ;
        RECT 1378.685 200.775 1379.015 200.790 ;
        RECT 1449.065 200.775 1449.395 200.790 ;
        RECT 1538.510 200.780 1538.890 200.790 ;
        RECT 1691.025 200.775 1691.355 200.790 ;
        RECT 1109.830 200.280 1161.650 200.410 ;
        RECT 1111.670 200.110 1161.650 200.280 ;
        RECT 1739.110 200.410 1739.410 200.790 ;
        RECT 1800.750 200.410 1801.050 201.470 ;
        RECT 1835.465 201.455 1835.795 201.470 ;
        RECT 2028.205 201.770 2028.535 201.785 ;
        RECT 2028.205 201.470 2063.250 201.770 ;
        RECT 2028.205 201.455 2028.535 201.470 ;
        RECT 1898.025 201.090 1898.355 201.105 ;
        RECT 1924.910 201.090 1925.290 201.100 ;
        RECT 1993.705 201.090 1994.035 201.105 ;
        RECT 1898.025 200.790 1925.290 201.090 ;
        RECT 1898.025 200.775 1898.355 200.790 ;
        RECT 1924.910 200.780 1925.290 200.790 ;
        RECT 1980.150 200.790 1994.035 201.090 ;
        RECT 2062.950 201.090 2063.250 201.470 ;
        RECT 2111.710 201.470 2159.850 201.770 ;
        RECT 2062.950 200.790 2111.090 201.090 ;
        RECT 1739.110 200.110 1801.050 200.410 ;
        RECT 1849.725 200.410 1850.055 200.425 ;
        RECT 1897.105 200.410 1897.435 200.425 ;
        RECT 1849.725 200.110 1897.435 200.410 ;
        RECT 1009.305 200.095 1009.635 200.110 ;
        RECT 1062.205 200.095 1062.535 200.110 ;
        RECT 1849.725 200.095 1850.055 200.110 ;
        RECT 1897.105 200.095 1897.435 200.110 ;
        RECT 1973.005 200.410 1973.335 200.425 ;
        RECT 1980.150 200.410 1980.450 200.790 ;
        RECT 1993.705 200.775 1994.035 200.790 ;
        RECT 1973.005 200.110 1980.450 200.410 ;
        RECT 2110.790 200.410 2111.090 200.790 ;
        RECT 2111.710 200.410 2112.010 201.470 ;
        RECT 2159.550 201.090 2159.850 201.470 ;
        RECT 2208.310 201.470 2256.450 201.770 ;
        RECT 2159.550 200.790 2207.690 201.090 ;
        RECT 2110.790 200.110 2112.010 200.410 ;
        RECT 2207.390 200.410 2207.690 200.790 ;
        RECT 2208.310 200.410 2208.610 201.470 ;
        RECT 2256.150 201.090 2256.450 201.470 ;
        RECT 2304.910 201.470 2353.050 201.770 ;
        RECT 2256.150 200.790 2304.290 201.090 ;
        RECT 2207.390 200.110 2208.610 200.410 ;
        RECT 2303.990 200.410 2304.290 200.790 ;
        RECT 2304.910 200.410 2305.210 201.470 ;
        RECT 2352.750 201.090 2353.050 201.470 ;
        RECT 2401.510 201.470 2449.650 201.770 ;
        RECT 2352.750 200.790 2400.890 201.090 ;
        RECT 2303.990 200.110 2305.210 200.410 ;
        RECT 2400.590 200.410 2400.890 200.790 ;
        RECT 2401.510 200.410 2401.810 201.470 ;
        RECT 2449.350 201.090 2449.650 201.470 ;
        RECT 2498.110 201.470 2546.250 201.770 ;
        RECT 2449.350 200.790 2497.490 201.090 ;
        RECT 2400.590 200.110 2401.810 200.410 ;
        RECT 2497.190 200.410 2497.490 200.790 ;
        RECT 2498.110 200.410 2498.410 201.470 ;
        RECT 2545.950 201.090 2546.250 201.470 ;
        RECT 2594.710 201.470 2642.850 201.770 ;
        RECT 2545.950 200.790 2594.090 201.090 ;
        RECT 2497.190 200.110 2498.410 200.410 ;
        RECT 2593.790 200.410 2594.090 200.790 ;
        RECT 2594.710 200.410 2595.010 201.470 ;
        RECT 2642.550 201.090 2642.850 201.470 ;
        RECT 2691.310 201.470 2739.450 201.770 ;
        RECT 2642.550 200.790 2690.690 201.090 ;
        RECT 2593.790 200.110 2595.010 200.410 ;
        RECT 2690.390 200.410 2690.690 200.790 ;
        RECT 2691.310 200.410 2691.610 201.470 ;
        RECT 2739.150 201.090 2739.450 201.470 ;
        RECT 2787.910 201.470 2836.050 201.770 ;
        RECT 2739.150 200.790 2787.290 201.090 ;
        RECT 2690.390 200.110 2691.610 200.410 ;
        RECT 2786.990 200.410 2787.290 200.790 ;
        RECT 2787.910 200.410 2788.210 201.470 ;
        RECT 2835.750 201.090 2836.050 201.470 ;
        RECT 2835.750 200.790 2883.890 201.090 ;
        RECT 2786.990 200.110 2788.210 200.410 ;
        RECT 2883.590 200.410 2883.890 200.790 ;
        RECT 2884.265 200.410 2884.595 200.425 ;
        RECT 2883.590 200.110 2884.595 200.410 ;
        RECT 1973.005 200.095 1973.335 200.110 ;
        RECT 2884.265 200.095 2884.595 200.110 ;
        RECT 1007.465 199.730 1007.795 199.745 ;
        RECT 959.870 199.430 1007.795 199.730 ;
        RECT 1007.465 199.415 1007.795 199.430 ;
      LAYER via3 ;
        RECT 866.940 2596.420 867.260 2596.740 ;
        RECT 1635.140 202.820 1635.460 203.140 ;
        RECT 1683.900 202.820 1684.220 203.140 ;
        RECT 1538.540 202.140 1538.860 202.460 ;
        RECT 866.940 201.460 867.260 201.780 ;
        RECT 1538.540 200.780 1538.860 201.100 ;
        RECT 1682.980 202.140 1683.300 202.460 ;
        RECT 1924.940 202.140 1925.260 202.460 ;
        RECT 1635.140 201.460 1635.460 201.780 ;
        RECT 1924.940 200.780 1925.260 201.100 ;
      LAYER met4 ;
        RECT 866.935 2596.415 867.265 2596.745 ;
        RECT 866.950 201.785 867.250 2596.415 ;
        RECT 1635.135 202.815 1635.465 203.145 ;
        RECT 1683.895 202.815 1684.225 203.145 ;
        RECT 1538.535 202.135 1538.865 202.465 ;
        RECT 866.935 201.455 867.265 201.785 ;
        RECT 1538.550 201.105 1538.850 202.135 ;
        RECT 1635.150 201.785 1635.450 202.815 ;
        RECT 1682.975 202.450 1683.305 202.465 ;
        RECT 1683.910 202.450 1684.210 202.815 ;
        RECT 1682.975 202.150 1684.210 202.450 ;
        RECT 1682.975 202.135 1683.305 202.150 ;
        RECT 1924.935 202.135 1925.265 202.465 ;
        RECT 1635.135 201.455 1635.465 201.785 ;
        RECT 1924.950 201.105 1925.250 202.135 ;
        RECT 1538.535 200.775 1538.865 201.105 ;
        RECT 1924.935 200.775 1925.265 201.105 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1121.090 2604.300 1121.410 2604.360 ;
        RECT 1848.810 2604.300 1849.130 2604.360 ;
        RECT 1121.090 2604.160 1849.130 2604.300 ;
        RECT 1121.090 2604.100 1121.410 2604.160 ;
        RECT 1848.810 2604.100 1849.130 2604.160 ;
        RECT 1848.810 2552.960 1849.130 2553.020 ;
        RECT 2899.910 2552.960 2900.230 2553.020 ;
        RECT 1848.810 2552.820 2900.230 2552.960 ;
        RECT 1848.810 2552.760 1849.130 2552.820 ;
        RECT 2899.910 2552.760 2900.230 2552.820 ;
      LAYER via ;
        RECT 1121.120 2604.100 1121.380 2604.360 ;
        RECT 1848.840 2604.100 1849.100 2604.360 ;
        RECT 1848.840 2552.760 1849.100 2553.020 ;
        RECT 2899.940 2552.760 2900.200 2553.020 ;
      LAYER met2 ;
        RECT 1121.120 2604.070 1121.380 2604.390 ;
        RECT 1848.840 2604.070 1849.100 2604.390 ;
        RECT 1119.190 2599.370 1119.470 2600.000 ;
        RECT 1121.180 2599.370 1121.320 2604.070 ;
        RECT 1119.190 2599.230 1121.320 2599.370 ;
        RECT 1119.190 2596.000 1119.470 2599.230 ;
        RECT 1848.900 2553.050 1849.040 2604.070 ;
        RECT 1848.840 2552.730 1849.100 2553.050 ;
        RECT 2899.940 2552.730 2900.200 2553.050 ;
        RECT 2900.000 2551.885 2900.140 2552.730 ;
        RECT 2899.930 2551.515 2900.210 2551.885 ;
      LAYER via2 ;
        RECT 2899.930 2551.560 2900.210 2551.840 ;
      LAYER met3 ;
        RECT 2899.905 2551.850 2900.235 2551.865 ;
        RECT 2918.000 2551.850 2924.000 2552.300 ;
        RECT 2899.905 2551.550 2924.000 2551.850 ;
        RECT 2899.905 2551.535 2900.235 2551.550 ;
        RECT 2918.000 2551.100 2924.000 2551.550 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1145.010 2781.100 1145.330 2781.160 ;
        RECT 2899.450 2781.100 2899.770 2781.160 ;
        RECT 1145.010 2780.960 2899.770 2781.100 ;
        RECT 1145.010 2780.900 1145.330 2780.960 ;
        RECT 2899.450 2780.900 2899.770 2780.960 ;
      LAYER via ;
        RECT 1145.040 2780.900 1145.300 2781.160 ;
        RECT 2899.480 2780.900 2899.740 2781.160 ;
      LAYER met2 ;
        RECT 2899.470 2786.115 2899.750 2786.485 ;
        RECT 2899.540 2781.190 2899.680 2786.115 ;
        RECT 1145.040 2780.870 1145.300 2781.190 ;
        RECT 2899.480 2780.870 2899.740 2781.190 ;
        RECT 1144.490 2599.370 1144.770 2600.000 ;
        RECT 1145.100 2599.370 1145.240 2780.870 ;
        RECT 1144.490 2599.230 1145.240 2599.370 ;
        RECT 1144.490 2596.000 1144.770 2599.230 ;
      LAYER via2 ;
        RECT 2899.470 2786.160 2899.750 2786.440 ;
      LAYER met3 ;
        RECT 2899.445 2786.450 2899.775 2786.465 ;
        RECT 2918.000 2786.450 2924.000 2786.900 ;
        RECT 2899.445 2786.150 2924.000 2786.450 ;
        RECT 2899.445 2786.135 2899.775 2786.150 ;
        RECT 2918.000 2785.700 2924.000 2786.150 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1172.610 3015.700 1172.930 3015.760 ;
        RECT 2899.450 3015.700 2899.770 3015.760 ;
        RECT 1172.610 3015.560 2899.770 3015.700 ;
        RECT 1172.610 3015.500 1172.930 3015.560 ;
        RECT 2899.450 3015.500 2899.770 3015.560 ;
        RECT 1166.170 2632.520 1166.490 2632.580 ;
        RECT 1172.610 2632.520 1172.930 2632.580 ;
        RECT 1166.170 2632.380 1172.930 2632.520 ;
        RECT 1166.170 2632.320 1166.490 2632.380 ;
        RECT 1172.610 2632.320 1172.930 2632.380 ;
      LAYER via ;
        RECT 1172.640 3015.500 1172.900 3015.760 ;
        RECT 2899.480 3015.500 2899.740 3015.760 ;
        RECT 1166.200 2632.320 1166.460 2632.580 ;
        RECT 1172.640 2632.320 1172.900 2632.580 ;
      LAYER met2 ;
        RECT 2899.470 3020.715 2899.750 3021.085 ;
        RECT 2899.540 3015.790 2899.680 3020.715 ;
        RECT 1172.640 3015.470 1172.900 3015.790 ;
        RECT 2899.480 3015.470 2899.740 3015.790 ;
        RECT 1172.700 2632.610 1172.840 3015.470 ;
        RECT 1166.200 2632.290 1166.460 2632.610 ;
        RECT 1172.640 2632.290 1172.900 2632.610 ;
        RECT 1166.260 2599.370 1166.400 2632.290 ;
        RECT 1170.250 2599.370 1170.530 2600.000 ;
        RECT 1166.260 2599.230 1170.530 2599.370 ;
        RECT 1170.250 2596.000 1170.530 2599.230 ;
      LAYER via2 ;
        RECT 2899.470 3020.760 2899.750 3021.040 ;
      LAYER met3 ;
        RECT 2899.445 3021.050 2899.775 3021.065 ;
        RECT 2918.000 3021.050 2924.000 3021.500 ;
        RECT 2899.445 3020.750 2924.000 3021.050 ;
        RECT 2899.445 3020.735 2899.775 3020.750 ;
        RECT 2918.000 3020.300 2924.000 3020.750 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1200.210 3250.300 1200.530 3250.360 ;
        RECT 2899.450 3250.300 2899.770 3250.360 ;
        RECT 1200.210 3250.160 2899.770 3250.300 ;
        RECT 1200.210 3250.100 1200.530 3250.160 ;
        RECT 2899.450 3250.100 2899.770 3250.160 ;
      LAYER via ;
        RECT 1200.240 3250.100 1200.500 3250.360 ;
        RECT 2899.480 3250.100 2899.740 3250.360 ;
      LAYER met2 ;
        RECT 2899.470 3255.315 2899.750 3255.685 ;
        RECT 2899.540 3250.390 2899.680 3255.315 ;
        RECT 1200.240 3250.070 1200.500 3250.390 ;
        RECT 2899.480 3250.070 2899.740 3250.390 ;
        RECT 1200.300 2600.730 1200.440 3250.070 ;
        RECT 1198.000 2600.590 1200.440 2600.730 ;
        RECT 1196.010 2599.370 1196.290 2600.000 ;
        RECT 1198.000 2599.370 1198.140 2600.590 ;
        RECT 1196.010 2599.230 1198.140 2599.370 ;
        RECT 1196.010 2596.000 1196.290 2599.230 ;
      LAYER via2 ;
        RECT 2899.470 3255.360 2899.750 3255.640 ;
      LAYER met3 ;
        RECT 2899.445 3255.650 2899.775 3255.665 ;
        RECT 2918.000 3255.650 2924.000 3256.100 ;
        RECT 2899.445 3255.350 2924.000 3255.650 ;
        RECT 2899.445 3255.335 2899.775 3255.350 ;
        RECT 2918.000 3254.900 2924.000 3255.350 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1227.810 3484.900 1228.130 3484.960 ;
        RECT 2899.450 3484.900 2899.770 3484.960 ;
        RECT 1227.810 3484.760 2899.770 3484.900 ;
        RECT 1227.810 3484.700 1228.130 3484.760 ;
        RECT 2899.450 3484.700 2899.770 3484.760 ;
      LAYER via ;
        RECT 1227.840 3484.700 1228.100 3484.960 ;
        RECT 2899.480 3484.700 2899.740 3484.960 ;
      LAYER met2 ;
        RECT 2899.470 3489.915 2899.750 3490.285 ;
        RECT 2899.540 3484.990 2899.680 3489.915 ;
        RECT 1227.840 3484.670 1228.100 3484.990 ;
        RECT 2899.480 3484.670 2899.740 3484.990 ;
        RECT 1227.900 2600.730 1228.040 3484.670 ;
        RECT 1223.300 2600.590 1228.040 2600.730 ;
        RECT 1221.310 2599.370 1221.590 2600.000 ;
        RECT 1223.300 2599.370 1223.440 2600.590 ;
        RECT 1221.310 2599.230 1223.440 2599.370 ;
        RECT 1221.310 2596.000 1221.590 2599.230 ;
      LAYER via2 ;
        RECT 2899.470 3489.960 2899.750 3490.240 ;
      LAYER met3 ;
        RECT 2899.445 3490.250 2899.775 3490.265 ;
        RECT 2918.000 3490.250 2924.000 3490.700 ;
        RECT 2899.445 3489.950 2924.000 3490.250 ;
        RECT 2899.445 3489.935 2899.775 3489.950 ;
        RECT 2918.000 3489.500 2924.000 3489.950 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1248.510 3501.900 1248.830 3501.960 ;
        RECT 2635.870 3501.900 2636.190 3501.960 ;
        RECT 1248.510 3501.760 2636.190 3501.900 ;
        RECT 1248.510 3501.700 1248.830 3501.760 ;
        RECT 2635.870 3501.700 2636.190 3501.760 ;
      LAYER via ;
        RECT 1248.540 3501.700 1248.800 3501.960 ;
        RECT 2635.900 3501.700 2636.160 3501.960 ;
      LAYER met2 ;
        RECT 2635.750 3518.000 2636.310 3524.000 ;
        RECT 2635.960 3501.990 2636.100 3518.000 ;
        RECT 1248.540 3501.670 1248.800 3501.990 ;
        RECT 2635.900 3501.670 2636.160 3501.990 ;
        RECT 1247.070 2599.370 1247.350 2600.000 ;
        RECT 1248.600 2599.370 1248.740 3501.670 ;
        RECT 1247.070 2599.230 1248.740 2599.370 ;
        RECT 1247.070 2596.000 1247.350 2599.230 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1276.110 3503.600 1276.430 3503.660 ;
        RECT 2311.570 3503.600 2311.890 3503.660 ;
        RECT 1276.110 3503.460 2311.890 3503.600 ;
        RECT 1276.110 3503.400 1276.430 3503.460 ;
        RECT 2311.570 3503.400 2311.890 3503.460 ;
      LAYER via ;
        RECT 1276.140 3503.400 1276.400 3503.660 ;
        RECT 2311.600 3503.400 2311.860 3503.660 ;
      LAYER met2 ;
        RECT 2311.450 3518.000 2312.010 3524.000 ;
        RECT 2311.660 3503.690 2311.800 3518.000 ;
        RECT 1276.140 3503.370 1276.400 3503.690 ;
        RECT 2311.600 3503.370 2311.860 3503.690 ;
        RECT 1276.200 2600.730 1276.340 3503.370 ;
        RECT 1274.820 2600.590 1276.340 2600.730 ;
        RECT 1272.830 2599.370 1273.110 2600.000 ;
        RECT 1274.820 2599.370 1274.960 2600.590 ;
        RECT 1272.830 2599.230 1274.960 2599.370 ;
        RECT 1272.830 2596.000 1273.110 2599.230 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1303.710 3501.220 1304.030 3501.280 ;
        RECT 1987.270 3501.220 1987.590 3501.280 ;
        RECT 1303.710 3501.080 1987.590 3501.220 ;
        RECT 1303.710 3501.020 1304.030 3501.080 ;
        RECT 1987.270 3501.020 1987.590 3501.080 ;
      LAYER via ;
        RECT 1303.740 3501.020 1304.000 3501.280 ;
        RECT 1987.300 3501.020 1987.560 3501.280 ;
      LAYER met2 ;
        RECT 1987.150 3518.000 1987.710 3524.000 ;
        RECT 1987.360 3501.310 1987.500 3518.000 ;
        RECT 1303.740 3500.990 1304.000 3501.310 ;
        RECT 1987.300 3500.990 1987.560 3501.310 ;
        RECT 1303.800 2600.730 1303.940 3500.990 ;
        RECT 1300.580 2600.590 1303.940 2600.730 ;
        RECT 1298.590 2599.370 1298.870 2600.000 ;
        RECT 1300.580 2599.370 1300.720 2600.590 ;
        RECT 1298.590 2599.230 1300.720 2599.370 ;
        RECT 1298.590 2596.000 1298.870 2599.230 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1324.410 3499.520 1324.730 3499.580 ;
        RECT 1662.510 3499.520 1662.830 3499.580 ;
        RECT 1324.410 3499.380 1662.830 3499.520 ;
        RECT 1324.410 3499.320 1324.730 3499.380 ;
        RECT 1662.510 3499.320 1662.830 3499.380 ;
      LAYER via ;
        RECT 1324.440 3499.320 1324.700 3499.580 ;
        RECT 1662.540 3499.320 1662.800 3499.580 ;
      LAYER met2 ;
        RECT 1662.390 3518.000 1662.950 3524.000 ;
        RECT 1662.600 3499.610 1662.740 3518.000 ;
        RECT 1324.440 3499.290 1324.700 3499.610 ;
        RECT 1662.540 3499.290 1662.800 3499.610 ;
        RECT 1323.890 2599.370 1324.170 2600.000 ;
        RECT 1324.500 2599.370 1324.640 3499.290 ;
        RECT 1323.890 2599.230 1324.640 2599.370 ;
        RECT 1323.890 2596.000 1324.170 2599.230 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1346.105 3429.665 1346.275 3477.435 ;
        RECT 1346.105 3381.045 1346.275 3422.355 ;
        RECT 1347.025 3249.465 1347.195 3318.655 ;
        RECT 1345.645 2946.525 1345.815 2994.635 ;
        RECT 1346.105 2911.845 1346.275 2939.215 ;
      LAYER mcon ;
        RECT 1346.105 3477.265 1346.275 3477.435 ;
        RECT 1346.105 3422.185 1346.275 3422.355 ;
        RECT 1347.025 3318.485 1347.195 3318.655 ;
        RECT 1345.645 2994.465 1345.815 2994.635 ;
        RECT 1346.105 2939.045 1346.275 2939.215 ;
      LAYER met1 ;
        RECT 1338.210 3500.200 1338.530 3500.260 ;
        RECT 1345.570 3500.200 1345.890 3500.260 ;
        RECT 1338.210 3500.060 1345.890 3500.200 ;
        RECT 1338.210 3500.000 1338.530 3500.060 ;
        RECT 1345.570 3500.000 1345.890 3500.060 ;
        RECT 1346.045 3477.420 1346.335 3477.465 ;
        RECT 1346.490 3477.420 1346.810 3477.480 ;
        RECT 1346.045 3477.280 1346.810 3477.420 ;
        RECT 1346.045 3477.235 1346.335 3477.280 ;
        RECT 1346.490 3477.220 1346.810 3477.280 ;
        RECT 1346.030 3429.820 1346.350 3429.880 ;
        RECT 1345.835 3429.680 1346.350 3429.820 ;
        RECT 1346.030 3429.620 1346.350 3429.680 ;
        RECT 1346.030 3422.340 1346.350 3422.400 ;
        RECT 1345.835 3422.200 1346.350 3422.340 ;
        RECT 1346.030 3422.140 1346.350 3422.200 ;
        RECT 1346.045 3381.200 1346.335 3381.245 ;
        RECT 1346.490 3381.200 1346.810 3381.260 ;
        RECT 1346.045 3381.060 1346.810 3381.200 ;
        RECT 1346.045 3381.015 1346.335 3381.060 ;
        RECT 1346.490 3381.000 1346.810 3381.060 ;
        RECT 1346.490 3346.660 1346.810 3346.920 ;
        RECT 1346.580 3346.180 1346.720 3346.660 ;
        RECT 1346.950 3346.180 1347.270 3346.240 ;
        RECT 1346.580 3346.040 1347.270 3346.180 ;
        RECT 1346.950 3345.980 1347.270 3346.040 ;
        RECT 1346.950 3318.640 1347.270 3318.700 ;
        RECT 1346.755 3318.500 1347.270 3318.640 ;
        RECT 1346.950 3318.440 1347.270 3318.500 ;
        RECT 1346.950 3249.620 1347.270 3249.680 ;
        RECT 1346.755 3249.480 1347.270 3249.620 ;
        RECT 1346.950 3249.420 1347.270 3249.480 ;
        RECT 1346.950 3202.020 1347.270 3202.080 ;
        RECT 1346.580 3201.880 1347.270 3202.020 ;
        RECT 1346.580 3201.400 1346.720 3201.880 ;
        RECT 1346.950 3201.820 1347.270 3201.880 ;
        RECT 1346.490 3201.140 1346.810 3201.400 ;
        RECT 1346.490 3056.980 1346.810 3057.240 ;
        RECT 1346.580 3056.560 1346.720 3056.980 ;
        RECT 1346.490 3056.300 1346.810 3056.560 ;
        RECT 1345.570 3008.560 1345.890 3008.620 ;
        RECT 1346.490 3008.560 1346.810 3008.620 ;
        RECT 1345.570 3008.420 1346.810 3008.560 ;
        RECT 1345.570 3008.360 1345.890 3008.420 ;
        RECT 1346.490 3008.360 1346.810 3008.420 ;
        RECT 1345.570 2994.620 1345.890 2994.680 ;
        RECT 1345.375 2994.480 1345.890 2994.620 ;
        RECT 1345.570 2994.420 1345.890 2994.480 ;
        RECT 1345.585 2946.680 1345.875 2946.725 ;
        RECT 1346.030 2946.680 1346.350 2946.740 ;
        RECT 1345.585 2946.540 1346.350 2946.680 ;
        RECT 1345.585 2946.495 1345.875 2946.540 ;
        RECT 1346.030 2946.480 1346.350 2946.540 ;
        RECT 1346.030 2939.200 1346.350 2939.260 ;
        RECT 1345.835 2939.060 1346.350 2939.200 ;
        RECT 1346.030 2939.000 1346.350 2939.060 ;
        RECT 1346.045 2912.000 1346.335 2912.045 ;
        RECT 1346.490 2912.000 1346.810 2912.060 ;
        RECT 1346.045 2911.860 1346.810 2912.000 ;
        RECT 1346.045 2911.815 1346.335 2911.860 ;
        RECT 1346.490 2911.800 1346.810 2911.860 ;
        RECT 1345.570 2842.980 1345.890 2843.040 ;
        RECT 1346.950 2842.980 1347.270 2843.040 ;
        RECT 1345.570 2842.840 1347.270 2842.980 ;
        RECT 1345.570 2842.780 1345.890 2842.840 ;
        RECT 1346.950 2842.780 1347.270 2842.840 ;
        RECT 1346.950 2815.780 1347.270 2815.840 ;
        RECT 1346.580 2815.640 1347.270 2815.780 ;
        RECT 1346.580 2815.160 1346.720 2815.640 ;
        RECT 1346.950 2815.580 1347.270 2815.640 ;
        RECT 1346.490 2814.900 1346.810 2815.160 ;
        RECT 1346.030 2744.380 1346.350 2744.440 ;
        RECT 1347.410 2744.380 1347.730 2744.440 ;
        RECT 1346.030 2744.240 1347.730 2744.380 ;
        RECT 1346.030 2744.180 1346.350 2744.240 ;
        RECT 1347.410 2744.180 1347.730 2744.240 ;
        RECT 1346.490 2656.660 1346.810 2656.720 ;
        RECT 1347.870 2656.660 1348.190 2656.720 ;
        RECT 1346.490 2656.520 1348.190 2656.660 ;
        RECT 1346.490 2656.460 1346.810 2656.520 ;
        RECT 1347.870 2656.460 1348.190 2656.520 ;
      LAYER via ;
        RECT 1338.240 3500.000 1338.500 3500.260 ;
        RECT 1345.600 3500.000 1345.860 3500.260 ;
        RECT 1346.520 3477.220 1346.780 3477.480 ;
        RECT 1346.060 3429.620 1346.320 3429.880 ;
        RECT 1346.060 3422.140 1346.320 3422.400 ;
        RECT 1346.520 3381.000 1346.780 3381.260 ;
        RECT 1346.520 3346.660 1346.780 3346.920 ;
        RECT 1346.980 3345.980 1347.240 3346.240 ;
        RECT 1346.980 3318.440 1347.240 3318.700 ;
        RECT 1346.980 3249.420 1347.240 3249.680 ;
        RECT 1346.980 3201.820 1347.240 3202.080 ;
        RECT 1346.520 3201.140 1346.780 3201.400 ;
        RECT 1346.520 3056.980 1346.780 3057.240 ;
        RECT 1346.520 3056.300 1346.780 3056.560 ;
        RECT 1345.600 3008.360 1345.860 3008.620 ;
        RECT 1346.520 3008.360 1346.780 3008.620 ;
        RECT 1345.600 2994.420 1345.860 2994.680 ;
        RECT 1346.060 2946.480 1346.320 2946.740 ;
        RECT 1346.060 2939.000 1346.320 2939.260 ;
        RECT 1346.520 2911.800 1346.780 2912.060 ;
        RECT 1345.600 2842.780 1345.860 2843.040 ;
        RECT 1346.980 2842.780 1347.240 2843.040 ;
        RECT 1346.980 2815.580 1347.240 2815.840 ;
        RECT 1346.520 2814.900 1346.780 2815.160 ;
        RECT 1346.060 2744.180 1346.320 2744.440 ;
        RECT 1347.440 2744.180 1347.700 2744.440 ;
        RECT 1346.520 2656.460 1346.780 2656.720 ;
        RECT 1347.900 2656.460 1348.160 2656.720 ;
      LAYER met2 ;
        RECT 1338.090 3518.000 1338.650 3524.000 ;
        RECT 1338.300 3500.290 1338.440 3518.000 ;
        RECT 1338.240 3499.970 1338.500 3500.290 ;
        RECT 1345.600 3499.970 1345.860 3500.290 ;
        RECT 1345.660 3491.530 1345.800 3499.970 ;
        RECT 1345.660 3491.390 1346.720 3491.530 ;
        RECT 1346.580 3477.510 1346.720 3491.390 ;
        RECT 1346.520 3477.190 1346.780 3477.510 ;
        RECT 1346.060 3429.590 1346.320 3429.910 ;
        RECT 1346.120 3422.430 1346.260 3429.590 ;
        RECT 1346.060 3422.110 1346.320 3422.430 ;
        RECT 1346.520 3380.970 1346.780 3381.290 ;
        RECT 1346.580 3346.950 1346.720 3380.970 ;
        RECT 1346.520 3346.630 1346.780 3346.950 ;
        RECT 1346.980 3345.950 1347.240 3346.270 ;
        RECT 1347.040 3318.730 1347.180 3345.950 ;
        RECT 1346.980 3318.410 1347.240 3318.730 ;
        RECT 1346.980 3249.390 1347.240 3249.710 ;
        RECT 1347.040 3202.110 1347.180 3249.390 ;
        RECT 1346.980 3201.790 1347.240 3202.110 ;
        RECT 1346.520 3201.110 1346.780 3201.430 ;
        RECT 1346.580 3057.270 1346.720 3201.110 ;
        RECT 1346.520 3056.950 1346.780 3057.270 ;
        RECT 1346.520 3056.270 1346.780 3056.590 ;
        RECT 1346.580 3008.650 1346.720 3056.270 ;
        RECT 1345.600 3008.330 1345.860 3008.650 ;
        RECT 1346.520 3008.330 1346.780 3008.650 ;
        RECT 1345.660 2994.710 1345.800 3008.330 ;
        RECT 1345.600 2994.390 1345.860 2994.710 ;
        RECT 1346.060 2946.450 1346.320 2946.770 ;
        RECT 1346.120 2939.290 1346.260 2946.450 ;
        RECT 1346.060 2938.970 1346.320 2939.290 ;
        RECT 1346.520 2911.770 1346.780 2912.090 ;
        RECT 1346.580 2891.205 1346.720 2911.770 ;
        RECT 1345.590 2890.835 1345.870 2891.205 ;
        RECT 1346.510 2890.835 1346.790 2891.205 ;
        RECT 1345.660 2843.070 1345.800 2890.835 ;
        RECT 1345.600 2842.750 1345.860 2843.070 ;
        RECT 1346.980 2842.750 1347.240 2843.070 ;
        RECT 1347.040 2815.870 1347.180 2842.750 ;
        RECT 1346.980 2815.550 1347.240 2815.870 ;
        RECT 1346.520 2814.870 1346.780 2815.190 ;
        RECT 1346.580 2766.650 1346.720 2814.870 ;
        RECT 1346.120 2766.510 1346.720 2766.650 ;
        RECT 1346.120 2744.470 1346.260 2766.510 ;
        RECT 1346.060 2744.150 1346.320 2744.470 ;
        RECT 1347.440 2744.150 1347.700 2744.470 ;
        RECT 1347.500 2704.885 1347.640 2744.150 ;
        RECT 1346.510 2704.515 1346.790 2704.885 ;
        RECT 1347.430 2704.515 1347.710 2704.885 ;
        RECT 1346.580 2656.750 1346.720 2704.515 ;
        RECT 1346.520 2656.430 1346.780 2656.750 ;
        RECT 1347.900 2656.430 1348.160 2656.750 ;
        RECT 1347.960 2632.010 1348.100 2656.430 ;
        RECT 1347.040 2631.870 1348.100 2632.010 ;
        RECT 1347.040 2600.050 1347.180 2631.870 ;
        RECT 1347.040 2600.000 1349.870 2600.050 ;
        RECT 1347.040 2599.910 1349.930 2600.000 ;
        RECT 1349.650 2596.000 1349.930 2599.910 ;
      LAYER via2 ;
        RECT 1345.590 2890.880 1345.870 2891.160 ;
        RECT 1346.510 2890.880 1346.790 2891.160 ;
        RECT 1346.510 2704.560 1346.790 2704.840 ;
        RECT 1347.430 2704.560 1347.710 2704.840 ;
      LAYER met3 ;
        RECT 1345.565 2891.170 1345.895 2891.185 ;
        RECT 1346.485 2891.170 1346.815 2891.185 ;
        RECT 1345.565 2890.870 1346.815 2891.170 ;
        RECT 1345.565 2890.855 1345.895 2890.870 ;
        RECT 1346.485 2890.855 1346.815 2890.870 ;
        RECT 1346.485 2704.850 1346.815 2704.865 ;
        RECT 1347.405 2704.850 1347.735 2704.865 ;
        RECT 1346.485 2704.550 1347.735 2704.850 ;
        RECT 1346.485 2704.535 1346.815 2704.550 ;
        RECT 1347.405 2704.535 1347.735 2704.550 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 889.730 2609.315 890.010 2609.685 ;
        RECT 2902.230 2609.315 2902.510 2609.685 ;
        RECT 888.270 2599.370 888.550 2600.000 ;
        RECT 889.800 2599.370 889.940 2609.315 ;
        RECT 888.270 2599.230 889.940 2599.370 ;
        RECT 888.270 2596.000 888.550 2599.230 ;
        RECT 2902.300 439.805 2902.440 2609.315 ;
        RECT 2902.230 439.435 2902.510 439.805 ;
      LAYER via2 ;
        RECT 889.730 2609.360 890.010 2609.640 ;
        RECT 2902.230 2609.360 2902.510 2609.640 ;
        RECT 2902.230 439.480 2902.510 439.760 ;
      LAYER met3 ;
        RECT 889.705 2609.650 890.035 2609.665 ;
        RECT 2902.205 2609.650 2902.535 2609.665 ;
        RECT 889.705 2609.350 2902.535 2609.650 ;
        RECT 889.705 2609.335 890.035 2609.350 ;
        RECT 2902.205 2609.335 2902.535 2609.350 ;
        RECT 2902.205 439.770 2902.535 439.785 ;
        RECT 2918.000 439.770 2924.000 440.220 ;
        RECT 2902.205 439.470 2924.000 439.770 ;
        RECT 2902.205 439.455 2902.535 439.470 ;
        RECT 2918.000 439.020 2924.000 439.470 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1013.910 3499.860 1014.230 3499.920 ;
        RECT 1373.170 3499.860 1373.490 3499.920 ;
        RECT 1013.910 3499.720 1373.490 3499.860 ;
        RECT 1013.910 3499.660 1014.230 3499.720 ;
        RECT 1373.170 3499.660 1373.490 3499.720 ;
      LAYER via ;
        RECT 1013.940 3499.660 1014.200 3499.920 ;
        RECT 1373.200 3499.660 1373.460 3499.920 ;
      LAYER met2 ;
        RECT 1013.790 3518.000 1014.350 3524.000 ;
        RECT 1014.000 3499.950 1014.140 3518.000 ;
        RECT 1013.940 3499.630 1014.200 3499.950 ;
        RECT 1373.200 3499.630 1373.460 3499.950 ;
        RECT 1373.260 2600.050 1373.400 3499.630 ;
        RECT 1373.260 2600.000 1375.630 2600.050 ;
        RECT 1373.260 2599.910 1375.690 2600.000 ;
        RECT 1375.410 2596.000 1375.690 2599.910 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 689.150 3504.960 689.470 3505.020 ;
        RECT 1400.770 3504.960 1401.090 3505.020 ;
        RECT 689.150 3504.820 1401.090 3504.960 ;
        RECT 689.150 3504.760 689.470 3504.820 ;
        RECT 1400.770 3504.760 1401.090 3504.820 ;
      LAYER via ;
        RECT 689.180 3504.760 689.440 3505.020 ;
        RECT 1400.800 3504.760 1401.060 3505.020 ;
      LAYER met2 ;
        RECT 689.030 3518.000 689.590 3524.000 ;
        RECT 689.240 3505.050 689.380 3518.000 ;
        RECT 689.180 3504.730 689.440 3505.050 ;
        RECT 1400.800 3504.730 1401.060 3505.050 ;
        RECT 1400.860 2600.050 1401.000 3504.730 ;
        RECT 1400.860 2600.000 1401.390 2600.050 ;
        RECT 1400.860 2599.910 1401.450 2600.000 ;
        RECT 1401.170 2596.000 1401.450 2599.910 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 364.850 3503.260 365.170 3503.320 ;
        RECT 1421.470 3503.260 1421.790 3503.320 ;
        RECT 364.850 3503.120 1421.790 3503.260 ;
        RECT 364.850 3503.060 365.170 3503.120 ;
        RECT 1421.470 3503.060 1421.790 3503.120 ;
      LAYER via ;
        RECT 364.880 3503.060 365.140 3503.320 ;
        RECT 1421.500 3503.060 1421.760 3503.320 ;
      LAYER met2 ;
        RECT 364.730 3518.000 365.290 3524.000 ;
        RECT 364.940 3503.350 365.080 3518.000 ;
        RECT 364.880 3503.030 365.140 3503.350 ;
        RECT 1421.500 3503.030 1421.760 3503.350 ;
        RECT 1421.560 2600.730 1421.700 3503.030 ;
        RECT 1421.560 2600.590 1424.920 2600.730 ;
        RECT 1424.780 2600.050 1424.920 2600.590 ;
        RECT 1424.780 2600.000 1426.690 2600.050 ;
        RECT 1424.780 2599.910 1426.750 2600.000 ;
        RECT 1426.470 2596.000 1426.750 2599.910 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1449.605 3442.925 1449.775 3477.435 ;
        RECT 1449.145 3284.485 1449.315 3332.595 ;
        RECT 1449.145 3187.925 1449.315 3236.035 ;
        RECT 1449.605 3091.365 1449.775 3139.475 ;
      LAYER mcon ;
        RECT 1449.605 3477.265 1449.775 3477.435 ;
        RECT 1449.145 3332.425 1449.315 3332.595 ;
        RECT 1449.145 3235.865 1449.315 3236.035 ;
        RECT 1449.605 3139.305 1449.775 3139.475 ;
      LAYER met1 ;
        RECT 40.550 3501.560 40.870 3501.620 ;
        RECT 1449.990 3501.560 1450.310 3501.620 ;
        RECT 40.550 3501.420 1450.310 3501.560 ;
        RECT 40.550 3501.360 40.870 3501.420 ;
        RECT 1449.990 3501.360 1450.310 3501.420 ;
        RECT 1449.545 3477.420 1449.835 3477.465 ;
        RECT 1449.990 3477.420 1450.310 3477.480 ;
        RECT 1449.545 3477.280 1450.310 3477.420 ;
        RECT 1449.545 3477.235 1449.835 3477.280 ;
        RECT 1449.990 3477.220 1450.310 3477.280 ;
        RECT 1449.530 3443.080 1449.850 3443.140 ;
        RECT 1449.335 3442.940 1449.850 3443.080 ;
        RECT 1449.530 3442.880 1449.850 3442.940 ;
        RECT 1449.070 3332.580 1449.390 3332.640 ;
        RECT 1449.070 3332.440 1449.585 3332.580 ;
        RECT 1449.070 3332.380 1449.390 3332.440 ;
        RECT 1449.070 3284.640 1449.390 3284.700 ;
        RECT 1449.070 3284.500 1449.585 3284.640 ;
        RECT 1449.070 3284.440 1449.390 3284.500 ;
        RECT 1449.070 3236.020 1449.390 3236.080 ;
        RECT 1449.070 3235.880 1449.585 3236.020 ;
        RECT 1449.070 3235.820 1449.390 3235.880 ;
        RECT 1449.070 3188.080 1449.390 3188.140 ;
        RECT 1449.070 3187.940 1449.585 3188.080 ;
        RECT 1449.070 3187.880 1449.390 3187.940 ;
        RECT 1449.530 3139.460 1449.850 3139.520 ;
        RECT 1449.335 3139.320 1449.850 3139.460 ;
        RECT 1449.530 3139.260 1449.850 3139.320 ;
        RECT 1449.545 3091.520 1449.835 3091.565 ;
        RECT 1449.990 3091.520 1450.310 3091.580 ;
        RECT 1449.545 3091.380 1450.310 3091.520 ;
        RECT 1449.545 3091.335 1449.835 3091.380 ;
        RECT 1449.990 3091.320 1450.310 3091.380 ;
        RECT 1449.070 3056.840 1449.390 3056.900 ;
        RECT 1449.990 3056.840 1450.310 3056.900 ;
        RECT 1449.070 3056.700 1450.310 3056.840 ;
        RECT 1449.070 3056.640 1449.390 3056.700 ;
        RECT 1449.990 3056.640 1450.310 3056.700 ;
        RECT 1449.070 2863.720 1449.390 2863.780 ;
        RECT 1449.990 2863.720 1450.310 2863.780 ;
        RECT 1449.070 2863.580 1450.310 2863.720 ;
        RECT 1449.070 2863.520 1449.390 2863.580 ;
        RECT 1449.990 2863.520 1450.310 2863.580 ;
        RECT 1449.070 2767.160 1449.390 2767.220 ;
        RECT 1449.990 2767.160 1450.310 2767.220 ;
        RECT 1449.070 2767.020 1450.310 2767.160 ;
        RECT 1449.070 2766.960 1449.390 2767.020 ;
        RECT 1449.990 2766.960 1450.310 2767.020 ;
      LAYER via ;
        RECT 40.580 3501.360 40.840 3501.620 ;
        RECT 1450.020 3501.360 1450.280 3501.620 ;
        RECT 1450.020 3477.220 1450.280 3477.480 ;
        RECT 1449.560 3442.880 1449.820 3443.140 ;
        RECT 1449.100 3332.380 1449.360 3332.640 ;
        RECT 1449.100 3284.440 1449.360 3284.700 ;
        RECT 1449.100 3235.820 1449.360 3236.080 ;
        RECT 1449.100 3187.880 1449.360 3188.140 ;
        RECT 1449.560 3139.260 1449.820 3139.520 ;
        RECT 1450.020 3091.320 1450.280 3091.580 ;
        RECT 1449.100 3056.640 1449.360 3056.900 ;
        RECT 1450.020 3056.640 1450.280 3056.900 ;
        RECT 1449.100 2863.520 1449.360 2863.780 ;
        RECT 1450.020 2863.520 1450.280 2863.780 ;
        RECT 1449.100 2766.960 1449.360 2767.220 ;
        RECT 1450.020 2766.960 1450.280 2767.220 ;
      LAYER met2 ;
        RECT 40.430 3518.000 40.990 3524.000 ;
        RECT 40.640 3501.650 40.780 3518.000 ;
        RECT 40.580 3501.330 40.840 3501.650 ;
        RECT 1450.020 3501.330 1450.280 3501.650 ;
        RECT 1450.080 3477.510 1450.220 3501.330 ;
        RECT 1450.020 3477.190 1450.280 3477.510 ;
        RECT 1449.560 3442.850 1449.820 3443.170 ;
        RECT 1449.620 3394.970 1449.760 3442.850 ;
        RECT 1449.620 3394.830 1450.220 3394.970 ;
        RECT 1450.080 3346.690 1450.220 3394.830 ;
        RECT 1449.160 3346.550 1450.220 3346.690 ;
        RECT 1449.160 3332.670 1449.300 3346.550 ;
        RECT 1449.100 3332.350 1449.360 3332.670 ;
        RECT 1449.100 3284.410 1449.360 3284.730 ;
        RECT 1449.160 3236.110 1449.300 3284.410 ;
        RECT 1449.100 3235.790 1449.360 3236.110 ;
        RECT 1449.100 3187.850 1449.360 3188.170 ;
        RECT 1449.160 3152.890 1449.300 3187.850 ;
        RECT 1449.160 3152.750 1449.760 3152.890 ;
        RECT 1449.620 3139.550 1449.760 3152.750 ;
        RECT 1449.560 3139.230 1449.820 3139.550 ;
        RECT 1450.020 3091.290 1450.280 3091.610 ;
        RECT 1450.080 3056.930 1450.220 3091.290 ;
        RECT 1449.100 3056.610 1449.360 3056.930 ;
        RECT 1450.020 3056.610 1450.280 3056.930 ;
        RECT 1449.160 2959.770 1449.300 3056.610 ;
        RECT 1449.160 2959.630 1450.220 2959.770 ;
        RECT 1450.080 2863.810 1450.220 2959.630 ;
        RECT 1449.100 2863.490 1449.360 2863.810 ;
        RECT 1450.020 2863.490 1450.280 2863.810 ;
        RECT 1449.160 2863.210 1449.300 2863.490 ;
        RECT 1449.160 2863.070 1449.760 2863.210 ;
        RECT 1449.620 2815.610 1449.760 2863.070 ;
        RECT 1449.620 2815.470 1450.220 2815.610 ;
        RECT 1450.080 2767.250 1450.220 2815.470 ;
        RECT 1449.100 2766.930 1449.360 2767.250 ;
        RECT 1450.020 2766.930 1450.280 2767.250 ;
        RECT 1449.160 2718.370 1449.300 2766.930 ;
        RECT 1449.160 2718.230 1449.760 2718.370 ;
        RECT 1449.620 2670.770 1449.760 2718.230 ;
        RECT 1449.620 2670.630 1450.220 2670.770 ;
        RECT 1450.080 2600.050 1450.220 2670.630 ;
        RECT 1450.080 2600.000 1452.450 2600.050 ;
        RECT 1450.080 2599.910 1452.510 2600.000 ;
        RECT 1452.230 2596.000 1452.510 2599.910 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.250 3263.900 15.570 3263.960 ;
        RECT 1476.670 3263.900 1476.990 3263.960 ;
        RECT 15.250 3263.760 1476.990 3263.900 ;
        RECT 15.250 3263.700 15.570 3263.760 ;
        RECT 1476.670 3263.700 1476.990 3263.760 ;
      LAYER via ;
        RECT 15.280 3263.700 15.540 3263.960 ;
        RECT 1476.700 3263.700 1476.960 3263.960 ;
      LAYER met2 ;
        RECT 15.270 3267.555 15.550 3267.925 ;
        RECT 15.340 3263.990 15.480 3267.555 ;
        RECT 15.280 3263.670 15.540 3263.990 ;
        RECT 1476.700 3263.670 1476.960 3263.990 ;
        RECT 1476.760 2600.050 1476.900 3263.670 ;
        RECT 1476.760 2600.000 1478.210 2600.050 ;
        RECT 1476.760 2599.910 1478.270 2600.000 ;
        RECT 1477.990 2596.000 1478.270 2599.910 ;
      LAYER via2 ;
        RECT 15.270 3267.600 15.550 3267.880 ;
      LAYER met3 ;
        RECT -4.000 3267.890 2.000 3268.340 ;
        RECT 15.245 3267.890 15.575 3267.905 ;
        RECT -4.000 3267.590 15.575 3267.890 ;
        RECT -4.000 3267.140 2.000 3267.590 ;
        RECT 15.245 3267.575 15.575 3267.590 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.170 2974.220 16.490 2974.280 ;
        RECT 1497.830 2974.220 1498.150 2974.280 ;
        RECT 16.170 2974.080 1498.150 2974.220 ;
        RECT 16.170 2974.020 16.490 2974.080 ;
        RECT 1497.830 2974.020 1498.150 2974.080 ;
      LAYER via ;
        RECT 16.200 2974.020 16.460 2974.280 ;
        RECT 1497.860 2974.020 1498.120 2974.280 ;
      LAYER met2 ;
        RECT 16.190 2979.915 16.470 2980.285 ;
        RECT 16.260 2974.310 16.400 2979.915 ;
        RECT 16.200 2973.990 16.460 2974.310 ;
        RECT 1497.860 2973.990 1498.120 2974.310 ;
        RECT 1497.920 2601.410 1498.060 2973.990 ;
        RECT 1497.920 2601.270 1502.200 2601.410 ;
        RECT 1502.060 2600.050 1502.200 2601.270 ;
        RECT 1502.060 2600.000 1503.970 2600.050 ;
        RECT 1502.060 2599.910 1504.030 2600.000 ;
        RECT 1503.750 2596.000 1504.030 2599.910 ;
      LAYER via2 ;
        RECT 16.190 2979.960 16.470 2980.240 ;
      LAYER met3 ;
        RECT -4.000 2980.250 2.000 2980.700 ;
        RECT 16.165 2980.250 16.495 2980.265 ;
        RECT -4.000 2979.950 16.495 2980.250 ;
        RECT -4.000 2979.500 2.000 2979.950 ;
        RECT 16.165 2979.935 16.495 2979.950 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 2691.340 17.410 2691.400 ;
        RECT 1524.970 2691.340 1525.290 2691.400 ;
        RECT 17.090 2691.200 1525.290 2691.340 ;
        RECT 17.090 2691.140 17.410 2691.200 ;
        RECT 1524.970 2691.140 1525.290 2691.200 ;
      LAYER via ;
        RECT 17.120 2691.140 17.380 2691.400 ;
        RECT 1525.000 2691.140 1525.260 2691.400 ;
      LAYER met2 ;
        RECT 17.110 2692.955 17.390 2693.325 ;
        RECT 17.180 2691.430 17.320 2692.955 ;
        RECT 17.120 2691.110 17.380 2691.430 ;
        RECT 1525.000 2691.110 1525.260 2691.430 ;
        RECT 1525.060 2600.730 1525.200 2691.110 ;
        RECT 1525.060 2600.590 1526.120 2600.730 ;
        RECT 1525.980 2600.050 1526.120 2600.590 ;
        RECT 1525.980 2600.000 1529.270 2600.050 ;
        RECT 1525.980 2599.910 1529.330 2600.000 ;
        RECT 1529.050 2596.000 1529.330 2599.910 ;
      LAYER via2 ;
        RECT 17.110 2693.000 17.390 2693.280 ;
      LAYER met3 ;
        RECT -4.000 2693.290 2.000 2693.740 ;
        RECT 17.085 2693.290 17.415 2693.305 ;
        RECT -4.000 2692.990 17.415 2693.290 ;
        RECT -4.000 2692.540 2.000 2692.990 ;
        RECT 17.085 2692.975 17.415 2692.990 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.250 2613.140 15.570 2613.200 ;
        RECT 1553.030 2613.140 1553.350 2613.200 ;
        RECT 15.250 2613.000 1553.350 2613.140 ;
        RECT 15.250 2612.940 15.570 2613.000 ;
        RECT 1553.030 2612.940 1553.350 2613.000 ;
      LAYER via ;
        RECT 15.280 2612.940 15.540 2613.200 ;
        RECT 1553.060 2612.940 1553.320 2613.200 ;
      LAYER met2 ;
        RECT 15.280 2612.910 15.540 2613.230 ;
        RECT 1553.060 2612.910 1553.320 2613.230 ;
        RECT 15.340 2405.685 15.480 2612.910 ;
        RECT 1553.120 2600.050 1553.260 2612.910 ;
        RECT 1553.120 2600.000 1555.030 2600.050 ;
        RECT 1553.120 2599.910 1555.090 2600.000 ;
        RECT 1554.810 2596.000 1555.090 2599.910 ;
        RECT 15.270 2405.315 15.550 2405.685 ;
      LAYER via2 ;
        RECT 15.270 2405.360 15.550 2405.640 ;
      LAYER met3 ;
        RECT -4.000 2405.650 2.000 2406.100 ;
        RECT 15.245 2405.650 15.575 2405.665 ;
        RECT -4.000 2405.350 15.575 2405.650 ;
        RECT -4.000 2404.900 2.000 2405.350 ;
        RECT 15.245 2405.335 15.575 2405.350 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 254.910 2589.340 255.230 2589.400 ;
        RECT 289.410 2589.340 289.730 2589.400 ;
        RECT 254.910 2589.200 289.730 2589.340 ;
        RECT 254.910 2589.140 255.230 2589.200 ;
        RECT 289.410 2589.140 289.730 2589.200 ;
        RECT 351.510 2589.340 351.830 2589.400 ;
        RECT 386.010 2589.340 386.330 2589.400 ;
        RECT 351.510 2589.200 386.330 2589.340 ;
        RECT 351.510 2589.140 351.830 2589.200 ;
        RECT 386.010 2589.140 386.330 2589.200 ;
        RECT 448.110 2589.340 448.430 2589.400 ;
        RECT 482.610 2589.340 482.930 2589.400 ;
        RECT 448.110 2589.200 482.930 2589.340 ;
        RECT 448.110 2589.140 448.430 2589.200 ;
        RECT 482.610 2589.140 482.930 2589.200 ;
        RECT 544.710 2589.340 545.030 2589.400 ;
        RECT 579.210 2589.340 579.530 2589.400 ;
        RECT 544.710 2589.200 579.530 2589.340 ;
        RECT 544.710 2589.140 545.030 2589.200 ;
        RECT 579.210 2589.140 579.530 2589.200 ;
        RECT 641.310 2589.340 641.630 2589.400 ;
        RECT 675.810 2589.340 676.130 2589.400 ;
        RECT 641.310 2589.200 676.130 2589.340 ;
        RECT 641.310 2589.140 641.630 2589.200 ;
        RECT 675.810 2589.140 676.130 2589.200 ;
        RECT 737.910 2589.340 738.230 2589.400 ;
        RECT 772.410 2589.340 772.730 2589.400 ;
        RECT 737.910 2589.200 772.730 2589.340 ;
        RECT 737.910 2589.140 738.230 2589.200 ;
        RECT 772.410 2589.140 772.730 2589.200 ;
        RECT 138.070 2587.980 138.390 2588.040 ;
        RECT 185.910 2587.980 186.230 2588.040 ;
        RECT 138.070 2587.840 186.230 2587.980 ;
        RECT 138.070 2587.780 138.390 2587.840 ;
        RECT 185.910 2587.780 186.230 2587.840 ;
        RECT 15.710 2120.480 16.030 2120.540 ;
        RECT 31.350 2120.480 31.670 2120.540 ;
        RECT 15.710 2120.340 31.670 2120.480 ;
        RECT 15.710 2120.280 16.030 2120.340 ;
        RECT 31.350 2120.280 31.670 2120.340 ;
      LAYER via ;
        RECT 254.940 2589.140 255.200 2589.400 ;
        RECT 289.440 2589.140 289.700 2589.400 ;
        RECT 351.540 2589.140 351.800 2589.400 ;
        RECT 386.040 2589.140 386.300 2589.400 ;
        RECT 448.140 2589.140 448.400 2589.400 ;
        RECT 482.640 2589.140 482.900 2589.400 ;
        RECT 544.740 2589.140 545.000 2589.400 ;
        RECT 579.240 2589.140 579.500 2589.400 ;
        RECT 641.340 2589.140 641.600 2589.400 ;
        RECT 675.840 2589.140 676.100 2589.400 ;
        RECT 737.940 2589.140 738.200 2589.400 ;
        RECT 772.440 2589.140 772.700 2589.400 ;
        RECT 138.100 2587.780 138.360 2588.040 ;
        RECT 185.940 2587.780 186.200 2588.040 ;
        RECT 15.740 2120.280 16.000 2120.540 ;
        RECT 31.380 2120.280 31.640 2120.540 ;
      LAYER met2 ;
        RECT 1578.810 2596.650 1579.090 2596.765 ;
        RECT 1580.570 2596.650 1580.850 2600.000 ;
        RECT 1578.810 2596.510 1580.850 2596.650 ;
        RECT 1578.810 2596.395 1579.090 2596.510 ;
        RECT 1580.570 2596.000 1580.850 2596.510 ;
        RECT 185.930 2589.595 186.210 2589.965 ;
        RECT 289.430 2589.595 289.710 2589.965 ;
        RECT 386.030 2589.595 386.310 2589.965 ;
        RECT 482.630 2589.595 482.910 2589.965 ;
        RECT 579.230 2589.595 579.510 2589.965 ;
        RECT 675.830 2589.595 676.110 2589.965 ;
        RECT 772.430 2589.595 772.710 2589.965 ;
        RECT 834.990 2589.595 835.270 2589.965 ;
        RECT 62.650 2588.490 62.930 2588.605 ;
        RECT 61.800 2588.350 62.930 2588.490 ;
        RECT 61.800 2587.925 61.940 2588.350 ;
        RECT 62.650 2588.235 62.930 2588.350 ;
        RECT 110.030 2588.490 110.310 2588.605 ;
        RECT 110.030 2588.350 111.160 2588.490 ;
        RECT 110.030 2588.235 110.310 2588.350 ;
        RECT 111.020 2587.925 111.160 2588.350 ;
        RECT 186.000 2588.070 186.140 2589.595 ;
        RECT 289.500 2589.430 289.640 2589.595 ;
        RECT 386.100 2589.430 386.240 2589.595 ;
        RECT 482.700 2589.430 482.840 2589.595 ;
        RECT 579.300 2589.430 579.440 2589.595 ;
        RECT 675.900 2589.430 676.040 2589.595 ;
        RECT 772.500 2589.430 772.640 2589.595 ;
        RECT 254.940 2589.285 255.200 2589.430 ;
        RECT 254.930 2588.915 255.210 2589.285 ;
        RECT 289.440 2589.110 289.700 2589.430 ;
        RECT 351.540 2589.285 351.800 2589.430 ;
        RECT 351.530 2588.915 351.810 2589.285 ;
        RECT 386.040 2589.110 386.300 2589.430 ;
        RECT 448.140 2589.285 448.400 2589.430 ;
        RECT 448.130 2588.915 448.410 2589.285 ;
        RECT 482.640 2589.110 482.900 2589.430 ;
        RECT 544.740 2589.285 545.000 2589.430 ;
        RECT 544.730 2588.915 545.010 2589.285 ;
        RECT 579.240 2589.110 579.500 2589.430 ;
        RECT 641.340 2589.285 641.600 2589.430 ;
        RECT 641.330 2588.915 641.610 2589.285 ;
        RECT 675.840 2589.110 676.100 2589.430 ;
        RECT 737.940 2589.285 738.200 2589.430 ;
        RECT 737.930 2588.915 738.210 2589.285 ;
        RECT 772.440 2589.110 772.700 2589.430 ;
        RECT 834.530 2589.170 834.810 2589.285 ;
        RECT 835.060 2589.170 835.200 2589.595 ;
        RECT 834.530 2589.030 835.200 2589.170 ;
        RECT 834.530 2588.915 834.810 2589.030 ;
        RECT 138.100 2587.925 138.360 2588.070 ;
        RECT 31.370 2587.555 31.650 2587.925 ;
        RECT 61.730 2587.555 62.010 2587.925 ;
        RECT 110.950 2587.555 111.230 2587.925 ;
        RECT 138.090 2587.555 138.370 2587.925 ;
        RECT 185.940 2587.750 186.200 2588.070 ;
        RECT 31.440 2120.570 31.580 2587.555 ;
        RECT 15.740 2120.250 16.000 2120.570 ;
        RECT 31.380 2120.250 31.640 2120.570 ;
        RECT 15.800 2118.725 15.940 2120.250 ;
        RECT 15.730 2118.355 16.010 2118.725 ;
      LAYER via2 ;
        RECT 1578.810 2596.440 1579.090 2596.720 ;
        RECT 185.930 2589.640 186.210 2589.920 ;
        RECT 289.430 2589.640 289.710 2589.920 ;
        RECT 386.030 2589.640 386.310 2589.920 ;
        RECT 482.630 2589.640 482.910 2589.920 ;
        RECT 579.230 2589.640 579.510 2589.920 ;
        RECT 675.830 2589.640 676.110 2589.920 ;
        RECT 772.430 2589.640 772.710 2589.920 ;
        RECT 834.990 2589.640 835.270 2589.920 ;
        RECT 62.650 2588.280 62.930 2588.560 ;
        RECT 110.030 2588.280 110.310 2588.560 ;
        RECT 254.930 2588.960 255.210 2589.240 ;
        RECT 351.530 2588.960 351.810 2589.240 ;
        RECT 448.130 2588.960 448.410 2589.240 ;
        RECT 544.730 2588.960 545.010 2589.240 ;
        RECT 641.330 2588.960 641.610 2589.240 ;
        RECT 737.930 2588.960 738.210 2589.240 ;
        RECT 834.530 2588.960 834.810 2589.240 ;
        RECT 31.370 2587.600 31.650 2587.880 ;
        RECT 61.730 2587.600 62.010 2587.880 ;
        RECT 110.950 2587.600 111.230 2587.880 ;
        RECT 138.090 2587.600 138.370 2587.880 ;
        RECT 15.730 2118.400 16.010 2118.680 ;
      LAYER met3 ;
        RECT 1563.350 2596.730 1563.730 2596.740 ;
        RECT 1578.785 2596.730 1579.115 2596.745 ;
        RECT 1563.350 2596.430 1579.115 2596.730 ;
        RECT 1563.350 2596.420 1563.730 2596.430 ;
        RECT 1578.785 2596.415 1579.115 2596.430 ;
        RECT 1513.670 2594.690 1514.050 2594.700 ;
        RECT 1563.350 2594.690 1563.730 2594.700 ;
        RECT 1513.670 2594.390 1563.730 2594.690 ;
        RECT 1513.670 2594.380 1514.050 2594.390 ;
        RECT 1563.350 2594.380 1563.730 2594.390 ;
        RECT 911.070 2592.650 911.450 2592.660 ;
        RECT 911.070 2592.350 958.330 2592.650 ;
        RECT 911.070 2592.340 911.450 2592.350 ;
        RECT 185.905 2589.930 186.235 2589.945 ;
        RECT 289.405 2589.930 289.735 2589.945 ;
        RECT 386.005 2589.930 386.335 2589.945 ;
        RECT 482.605 2589.930 482.935 2589.945 ;
        RECT 579.205 2589.930 579.535 2589.945 ;
        RECT 675.805 2589.930 676.135 2589.945 ;
        RECT 772.405 2589.930 772.735 2589.945 ;
        RECT 834.965 2589.930 835.295 2589.945 ;
        RECT 882.550 2589.930 882.930 2589.940 ;
        RECT 185.905 2589.630 207.610 2589.930 ;
        RECT 185.905 2589.615 186.235 2589.630 ;
        RECT 207.310 2589.250 207.610 2589.630 ;
        RECT 289.405 2589.630 304.210 2589.930 ;
        RECT 289.405 2589.615 289.735 2589.630 ;
        RECT 254.905 2589.250 255.235 2589.265 ;
        RECT 207.310 2588.950 255.235 2589.250 ;
        RECT 303.910 2589.250 304.210 2589.630 ;
        RECT 386.005 2589.630 400.810 2589.930 ;
        RECT 386.005 2589.615 386.335 2589.630 ;
        RECT 351.505 2589.250 351.835 2589.265 ;
        RECT 303.910 2588.950 351.835 2589.250 ;
        RECT 400.510 2589.250 400.810 2589.630 ;
        RECT 482.605 2589.630 497.410 2589.930 ;
        RECT 482.605 2589.615 482.935 2589.630 ;
        RECT 448.105 2589.250 448.435 2589.265 ;
        RECT 400.510 2588.950 448.435 2589.250 ;
        RECT 497.110 2589.250 497.410 2589.630 ;
        RECT 579.205 2589.630 594.010 2589.930 ;
        RECT 579.205 2589.615 579.535 2589.630 ;
        RECT 544.705 2589.250 545.035 2589.265 ;
        RECT 497.110 2588.950 545.035 2589.250 ;
        RECT 593.710 2589.250 594.010 2589.630 ;
        RECT 675.805 2589.630 690.610 2589.930 ;
        RECT 675.805 2589.615 676.135 2589.630 ;
        RECT 641.305 2589.250 641.635 2589.265 ;
        RECT 593.710 2588.950 641.635 2589.250 ;
        RECT 690.310 2589.250 690.610 2589.630 ;
        RECT 772.405 2589.630 787.210 2589.930 ;
        RECT 772.405 2589.615 772.735 2589.630 ;
        RECT 737.905 2589.250 738.235 2589.265 ;
        RECT 690.310 2588.950 738.235 2589.250 ;
        RECT 786.910 2589.250 787.210 2589.630 ;
        RECT 834.965 2589.630 882.930 2589.930 ;
        RECT 834.965 2589.615 835.295 2589.630 ;
        RECT 882.550 2589.620 882.930 2589.630 ;
        RECT 883.470 2589.930 883.850 2589.940 ;
        RECT 883.470 2589.630 910.490 2589.930 ;
        RECT 883.470 2589.620 883.850 2589.630 ;
        RECT 834.505 2589.250 834.835 2589.265 ;
        RECT 786.910 2588.950 834.835 2589.250 ;
        RECT 910.190 2589.250 910.490 2589.630 ;
        RECT 911.070 2589.620 911.450 2589.940 ;
        RECT 911.110 2589.250 911.410 2589.620 ;
        RECT 910.190 2588.950 911.410 2589.250 ;
        RECT 958.030 2589.250 958.330 2592.350 ;
        RECT 980.070 2589.930 980.450 2589.940 ;
        RECT 1051.830 2589.930 1052.210 2589.940 ;
        RECT 980.070 2589.630 1052.210 2589.930 ;
        RECT 980.070 2589.620 980.450 2589.630 ;
        RECT 1051.830 2589.620 1052.210 2589.630 ;
        RECT 1095.990 2589.930 1096.370 2589.940 ;
        RECT 1172.350 2589.930 1172.730 2589.940 ;
        RECT 1095.990 2589.630 1172.730 2589.930 ;
        RECT 1095.990 2589.620 1096.370 2589.630 ;
        RECT 1172.350 2589.620 1172.730 2589.630 ;
        RECT 1218.350 2589.930 1218.730 2589.940 ;
        RECT 1221.110 2589.930 1221.490 2589.940 ;
        RECT 1218.350 2589.630 1221.490 2589.930 ;
        RECT 1218.350 2589.620 1218.730 2589.630 ;
        RECT 1221.110 2589.620 1221.490 2589.630 ;
        RECT 1270.790 2589.930 1271.170 2589.940 ;
        RECT 1322.310 2589.930 1322.690 2589.940 ;
        RECT 1270.790 2589.630 1322.690 2589.930 ;
        RECT 1270.790 2589.620 1271.170 2589.630 ;
        RECT 1322.310 2589.620 1322.690 2589.630 ;
        RECT 1367.390 2589.930 1367.770 2589.940 ;
        RECT 1414.310 2589.930 1414.690 2589.940 ;
        RECT 1367.390 2589.630 1414.690 2589.930 ;
        RECT 1367.390 2589.620 1367.770 2589.630 ;
        RECT 1414.310 2589.620 1414.690 2589.630 ;
        RECT 979.150 2589.250 979.530 2589.260 ;
        RECT 958.030 2588.950 979.530 2589.250 ;
        RECT 254.905 2588.935 255.235 2588.950 ;
        RECT 351.505 2588.935 351.835 2588.950 ;
        RECT 448.105 2588.935 448.435 2588.950 ;
        RECT 544.705 2588.935 545.035 2588.950 ;
        RECT 641.305 2588.935 641.635 2588.950 ;
        RECT 737.905 2588.935 738.235 2588.950 ;
        RECT 834.505 2588.935 834.835 2588.950 ;
        RECT 979.150 2588.940 979.530 2588.950 ;
        RECT 62.625 2588.570 62.955 2588.585 ;
        RECT 110.005 2588.570 110.335 2588.585 ;
        RECT 62.625 2588.270 110.335 2588.570 ;
        RECT 62.625 2588.255 62.955 2588.270 ;
        RECT 110.005 2588.255 110.335 2588.270 ;
        RECT 31.345 2587.890 31.675 2587.905 ;
        RECT 61.705 2587.890 62.035 2587.905 ;
        RECT 31.345 2587.590 62.035 2587.890 ;
        RECT 31.345 2587.575 31.675 2587.590 ;
        RECT 61.705 2587.575 62.035 2587.590 ;
        RECT 110.925 2587.890 111.255 2587.905 ;
        RECT 138.065 2587.890 138.395 2587.905 ;
        RECT 110.925 2587.590 138.395 2587.890 ;
        RECT 110.925 2587.575 111.255 2587.590 ;
        RECT 138.065 2587.575 138.395 2587.590 ;
        RECT -4.000 2118.690 2.000 2119.140 ;
        RECT 15.705 2118.690 16.035 2118.705 ;
        RECT -4.000 2118.390 16.035 2118.690 ;
        RECT -4.000 2117.940 2.000 2118.390 ;
        RECT 15.705 2118.375 16.035 2118.390 ;
      LAYER via3 ;
        RECT 1563.380 2596.420 1563.700 2596.740 ;
        RECT 1513.700 2594.380 1514.020 2594.700 ;
        RECT 1563.380 2594.380 1563.700 2594.700 ;
        RECT 911.100 2592.340 911.420 2592.660 ;
        RECT 882.580 2589.620 882.900 2589.940 ;
        RECT 883.500 2589.620 883.820 2589.940 ;
        RECT 911.100 2589.620 911.420 2589.940 ;
        RECT 980.100 2589.620 980.420 2589.940 ;
        RECT 1051.860 2589.620 1052.180 2589.940 ;
        RECT 1096.020 2589.620 1096.340 2589.940 ;
        RECT 1172.380 2589.620 1172.700 2589.940 ;
        RECT 1218.380 2589.620 1218.700 2589.940 ;
        RECT 1221.140 2589.620 1221.460 2589.940 ;
        RECT 1270.820 2589.620 1271.140 2589.940 ;
        RECT 1322.340 2589.620 1322.660 2589.940 ;
        RECT 1367.420 2589.620 1367.740 2589.940 ;
        RECT 1414.340 2589.620 1414.660 2589.940 ;
        RECT 979.180 2588.940 979.500 2589.260 ;
      LAYER met4 ;
        RECT 1563.375 2596.415 1563.705 2596.745 ;
        RECT 1563.390 2594.705 1563.690 2596.415 ;
        RECT 1513.695 2594.375 1514.025 2594.705 ;
        RECT 1563.375 2594.375 1563.705 2594.705 ;
        RECT 911.095 2592.335 911.425 2592.665 ;
        RECT 911.110 2589.945 911.410 2592.335 ;
        RECT 882.575 2589.615 882.905 2589.945 ;
        RECT 883.495 2589.615 883.825 2589.945 ;
        RECT 911.095 2589.615 911.425 2589.945 ;
        RECT 980.095 2589.615 980.425 2589.945 ;
        RECT 1051.855 2589.690 1052.185 2589.945 ;
        RECT 1096.015 2589.690 1096.345 2589.945 ;
        RECT 1172.375 2589.690 1172.705 2589.945 ;
        RECT 1218.375 2589.690 1218.705 2589.945 ;
        RECT 882.590 2589.250 882.890 2589.615 ;
        RECT 883.510 2589.250 883.810 2589.615 ;
        RECT 882.590 2588.950 883.810 2589.250 ;
        RECT 979.175 2589.250 979.505 2589.265 ;
        RECT 980.110 2589.250 980.410 2589.615 ;
        RECT 979.175 2588.950 980.410 2589.250 ;
        RECT 979.175 2588.935 979.505 2588.950 ;
        RECT 1051.430 2588.510 1052.610 2589.690 ;
        RECT 1095.590 2588.510 1096.770 2589.690 ;
        RECT 1171.950 2588.510 1173.130 2589.690 ;
        RECT 1217.950 2588.510 1219.130 2589.690 ;
        RECT 1221.135 2589.615 1221.465 2589.945 ;
        RECT 1270.815 2589.690 1271.145 2589.945 ;
        RECT 1322.335 2589.690 1322.665 2589.945 ;
        RECT 1367.415 2589.690 1367.745 2589.945 ;
        RECT 1221.150 2589.250 1221.450 2589.615 ;
        RECT 1223.470 2589.250 1224.650 2589.690 ;
        RECT 1221.150 2588.950 1224.650 2589.250 ;
        RECT 1223.470 2588.510 1224.650 2588.950 ;
        RECT 1270.390 2588.510 1271.570 2589.690 ;
        RECT 1321.910 2588.510 1323.090 2589.690 ;
        RECT 1366.990 2588.510 1368.170 2589.690 ;
        RECT 1414.335 2589.615 1414.665 2589.945 ;
        RECT 1513.710 2589.690 1514.010 2594.375 ;
        RECT 1414.350 2589.250 1414.650 2589.615 ;
        RECT 1416.670 2589.250 1417.850 2589.690 ;
        RECT 1414.350 2588.950 1417.850 2589.250 ;
        RECT 1416.670 2588.510 1417.850 2588.950 ;
        RECT 1513.270 2588.510 1514.450 2589.690 ;
      LAYER met5 ;
        RECT 1051.220 2588.300 1096.980 2589.900 ;
        RECT 1171.740 2588.300 1219.340 2589.900 ;
        RECT 1223.260 2588.300 1271.780 2589.900 ;
        RECT 1321.700 2588.300 1368.380 2589.900 ;
        RECT 1416.460 2588.300 1514.660 2589.900 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 26.750 2597.160 27.070 2597.220 ;
        RECT 1604.550 2597.160 1604.870 2597.220 ;
        RECT 26.750 2597.020 1604.870 2597.160 ;
        RECT 26.750 2596.960 27.070 2597.020 ;
        RECT 1604.550 2596.960 1604.870 2597.020 ;
        RECT 13.870 1834.880 14.190 1834.940 ;
        RECT 26.750 1834.880 27.070 1834.940 ;
        RECT 13.870 1834.740 27.070 1834.880 ;
        RECT 13.870 1834.680 14.190 1834.740 ;
        RECT 26.750 1834.680 27.070 1834.740 ;
      LAYER via ;
        RECT 26.780 2596.960 27.040 2597.220 ;
        RECT 1604.580 2596.960 1604.840 2597.220 ;
        RECT 13.900 1834.680 14.160 1834.940 ;
        RECT 26.780 1834.680 27.040 1834.940 ;
      LAYER met2 ;
        RECT 1606.330 2597.330 1606.610 2600.000 ;
        RECT 1604.640 2597.250 1606.610 2597.330 ;
        RECT 26.780 2596.930 27.040 2597.250 ;
        RECT 1604.580 2597.190 1606.610 2597.250 ;
        RECT 1604.580 2596.930 1604.840 2597.190 ;
        RECT 26.840 1834.970 26.980 2596.930 ;
        RECT 1606.330 2596.000 1606.610 2597.190 ;
        RECT 13.900 1834.650 14.160 1834.970 ;
        RECT 26.780 1834.650 27.040 1834.970 ;
        RECT 13.960 1831.085 14.100 1834.650 ;
        RECT 13.890 1830.715 14.170 1831.085 ;
      LAYER via2 ;
        RECT 13.890 1830.760 14.170 1831.040 ;
      LAYER met3 ;
        RECT -4.000 1831.050 2.000 1831.500 ;
        RECT 13.865 1831.050 14.195 1831.065 ;
        RECT -4.000 1830.750 14.195 1831.050 ;
        RECT -4.000 1830.300 2.000 1830.750 ;
        RECT 13.865 1830.735 14.195 1830.750 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 915.930 2601.580 916.250 2601.640 ;
        RECT 2902.670 2601.580 2902.990 2601.640 ;
        RECT 915.930 2601.440 2902.990 2601.580 ;
        RECT 915.930 2601.380 916.250 2601.440 ;
        RECT 2902.670 2601.380 2902.990 2601.440 ;
      LAYER via ;
        RECT 915.960 2601.380 916.220 2601.640 ;
        RECT 2902.700 2601.380 2902.960 2601.640 ;
      LAYER met2 ;
        RECT 915.960 2601.350 916.220 2601.670 ;
        RECT 2902.700 2601.350 2902.960 2601.670 ;
        RECT 914.030 2599.370 914.310 2600.000 ;
        RECT 916.020 2599.370 916.160 2601.350 ;
        RECT 914.030 2599.230 916.160 2599.370 ;
        RECT 914.030 2596.000 914.310 2599.230 ;
        RECT 2902.760 674.405 2902.900 2601.350 ;
        RECT 2902.690 674.035 2902.970 674.405 ;
      LAYER via2 ;
        RECT 2902.690 674.080 2902.970 674.360 ;
      LAYER met3 ;
        RECT 2902.665 674.370 2902.995 674.385 ;
        RECT 2918.000 674.370 2924.000 674.820 ;
        RECT 2902.665 674.070 2924.000 674.370 ;
        RECT 2902.665 674.055 2902.995 674.070 ;
        RECT 2918.000 673.620 2924.000 674.070 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 20.310 2611.440 20.630 2611.500 ;
        RECT 1630.310 2611.440 1630.630 2611.500 ;
        RECT 20.310 2611.300 1630.630 2611.440 ;
        RECT 20.310 2611.240 20.630 2611.300 ;
        RECT 1630.310 2611.240 1630.630 2611.300 ;
      LAYER via ;
        RECT 20.340 2611.240 20.600 2611.500 ;
        RECT 1630.340 2611.240 1630.600 2611.500 ;
      LAYER met2 ;
        RECT 20.340 2611.210 20.600 2611.530 ;
        RECT 1630.340 2611.210 1630.600 2611.530 ;
        RECT 20.400 1544.125 20.540 2611.210 ;
        RECT 1630.400 2600.050 1630.540 2611.210 ;
        RECT 1630.400 2600.000 1631.850 2600.050 ;
        RECT 1630.400 2599.910 1631.910 2600.000 ;
        RECT 1631.630 2596.000 1631.910 2599.910 ;
        RECT 20.330 1543.755 20.610 1544.125 ;
      LAYER via2 ;
        RECT 20.330 1543.800 20.610 1544.080 ;
      LAYER met3 ;
        RECT -4.000 1544.090 2.000 1544.540 ;
        RECT 20.305 1544.090 20.635 1544.105 ;
        RECT -4.000 1543.790 20.635 1544.090 ;
        RECT -4.000 1543.340 2.000 1543.790 ;
        RECT 20.305 1543.775 20.635 1543.790 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 26.290 2610.080 26.610 2610.140 ;
        RECT 1656.070 2610.080 1656.390 2610.140 ;
        RECT 26.290 2609.940 1656.390 2610.080 ;
        RECT 26.290 2609.880 26.610 2609.940 ;
        RECT 1656.070 2609.880 1656.390 2609.940 ;
        RECT 13.870 1330.320 14.190 1330.380 ;
        RECT 26.290 1330.320 26.610 1330.380 ;
        RECT 13.870 1330.180 26.610 1330.320 ;
        RECT 13.870 1330.120 14.190 1330.180 ;
        RECT 26.290 1330.120 26.610 1330.180 ;
      LAYER via ;
        RECT 26.320 2609.880 26.580 2610.140 ;
        RECT 1656.100 2609.880 1656.360 2610.140 ;
        RECT 13.900 1330.120 14.160 1330.380 ;
        RECT 26.320 1330.120 26.580 1330.380 ;
      LAYER met2 ;
        RECT 26.320 2609.850 26.580 2610.170 ;
        RECT 1656.100 2609.850 1656.360 2610.170 ;
        RECT 26.380 1330.410 26.520 2609.850 ;
        RECT 1656.160 2600.050 1656.300 2609.850 ;
        RECT 1656.160 2600.000 1657.610 2600.050 ;
        RECT 1656.160 2599.910 1657.670 2600.000 ;
        RECT 1657.390 2596.000 1657.670 2599.910 ;
        RECT 13.900 1330.090 14.160 1330.410 ;
        RECT 26.320 1330.090 26.580 1330.410 ;
        RECT 13.960 1328.565 14.100 1330.090 ;
        RECT 13.890 1328.195 14.170 1328.565 ;
      LAYER via2 ;
        RECT 13.890 1328.240 14.170 1328.520 ;
      LAYER met3 ;
        RECT -4.000 1328.530 2.000 1328.980 ;
        RECT 13.865 1328.530 14.195 1328.545 ;
        RECT -4.000 1328.230 14.195 1328.530 ;
        RECT -4.000 1327.780 2.000 1328.230 ;
        RECT 13.865 1328.215 14.195 1328.230 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.930 2609.060 19.250 2609.120 ;
        RECT 1681.830 2609.060 1682.150 2609.120 ;
        RECT 18.930 2608.920 1682.150 2609.060 ;
        RECT 18.930 2608.860 19.250 2608.920 ;
        RECT 1681.830 2608.860 1682.150 2608.920 ;
      LAYER via ;
        RECT 18.960 2608.860 19.220 2609.120 ;
        RECT 1681.860 2608.860 1682.120 2609.120 ;
      LAYER met2 ;
        RECT 18.960 2608.830 19.220 2609.150 ;
        RECT 1681.860 2608.830 1682.120 2609.150 ;
        RECT 19.020 1113.005 19.160 2608.830 ;
        RECT 1681.920 2600.050 1682.060 2608.830 ;
        RECT 1681.920 2600.000 1683.370 2600.050 ;
        RECT 1681.920 2599.910 1683.430 2600.000 ;
        RECT 1683.150 2596.000 1683.430 2599.910 ;
        RECT 18.950 1112.635 19.230 1113.005 ;
      LAYER via2 ;
        RECT 18.950 1112.680 19.230 1112.960 ;
      LAYER met3 ;
        RECT -4.000 1112.970 2.000 1113.420 ;
        RECT 18.925 1112.970 19.255 1112.985 ;
        RECT -4.000 1112.670 19.255 1112.970 ;
        RECT -4.000 1112.220 2.000 1112.670 ;
        RECT 18.925 1112.655 19.255 1112.670 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1708.070 2596.650 1708.350 2596.765 ;
        RECT 1708.910 2596.650 1709.190 2600.000 ;
        RECT 1708.070 2596.510 1709.190 2596.650 ;
        RECT 1708.070 2596.395 1708.350 2596.510 ;
        RECT 1708.910 2596.000 1709.190 2596.510 ;
        RECT 18.030 2593.675 18.310 2594.045 ;
        RECT 18.100 897.445 18.240 2593.675 ;
        RECT 18.030 897.075 18.310 897.445 ;
      LAYER via2 ;
        RECT 1708.070 2596.440 1708.350 2596.720 ;
        RECT 18.030 2593.720 18.310 2594.000 ;
        RECT 18.030 897.120 18.310 897.400 ;
      LAYER met3 ;
        RECT 1708.045 2596.730 1708.375 2596.745 ;
        RECT 1707.830 2596.415 1708.375 2596.730 ;
        RECT 1207.310 2596.050 1207.690 2596.060 ;
        RECT 1232.150 2596.050 1232.530 2596.060 ;
        RECT 1207.310 2595.750 1232.530 2596.050 ;
        RECT 1207.310 2595.740 1207.690 2595.750 ;
        RECT 1232.150 2595.740 1232.530 2595.750 ;
        RECT 1316.790 2595.370 1317.170 2595.380 ;
        RECT 1316.790 2595.070 1325.410 2595.370 ;
        RECT 1316.790 2595.060 1317.170 2595.070 ;
        RECT 18.005 2594.010 18.335 2594.025 ;
        RECT 1207.310 2594.010 1207.690 2594.020 ;
        RECT 18.005 2593.710 1207.690 2594.010 ;
        RECT 18.005 2593.695 18.335 2593.710 ;
        RECT 1207.310 2593.700 1207.690 2593.710 ;
        RECT 1232.150 2594.010 1232.530 2594.020 ;
        RECT 1316.790 2594.010 1317.170 2594.020 ;
        RECT 1232.150 2593.710 1317.170 2594.010 ;
        RECT 1325.110 2594.010 1325.410 2595.070 ;
        RECT 1508.190 2594.390 1510.330 2594.690 ;
        RECT 1508.190 2594.010 1508.490 2594.390 ;
        RECT 1325.110 2593.710 1416.490 2594.010 ;
        RECT 1232.150 2593.700 1232.530 2593.710 ;
        RECT 1316.790 2593.700 1317.170 2593.710 ;
        RECT 1416.190 2593.330 1416.490 2593.710 ;
        RECT 1418.030 2593.710 1508.490 2594.010 ;
        RECT 1510.030 2594.010 1510.330 2594.390 ;
        RECT 1608.430 2594.010 1608.810 2594.020 ;
        RECT 1676.510 2594.010 1676.890 2594.020 ;
        RECT 1510.030 2593.710 1590.370 2594.010 ;
        RECT 1418.030 2593.330 1418.330 2593.710 ;
        RECT 1416.190 2593.030 1418.330 2593.330 ;
        RECT 1590.070 2593.330 1590.370 2593.710 ;
        RECT 1608.430 2593.710 1676.890 2594.010 ;
        RECT 1608.430 2593.700 1608.810 2593.710 ;
        RECT 1676.510 2593.700 1676.890 2593.710 ;
        RECT 1682.030 2594.010 1682.410 2594.020 ;
        RECT 1707.830 2594.010 1708.130 2596.415 ;
        RECT 1682.030 2593.710 1708.130 2594.010 ;
        RECT 1682.030 2593.700 1682.410 2593.710 ;
        RECT 1607.510 2593.330 1607.890 2593.340 ;
        RECT 1590.070 2593.030 1607.890 2593.330 ;
        RECT 1607.510 2593.020 1607.890 2593.030 ;
        RECT -4.000 897.410 2.000 897.860 ;
        RECT 18.005 897.410 18.335 897.425 ;
        RECT -4.000 897.110 18.335 897.410 ;
        RECT -4.000 896.660 2.000 897.110 ;
        RECT 18.005 897.095 18.335 897.110 ;
      LAYER via3 ;
        RECT 1207.340 2595.740 1207.660 2596.060 ;
        RECT 1232.180 2595.740 1232.500 2596.060 ;
        RECT 1316.820 2595.060 1317.140 2595.380 ;
        RECT 1207.340 2593.700 1207.660 2594.020 ;
        RECT 1232.180 2593.700 1232.500 2594.020 ;
        RECT 1316.820 2593.700 1317.140 2594.020 ;
        RECT 1608.460 2593.700 1608.780 2594.020 ;
        RECT 1676.540 2593.700 1676.860 2594.020 ;
        RECT 1682.060 2593.700 1682.380 2594.020 ;
        RECT 1607.540 2593.020 1607.860 2593.340 ;
      LAYER met4 ;
        RECT 1207.335 2595.735 1207.665 2596.065 ;
        RECT 1232.175 2595.735 1232.505 2596.065 ;
        RECT 1207.350 2594.025 1207.650 2595.735 ;
        RECT 1232.190 2594.025 1232.490 2595.735 ;
        RECT 1316.815 2595.055 1317.145 2595.385 ;
        RECT 1316.830 2594.025 1317.130 2595.055 ;
        RECT 1207.335 2593.695 1207.665 2594.025 ;
        RECT 1232.175 2593.695 1232.505 2594.025 ;
        RECT 1316.815 2593.695 1317.145 2594.025 ;
        RECT 1608.455 2593.695 1608.785 2594.025 ;
        RECT 1676.535 2593.695 1676.865 2594.025 ;
        RECT 1682.055 2593.695 1682.385 2594.025 ;
        RECT 1607.535 2593.015 1607.865 2593.345 ;
        RECT 1607.550 2592.650 1607.850 2593.015 ;
        RECT 1608.470 2592.650 1608.770 2593.695 ;
        RECT 1607.550 2592.350 1608.770 2592.650 ;
        RECT 1676.550 2589.690 1676.850 2593.695 ;
        RECT 1682.070 2589.690 1682.370 2593.695 ;
        RECT 1676.110 2588.510 1677.290 2589.690 ;
        RECT 1681.630 2588.510 1682.810 2589.690 ;
      LAYER met5 ;
        RECT 1675.900 2588.300 1683.020 2589.900 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 25.370 2608.720 25.690 2608.780 ;
        RECT 1732.430 2608.720 1732.750 2608.780 ;
        RECT 25.370 2608.580 1732.750 2608.720 ;
        RECT 25.370 2608.520 25.690 2608.580 ;
        RECT 1732.430 2608.520 1732.750 2608.580 ;
        RECT 13.870 682.620 14.190 682.680 ;
        RECT 25.370 682.620 25.690 682.680 ;
        RECT 13.870 682.480 25.690 682.620 ;
        RECT 13.870 682.420 14.190 682.480 ;
        RECT 25.370 682.420 25.690 682.480 ;
      LAYER via ;
        RECT 25.400 2608.520 25.660 2608.780 ;
        RECT 1732.460 2608.520 1732.720 2608.780 ;
        RECT 13.900 682.420 14.160 682.680 ;
        RECT 25.400 682.420 25.660 682.680 ;
      LAYER met2 ;
        RECT 25.400 2608.490 25.660 2608.810 ;
        RECT 1732.460 2608.490 1732.720 2608.810 ;
        RECT 25.460 682.710 25.600 2608.490 ;
        RECT 1732.520 2600.050 1732.660 2608.490 ;
        RECT 1732.520 2600.000 1734.430 2600.050 ;
        RECT 1732.520 2599.910 1734.490 2600.000 ;
        RECT 1734.210 2596.000 1734.490 2599.910 ;
        RECT 13.900 682.390 14.160 682.710 ;
        RECT 25.400 682.390 25.660 682.710 ;
        RECT 13.960 681.885 14.100 682.390 ;
        RECT 13.890 681.515 14.170 681.885 ;
      LAYER via2 ;
        RECT 13.890 681.560 14.170 681.840 ;
      LAYER met3 ;
        RECT -4.000 681.850 2.000 682.300 ;
        RECT 13.865 681.850 14.195 681.865 ;
        RECT -4.000 681.550 14.195 681.850 ;
        RECT -4.000 681.100 2.000 681.550 ;
        RECT 13.865 681.535 14.195 681.550 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1759.185 2591.225 1759.355 2596.495 ;
      LAYER mcon ;
        RECT 1759.185 2596.325 1759.355 2596.495 ;
      LAYER met1 ;
        RECT 1759.110 2596.480 1759.430 2596.540 ;
        RECT 1758.915 2596.340 1759.430 2596.480 ;
        RECT 1759.110 2596.280 1759.430 2596.340 ;
        RECT 17.550 2591.380 17.870 2591.440 ;
        RECT 1759.125 2591.380 1759.415 2591.425 ;
        RECT 17.550 2591.240 1759.415 2591.380 ;
        RECT 17.550 2591.180 17.870 2591.240 ;
        RECT 1759.125 2591.195 1759.415 2591.240 ;
      LAYER via ;
        RECT 1759.140 2596.280 1759.400 2596.540 ;
        RECT 17.580 2591.180 17.840 2591.440 ;
      LAYER met2 ;
        RECT 1759.970 2596.650 1760.250 2600.000 ;
        RECT 1759.200 2596.570 1760.250 2596.650 ;
        RECT 1759.140 2596.510 1760.250 2596.570 ;
        RECT 1759.140 2596.250 1759.400 2596.510 ;
        RECT 1759.970 2596.000 1760.250 2596.510 ;
        RECT 17.580 2591.150 17.840 2591.470 ;
        RECT 17.640 466.325 17.780 2591.150 ;
        RECT 17.570 465.955 17.850 466.325 ;
      LAYER via2 ;
        RECT 17.570 466.000 17.850 466.280 ;
      LAYER met3 ;
        RECT -4.000 466.290 2.000 466.740 ;
        RECT 17.545 466.290 17.875 466.305 ;
        RECT -4.000 465.990 17.875 466.290 ;
        RECT -4.000 465.540 2.000 465.990 ;
        RECT 17.545 465.975 17.875 465.990 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 13.870 250.820 14.190 250.880 ;
        RECT 24.450 250.820 24.770 250.880 ;
        RECT 13.870 250.680 24.770 250.820 ;
        RECT 13.870 250.620 14.190 250.680 ;
        RECT 24.450 250.620 24.770 250.680 ;
      LAYER via ;
        RECT 13.900 250.620 14.160 250.880 ;
        RECT 24.480 250.620 24.740 250.880 ;
      LAYER met2 ;
        RECT 24.470 2611.355 24.750 2611.725 ;
        RECT 1783.970 2611.355 1784.250 2611.725 ;
        RECT 24.540 250.910 24.680 2611.355 ;
        RECT 1784.040 2600.050 1784.180 2611.355 ;
        RECT 1784.040 2600.000 1785.950 2600.050 ;
        RECT 1784.040 2599.910 1786.010 2600.000 ;
        RECT 1785.730 2596.000 1786.010 2599.910 ;
        RECT 13.900 250.765 14.160 250.910 ;
        RECT 13.890 250.395 14.170 250.765 ;
        RECT 24.480 250.590 24.740 250.910 ;
      LAYER via2 ;
        RECT 24.470 2611.400 24.750 2611.680 ;
        RECT 1783.970 2611.400 1784.250 2611.680 ;
        RECT 13.890 250.440 14.170 250.720 ;
      LAYER met3 ;
        RECT 24.445 2611.690 24.775 2611.705 ;
        RECT 1783.945 2611.690 1784.275 2611.705 ;
        RECT 24.445 2611.390 1784.275 2611.690 ;
        RECT 24.445 2611.375 24.775 2611.390 ;
        RECT 1783.945 2611.375 1784.275 2611.390 ;
        RECT -4.000 250.730 2.000 251.180 ;
        RECT 13.865 250.730 14.195 250.745 ;
        RECT -4.000 250.430 14.195 250.730 ;
        RECT -4.000 249.980 2.000 250.430 ;
        RECT 13.865 250.415 14.195 250.430 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1809.730 2596.650 1810.010 2596.765 ;
        RECT 1811.490 2596.650 1811.770 2600.000 ;
        RECT 1809.730 2596.510 1811.770 2596.650 ;
        RECT 1809.730 2596.395 1810.010 2596.510 ;
        RECT 1811.490 2596.000 1811.770 2596.510 ;
        RECT 14.810 51.155 15.090 51.525 ;
        RECT 14.880 35.885 15.020 51.155 ;
        RECT 14.810 35.515 15.090 35.885 ;
      LAYER via2 ;
        RECT 1809.730 2596.440 1810.010 2596.720 ;
        RECT 14.810 51.200 15.090 51.480 ;
        RECT 14.810 35.560 15.090 35.840 ;
      LAYER met3 ;
        RECT 1808.070 2596.730 1808.450 2596.740 ;
        RECT 1809.705 2596.730 1810.035 2596.745 ;
        RECT 1808.070 2596.430 1810.035 2596.730 ;
        RECT 1808.070 2596.420 1808.450 2596.430 ;
        RECT 1809.705 2596.415 1810.035 2596.430 ;
        RECT 14.785 51.490 15.115 51.505 ;
        RECT 1808.070 51.490 1808.450 51.500 ;
        RECT 14.785 51.190 1808.450 51.490 ;
        RECT 14.785 51.175 15.115 51.190 ;
        RECT 1808.070 51.180 1808.450 51.190 ;
        RECT -4.000 35.850 2.000 36.300 ;
        RECT 14.785 35.850 15.115 35.865 ;
        RECT -4.000 35.550 15.115 35.850 ;
        RECT -4.000 35.100 2.000 35.550 ;
        RECT 14.785 35.535 15.115 35.550 ;
      LAYER via3 ;
        RECT 1808.100 2596.420 1808.420 2596.740 ;
        RECT 1808.100 51.180 1808.420 51.500 ;
      LAYER met4 ;
        RECT 1808.095 2596.415 1808.425 2596.745 ;
        RECT 1808.110 51.505 1808.410 2596.415 ;
        RECT 1808.095 51.175 1808.425 51.505 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 940.770 2601.920 941.090 2601.980 ;
        RECT 2904.510 2601.920 2904.830 2601.980 ;
        RECT 940.770 2601.780 2904.830 2601.920 ;
        RECT 940.770 2601.720 941.090 2601.780 ;
        RECT 2904.510 2601.720 2904.830 2601.780 ;
      LAYER via ;
        RECT 940.800 2601.720 941.060 2601.980 ;
        RECT 2904.540 2601.720 2904.800 2601.980 ;
      LAYER met2 ;
        RECT 940.800 2601.690 941.060 2602.010 ;
        RECT 2904.540 2601.690 2904.800 2602.010 ;
        RECT 939.330 2599.370 939.610 2600.000 ;
        RECT 940.860 2599.370 941.000 2601.690 ;
        RECT 939.330 2599.230 941.000 2599.370 ;
        RECT 939.330 2596.000 939.610 2599.230 ;
        RECT 2904.600 909.685 2904.740 2601.690 ;
        RECT 2904.530 909.315 2904.810 909.685 ;
      LAYER via2 ;
        RECT 2904.530 909.360 2904.810 909.640 ;
      LAYER met3 ;
        RECT 2904.505 909.650 2904.835 909.665 ;
        RECT 2918.000 909.650 2924.000 910.100 ;
        RECT 2904.505 909.350 2924.000 909.650 ;
        RECT 2904.505 909.335 2904.835 909.350 ;
        RECT 2918.000 908.900 2924.000 909.350 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2898.530 2551.260 2898.850 2551.320 ;
        RECT 2899.910 2551.260 2900.230 2551.320 ;
        RECT 2898.530 2551.120 2900.230 2551.260 ;
        RECT 2898.530 2551.060 2898.850 2551.120 ;
        RECT 2899.910 2551.060 2900.230 2551.120 ;
      LAYER via ;
        RECT 2898.560 2551.060 2898.820 2551.320 ;
        RECT 2899.940 2551.060 2900.200 2551.320 ;
      LAYER met2 ;
        RECT 965.090 2596.650 965.370 2600.000 ;
        RECT 965.630 2596.650 965.910 2596.765 ;
        RECT 965.090 2596.510 965.910 2596.650 ;
        RECT 965.090 2596.000 965.370 2596.510 ;
        RECT 965.630 2596.395 965.910 2596.510 ;
        RECT 1860.330 2594.355 1860.610 2594.725 ;
        RECT 1860.400 2590.645 1860.540 2594.355 ;
        RECT 1860.330 2590.275 1860.610 2590.645 ;
        RECT 2898.550 2590.275 2898.830 2590.645 ;
        RECT 2898.620 2551.350 2898.760 2590.275 ;
        RECT 2898.560 2551.030 2898.820 2551.350 ;
        RECT 2899.940 2551.030 2900.200 2551.350 ;
        RECT 2900.000 1144.285 2900.140 2551.030 ;
        RECT 2899.930 1143.915 2900.210 1144.285 ;
      LAYER via2 ;
        RECT 965.630 2596.440 965.910 2596.720 ;
        RECT 1860.330 2594.400 1860.610 2594.680 ;
        RECT 1860.330 2590.320 1860.610 2590.600 ;
        RECT 2898.550 2590.320 2898.830 2590.600 ;
        RECT 2899.930 1143.960 2900.210 1144.240 ;
      LAYER met3 ;
        RECT 965.605 2596.740 965.935 2596.745 ;
        RECT 965.350 2596.730 965.935 2596.740 ;
        RECT 965.150 2596.430 965.935 2596.730 ;
        RECT 965.350 2596.420 965.935 2596.430 ;
        RECT 965.605 2596.415 965.935 2596.420 ;
        RECT 1836.590 2594.690 1836.970 2594.700 ;
        RECT 1860.305 2594.690 1860.635 2594.705 ;
        RECT 1836.590 2594.390 1860.635 2594.690 ;
        RECT 1836.590 2594.380 1836.970 2594.390 ;
        RECT 1860.305 2594.375 1860.635 2594.390 ;
        RECT 1173.270 2591.970 1173.650 2591.980 ;
        RECT 1181.550 2591.970 1181.930 2591.980 ;
        RECT 1173.270 2591.670 1181.930 2591.970 ;
        RECT 1173.270 2591.660 1173.650 2591.670 ;
        RECT 1181.550 2591.660 1181.930 2591.670 ;
        RECT 1495.270 2591.290 1495.650 2591.300 ;
        RECT 1475.990 2590.990 1495.650 2591.290 ;
        RECT 965.350 2590.610 965.730 2590.620 ;
        RECT 1173.270 2590.610 1173.650 2590.620 ;
        RECT 965.350 2590.310 1173.650 2590.610 ;
        RECT 965.350 2590.300 965.730 2590.310 ;
        RECT 1173.270 2590.300 1173.650 2590.310 ;
        RECT 1181.550 2590.610 1181.930 2590.620 ;
        RECT 1475.990 2590.610 1476.290 2590.990 ;
        RECT 1495.270 2590.980 1495.650 2590.990 ;
        RECT 1181.550 2590.310 1476.290 2590.610 ;
        RECT 1496.190 2590.610 1496.570 2590.620 ;
        RECT 1835.670 2590.610 1836.050 2590.620 ;
        RECT 1496.190 2590.310 1836.050 2590.610 ;
        RECT 1181.550 2590.300 1181.930 2590.310 ;
        RECT 1496.190 2590.300 1496.570 2590.310 ;
        RECT 1835.670 2590.300 1836.050 2590.310 ;
        RECT 1860.305 2590.610 1860.635 2590.625 ;
        RECT 2898.525 2590.610 2898.855 2590.625 ;
        RECT 1860.305 2590.310 2898.855 2590.610 ;
        RECT 1860.305 2590.295 1860.635 2590.310 ;
        RECT 2898.525 2590.295 2898.855 2590.310 ;
        RECT 2899.905 1144.250 2900.235 1144.265 ;
        RECT 2918.000 1144.250 2924.000 1144.700 ;
        RECT 2899.905 1143.950 2924.000 1144.250 ;
        RECT 2899.905 1143.935 2900.235 1143.950 ;
        RECT 2918.000 1143.500 2924.000 1143.950 ;
      LAYER via3 ;
        RECT 965.380 2596.420 965.700 2596.740 ;
        RECT 1836.620 2594.380 1836.940 2594.700 ;
        RECT 1173.300 2591.660 1173.620 2591.980 ;
        RECT 1181.580 2591.660 1181.900 2591.980 ;
        RECT 965.380 2590.300 965.700 2590.620 ;
        RECT 1173.300 2590.300 1173.620 2590.620 ;
        RECT 1181.580 2590.300 1181.900 2590.620 ;
        RECT 1495.300 2590.980 1495.620 2591.300 ;
        RECT 1496.220 2590.300 1496.540 2590.620 ;
        RECT 1835.700 2590.300 1836.020 2590.620 ;
      LAYER met4 ;
        RECT 965.375 2596.415 965.705 2596.745 ;
        RECT 965.390 2590.625 965.690 2596.415 ;
        RECT 1836.615 2594.375 1836.945 2594.705 ;
        RECT 1836.630 2592.650 1836.930 2594.375 ;
        RECT 1835.710 2592.350 1836.930 2592.650 ;
        RECT 1173.295 2591.655 1173.625 2591.985 ;
        RECT 1181.575 2591.655 1181.905 2591.985 ;
        RECT 1173.310 2590.625 1173.610 2591.655 ;
        RECT 1181.590 2590.625 1181.890 2591.655 ;
        RECT 1495.295 2590.975 1495.625 2591.305 ;
        RECT 965.375 2590.295 965.705 2590.625 ;
        RECT 1173.295 2590.295 1173.625 2590.625 ;
        RECT 1181.575 2590.295 1181.905 2590.625 ;
        RECT 1495.310 2589.250 1495.610 2590.975 ;
        RECT 1835.710 2590.625 1836.010 2592.350 ;
        RECT 1496.215 2590.295 1496.545 2590.625 ;
        RECT 1835.695 2590.295 1836.025 2590.625 ;
        RECT 1496.230 2589.250 1496.530 2590.295 ;
        RECT 1495.310 2588.950 1496.530 2589.250 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 990.850 2596.650 991.130 2600.000 ;
        RECT 991.850 2596.650 992.130 2596.765 ;
        RECT 990.850 2596.510 992.130 2596.650 ;
        RECT 990.850 2596.000 991.130 2596.510 ;
        RECT 991.850 2596.395 992.130 2596.510 ;
        RECT 1859.410 2591.635 1859.690 2592.005 ;
        RECT 2898.090 2591.635 2898.370 2592.005 ;
        RECT 1859.480 2590.645 1859.620 2591.635 ;
        RECT 1859.410 2590.275 1859.690 2590.645 ;
        RECT 2898.160 1378.885 2898.300 2591.635 ;
        RECT 2898.090 1378.515 2898.370 1378.885 ;
      LAYER via2 ;
        RECT 991.850 2596.440 992.130 2596.720 ;
        RECT 1859.410 2591.680 1859.690 2591.960 ;
        RECT 2898.090 2591.680 2898.370 2591.960 ;
        RECT 1859.410 2590.320 1859.690 2590.600 ;
        RECT 2898.090 1378.560 2898.370 1378.840 ;
      LAYER met3 ;
        RECT 991.825 2596.740 992.155 2596.745 ;
        RECT 991.825 2596.730 992.410 2596.740 ;
        RECT 1171.430 2596.730 1171.810 2596.740 ;
        RECT 1182.470 2596.730 1182.850 2596.740 ;
        RECT 991.825 2596.430 992.610 2596.730 ;
        RECT 1171.430 2596.430 1182.850 2596.730 ;
        RECT 991.825 2596.420 992.410 2596.430 ;
        RECT 1171.430 2596.420 1171.810 2596.430 ;
        RECT 1182.470 2596.420 1182.850 2596.430 ;
        RECT 991.825 2596.415 992.155 2596.420 ;
        RECT 992.030 2591.970 992.410 2591.980 ;
        RECT 1171.430 2591.970 1171.810 2591.980 ;
        RECT 992.030 2591.670 1171.810 2591.970 ;
        RECT 992.030 2591.660 992.410 2591.670 ;
        RECT 1171.430 2591.660 1171.810 2591.670 ;
        RECT 1182.470 2591.970 1182.850 2591.980 ;
        RECT 1836.590 2591.970 1836.970 2591.980 ;
        RECT 1182.470 2591.670 1836.970 2591.970 ;
        RECT 1182.470 2591.660 1182.850 2591.670 ;
        RECT 1836.590 2591.660 1836.970 2591.670 ;
        RECT 1859.385 2591.970 1859.715 2591.985 ;
        RECT 2898.065 2591.970 2898.395 2591.985 ;
        RECT 1859.385 2591.670 2898.395 2591.970 ;
        RECT 1859.385 2591.655 1859.715 2591.670 ;
        RECT 2898.065 2591.655 2898.395 2591.670 ;
        RECT 1836.590 2590.610 1836.970 2590.620 ;
        RECT 1859.385 2590.610 1859.715 2590.625 ;
        RECT 1836.590 2590.310 1859.715 2590.610 ;
        RECT 1836.590 2590.300 1836.970 2590.310 ;
        RECT 1859.385 2590.295 1859.715 2590.310 ;
        RECT 2898.065 1378.850 2898.395 1378.865 ;
        RECT 2918.000 1378.850 2924.000 1379.300 ;
        RECT 2898.065 1378.550 2924.000 1378.850 ;
        RECT 2898.065 1378.535 2898.395 1378.550 ;
        RECT 2918.000 1378.100 2924.000 1378.550 ;
      LAYER via3 ;
        RECT 992.060 2596.420 992.380 2596.740 ;
        RECT 1171.460 2596.420 1171.780 2596.740 ;
        RECT 1182.500 2596.420 1182.820 2596.740 ;
        RECT 992.060 2591.660 992.380 2591.980 ;
        RECT 1171.460 2591.660 1171.780 2591.980 ;
        RECT 1182.500 2591.660 1182.820 2591.980 ;
        RECT 1836.620 2591.660 1836.940 2591.980 ;
        RECT 1836.620 2590.300 1836.940 2590.620 ;
      LAYER met4 ;
        RECT 992.055 2596.415 992.385 2596.745 ;
        RECT 1171.455 2596.415 1171.785 2596.745 ;
        RECT 1182.495 2596.415 1182.825 2596.745 ;
        RECT 992.070 2591.985 992.370 2596.415 ;
        RECT 1171.470 2591.985 1171.770 2596.415 ;
        RECT 1182.510 2591.985 1182.810 2596.415 ;
        RECT 992.055 2591.655 992.385 2591.985 ;
        RECT 1171.455 2591.655 1171.785 2591.985 ;
        RECT 1182.495 2591.655 1182.825 2591.985 ;
        RECT 1836.615 2591.655 1836.945 2591.985 ;
        RECT 1836.630 2590.625 1836.930 2591.655 ;
        RECT 1836.615 2590.295 1836.945 2590.625 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1018.050 2602.260 1018.370 2602.320 ;
        RECT 1847.430 2602.260 1847.750 2602.320 ;
        RECT 1018.050 2602.120 1847.750 2602.260 ;
        RECT 1018.050 2602.060 1018.370 2602.120 ;
        RECT 1847.430 2602.060 1847.750 2602.120 ;
        RECT 1848.350 1614.560 1848.670 1614.620 ;
        RECT 2900.370 1614.560 2900.690 1614.620 ;
        RECT 1848.350 1614.420 2900.690 1614.560 ;
        RECT 1848.350 1614.360 1848.670 1614.420 ;
        RECT 2900.370 1614.360 2900.690 1614.420 ;
      LAYER via ;
        RECT 1018.080 2602.060 1018.340 2602.320 ;
        RECT 1847.460 2602.060 1847.720 2602.320 ;
        RECT 1848.380 1614.360 1848.640 1614.620 ;
        RECT 2900.400 1614.360 2900.660 1614.620 ;
      LAYER met2 ;
        RECT 1018.080 2602.030 1018.340 2602.350 ;
        RECT 1847.460 2602.030 1847.720 2602.350 ;
        RECT 1016.610 2599.370 1016.890 2600.000 ;
        RECT 1018.140 2599.370 1018.280 2602.030 ;
        RECT 1016.610 2599.230 1018.280 2599.370 ;
        RECT 1016.610 2596.000 1016.890 2599.230 ;
        RECT 1847.520 1614.050 1847.660 2602.030 ;
        RECT 1848.380 1614.330 1848.640 1614.650 ;
        RECT 2900.400 1614.330 2900.660 1614.650 ;
        RECT 1848.440 1614.050 1848.580 1614.330 ;
        RECT 1847.520 1613.910 1848.580 1614.050 ;
        RECT 2900.460 1613.485 2900.600 1614.330 ;
        RECT 2900.390 1613.115 2900.670 1613.485 ;
      LAYER via2 ;
        RECT 2900.390 1613.160 2900.670 1613.440 ;
      LAYER met3 ;
        RECT 2900.365 1613.450 2900.695 1613.465 ;
        RECT 2918.000 1613.450 2924.000 1613.900 ;
        RECT 2900.365 1613.150 2924.000 1613.450 ;
        RECT 2900.365 1613.135 2900.695 1613.150 ;
        RECT 2918.000 1612.700 2924.000 1613.150 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1043.810 2602.940 1044.130 2603.000 ;
        RECT 1848.350 2602.940 1848.670 2603.000 ;
        RECT 1043.810 2602.800 1848.670 2602.940 ;
        RECT 1043.810 2602.740 1044.130 2602.800 ;
        RECT 1848.350 2602.740 1848.670 2602.800 ;
        RECT 1848.350 1849.160 1848.670 1849.220 ;
        RECT 2899.450 1849.160 2899.770 1849.220 ;
        RECT 1848.350 1849.020 2899.770 1849.160 ;
        RECT 1848.350 1848.960 1848.670 1849.020 ;
        RECT 2899.450 1848.960 2899.770 1849.020 ;
      LAYER via ;
        RECT 1043.840 2602.740 1044.100 2603.000 ;
        RECT 1848.380 2602.740 1848.640 2603.000 ;
        RECT 1848.380 1848.960 1848.640 1849.220 ;
        RECT 2899.480 1848.960 2899.740 1849.220 ;
      LAYER met2 ;
        RECT 1043.840 2602.710 1044.100 2603.030 ;
        RECT 1848.380 2602.710 1848.640 2603.030 ;
        RECT 1041.910 2599.370 1042.190 2600.000 ;
        RECT 1043.900 2599.370 1044.040 2602.710 ;
        RECT 1041.910 2599.230 1044.040 2599.370 ;
        RECT 1041.910 2596.000 1042.190 2599.230 ;
        RECT 1848.440 1849.250 1848.580 2602.710 ;
        RECT 1848.380 1848.930 1848.640 1849.250 ;
        RECT 2899.480 1848.930 2899.740 1849.250 ;
        RECT 2899.540 1848.085 2899.680 1848.930 ;
        RECT 2899.470 1847.715 2899.750 1848.085 ;
      LAYER via2 ;
        RECT 2899.470 1847.760 2899.750 1848.040 ;
      LAYER met3 ;
        RECT 2899.445 1848.050 2899.775 1848.065 ;
        RECT 2918.000 1848.050 2924.000 1848.500 ;
        RECT 2899.445 1847.750 2924.000 1848.050 ;
        RECT 2899.445 1847.735 2899.775 1847.750 ;
        RECT 2918.000 1847.300 2924.000 1847.750 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1069.110 2614.500 1069.430 2614.560 ;
        RECT 1853.870 2614.500 1854.190 2614.560 ;
        RECT 1069.110 2614.360 1854.190 2614.500 ;
        RECT 1069.110 2614.300 1069.430 2614.360 ;
        RECT 1853.870 2614.300 1854.190 2614.360 ;
        RECT 1853.870 2083.760 1854.190 2083.820 ;
        RECT 2899.450 2083.760 2899.770 2083.820 ;
        RECT 1853.870 2083.620 2899.770 2083.760 ;
        RECT 1853.870 2083.560 1854.190 2083.620 ;
        RECT 2899.450 2083.560 2899.770 2083.620 ;
      LAYER via ;
        RECT 1069.140 2614.300 1069.400 2614.560 ;
        RECT 1853.900 2614.300 1854.160 2614.560 ;
        RECT 1853.900 2083.560 1854.160 2083.820 ;
        RECT 2899.480 2083.560 2899.740 2083.820 ;
      LAYER met2 ;
        RECT 1069.140 2614.270 1069.400 2614.590 ;
        RECT 1853.900 2614.270 1854.160 2614.590 ;
        RECT 1067.670 2599.370 1067.950 2600.000 ;
        RECT 1069.200 2599.370 1069.340 2614.270 ;
        RECT 1067.670 2599.230 1069.340 2599.370 ;
        RECT 1067.670 2596.000 1067.950 2599.230 ;
        RECT 1853.960 2083.850 1854.100 2614.270 ;
        RECT 1853.900 2083.530 1854.160 2083.850 ;
        RECT 2899.480 2083.530 2899.740 2083.850 ;
        RECT 2899.540 2082.685 2899.680 2083.530 ;
        RECT 2899.470 2082.315 2899.750 2082.685 ;
      LAYER via2 ;
        RECT 2899.470 2082.360 2899.750 2082.640 ;
      LAYER met3 ;
        RECT 2899.445 2082.650 2899.775 2082.665 ;
        RECT 2918.000 2082.650 2924.000 2083.100 ;
        RECT 2899.445 2082.350 2924.000 2082.650 ;
        RECT 2899.445 2082.335 2899.775 2082.350 ;
        RECT 2918.000 2081.900 2924.000 2082.350 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1095.330 2614.840 1095.650 2614.900 ;
        RECT 1855.250 2614.840 1855.570 2614.900 ;
        RECT 1095.330 2614.700 1855.570 2614.840 ;
        RECT 1095.330 2614.640 1095.650 2614.700 ;
        RECT 1855.250 2614.640 1855.570 2614.700 ;
        RECT 1855.250 2318.360 1855.570 2318.420 ;
        RECT 2899.450 2318.360 2899.770 2318.420 ;
        RECT 1855.250 2318.220 2899.770 2318.360 ;
        RECT 1855.250 2318.160 1855.570 2318.220 ;
        RECT 2899.450 2318.160 2899.770 2318.220 ;
      LAYER via ;
        RECT 1095.360 2614.640 1095.620 2614.900 ;
        RECT 1855.280 2614.640 1855.540 2614.900 ;
        RECT 1855.280 2318.160 1855.540 2318.420 ;
        RECT 2899.480 2318.160 2899.740 2318.420 ;
      LAYER met2 ;
        RECT 1095.360 2614.610 1095.620 2614.930 ;
        RECT 1855.280 2614.610 1855.540 2614.930 ;
        RECT 1093.430 2599.370 1093.710 2600.000 ;
        RECT 1095.420 2599.370 1095.560 2614.610 ;
        RECT 1093.430 2599.230 1095.560 2599.370 ;
        RECT 1093.430 2596.000 1093.710 2599.230 ;
        RECT 1855.340 2318.450 1855.480 2614.610 ;
        RECT 1855.280 2318.130 1855.540 2318.450 ;
        RECT 2899.480 2318.130 2899.740 2318.450 ;
        RECT 2899.540 2317.285 2899.680 2318.130 ;
        RECT 2899.470 2316.915 2899.750 2317.285 ;
      LAYER via2 ;
        RECT 2899.470 2316.960 2899.750 2317.240 ;
      LAYER met3 ;
        RECT 2899.445 2317.250 2899.775 2317.265 ;
        RECT 2918.000 2317.250 2924.000 2317.700 ;
        RECT 2899.445 2316.950 2924.000 2317.250 ;
        RECT 2899.445 2316.935 2899.775 2316.950 ;
        RECT 2918.000 2316.500 2924.000 2316.950 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1852.490 151.540 1852.810 151.600 ;
        RECT 2901.290 151.540 2901.610 151.600 ;
        RECT 1852.490 151.400 2901.610 151.540 ;
        RECT 1852.490 151.340 1852.810 151.400 ;
        RECT 2901.290 151.340 2901.610 151.400 ;
      LAYER via ;
        RECT 1852.520 151.340 1852.780 151.600 ;
        RECT 2901.320 151.340 2901.580 151.600 ;
      LAYER met2 ;
        RECT 872.710 2612.715 872.990 2613.085 ;
        RECT 1852.510 2612.715 1852.790 2613.085 ;
        RECT 871.250 2599.370 871.530 2600.000 ;
        RECT 872.780 2599.370 872.920 2612.715 ;
        RECT 871.250 2599.230 872.920 2599.370 ;
        RECT 871.250 2596.000 871.530 2599.230 ;
        RECT 1852.580 151.630 1852.720 2612.715 ;
        RECT 1852.520 151.310 1852.780 151.630 ;
        RECT 2901.320 151.310 2901.580 151.630 ;
        RECT 2901.380 146.725 2901.520 151.310 ;
        RECT 2901.310 146.355 2901.590 146.725 ;
      LAYER via2 ;
        RECT 872.710 2612.760 872.990 2613.040 ;
        RECT 1852.510 2612.760 1852.790 2613.040 ;
        RECT 2901.310 146.400 2901.590 146.680 ;
      LAYER met3 ;
        RECT 872.685 2613.050 873.015 2613.065 ;
        RECT 1852.485 2613.050 1852.815 2613.065 ;
        RECT 872.685 2612.750 1852.815 2613.050 ;
        RECT 872.685 2612.735 873.015 2612.750 ;
        RECT 1852.485 2612.735 1852.815 2612.750 ;
        RECT 2901.285 146.690 2901.615 146.705 ;
        RECT 2918.000 146.690 2924.000 147.140 ;
        RECT 2901.285 146.390 2924.000 146.690 ;
        RECT 2901.285 146.375 2901.615 146.390 ;
        RECT 2918.000 145.940 2924.000 146.390 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1855.710 2497.540 1856.030 2497.600 ;
        RECT 2899.450 2497.540 2899.770 2497.600 ;
        RECT 1855.710 2497.400 2899.770 2497.540 ;
        RECT 1855.710 2497.340 1856.030 2497.400 ;
        RECT 2899.450 2497.340 2899.770 2497.400 ;
      LAYER via ;
        RECT 1855.740 2497.340 1856.000 2497.600 ;
        RECT 2899.480 2497.340 2899.740 2497.600 ;
      LAYER met2 ;
        RECT 1127.470 2596.650 1127.750 2600.000 ;
        RECT 1128.930 2596.650 1129.210 2596.765 ;
        RECT 1127.470 2596.510 1129.210 2596.650 ;
        RECT 1127.470 2596.000 1127.750 2596.510 ;
        RECT 1128.930 2596.395 1129.210 2596.510 ;
        RECT 1855.730 2589.595 1856.010 2589.965 ;
        RECT 1855.800 2497.630 1855.940 2589.595 ;
        RECT 1855.740 2497.310 1856.000 2497.630 ;
        RECT 2899.480 2497.310 2899.740 2497.630 ;
        RECT 2899.540 2493.405 2899.680 2497.310 ;
        RECT 2899.470 2493.035 2899.750 2493.405 ;
      LAYER via2 ;
        RECT 1128.930 2596.440 1129.210 2596.720 ;
        RECT 1855.730 2589.640 1856.010 2589.920 ;
        RECT 2899.470 2493.080 2899.750 2493.360 ;
      LAYER met3 ;
        RECT 1128.905 2596.730 1129.235 2596.745 ;
        RECT 1400.510 2596.730 1400.890 2596.740 ;
        RECT 1424.430 2596.730 1424.810 2596.740 ;
        RECT 1128.905 2596.415 1129.450 2596.730 ;
        RECT 1400.510 2596.430 1424.810 2596.730 ;
        RECT 1400.510 2596.420 1400.890 2596.430 ;
        RECT 1424.430 2596.420 1424.810 2596.430 ;
        RECT 1129.150 2595.370 1129.450 2596.415 ;
        RECT 1184.310 2595.370 1184.690 2595.380 ;
        RECT 1129.150 2595.070 1184.690 2595.370 ;
        RECT 1184.310 2595.060 1184.690 2595.070 ;
        RECT 1364.630 2595.370 1365.010 2595.380 ;
        RECT 1400.510 2595.370 1400.890 2595.380 ;
        RECT 1364.630 2595.070 1400.890 2595.370 ;
        RECT 1364.630 2595.060 1365.010 2595.070 ;
        RECT 1400.510 2595.060 1400.890 2595.070 ;
        RECT 1268.030 2594.690 1268.410 2594.700 ;
        RECT 1471.350 2594.690 1471.730 2594.700 ;
        RECT 1494.350 2594.690 1494.730 2594.700 ;
        RECT 1217.470 2594.390 1222.370 2594.690 ;
        RECT 1184.310 2593.330 1184.690 2593.340 ;
        RECT 1217.470 2593.330 1217.770 2594.390 ;
        RECT 1184.310 2593.030 1217.770 2593.330 ;
        RECT 1222.070 2593.330 1222.370 2594.390 ;
        RECT 1268.030 2594.390 1324.490 2594.690 ;
        RECT 1268.030 2594.380 1268.410 2594.390 ;
        RECT 1268.030 2593.330 1268.410 2593.340 ;
        RECT 1222.070 2593.030 1268.410 2593.330 ;
        RECT 1324.190 2593.330 1324.490 2594.390 ;
        RECT 1471.350 2594.390 1494.730 2594.690 ;
        RECT 1471.350 2594.380 1471.730 2594.390 ;
        RECT 1494.350 2594.380 1494.730 2594.390 ;
        RECT 1364.630 2593.330 1365.010 2593.340 ;
        RECT 1324.190 2593.030 1365.010 2593.330 ;
        RECT 1184.310 2593.020 1184.690 2593.030 ;
        RECT 1268.030 2593.020 1268.410 2593.030 ;
        RECT 1364.630 2593.020 1365.010 2593.030 ;
        RECT 1424.430 2593.330 1424.810 2593.340 ;
        RECT 1471.350 2593.330 1471.730 2593.340 ;
        RECT 1424.430 2593.030 1471.730 2593.330 ;
        RECT 1424.430 2593.020 1424.810 2593.030 ;
        RECT 1471.350 2593.020 1471.730 2593.030 ;
        RECT 1494.350 2593.330 1494.730 2593.340 ;
        RECT 1509.070 2593.330 1509.450 2593.340 ;
        RECT 1494.350 2593.030 1509.450 2593.330 ;
        RECT 1494.350 2593.020 1494.730 2593.030 ;
        RECT 1509.070 2593.020 1509.450 2593.030 ;
        RECT 1510.910 2589.930 1511.290 2589.940 ;
        RECT 1855.705 2589.930 1856.035 2589.945 ;
        RECT 1510.910 2589.630 1856.035 2589.930 ;
        RECT 1510.910 2589.620 1511.290 2589.630 ;
        RECT 1855.705 2589.615 1856.035 2589.630 ;
        RECT 2899.445 2493.370 2899.775 2493.385 ;
        RECT 2918.000 2493.370 2924.000 2493.820 ;
        RECT 2899.445 2493.070 2924.000 2493.370 ;
        RECT 2899.445 2493.055 2899.775 2493.070 ;
        RECT 2918.000 2492.620 2924.000 2493.070 ;
      LAYER via3 ;
        RECT 1400.540 2596.420 1400.860 2596.740 ;
        RECT 1424.460 2596.420 1424.780 2596.740 ;
        RECT 1184.340 2595.060 1184.660 2595.380 ;
        RECT 1364.660 2595.060 1364.980 2595.380 ;
        RECT 1400.540 2595.060 1400.860 2595.380 ;
        RECT 1184.340 2593.020 1184.660 2593.340 ;
        RECT 1268.060 2594.380 1268.380 2594.700 ;
        RECT 1268.060 2593.020 1268.380 2593.340 ;
        RECT 1471.380 2594.380 1471.700 2594.700 ;
        RECT 1494.380 2594.380 1494.700 2594.700 ;
        RECT 1364.660 2593.020 1364.980 2593.340 ;
        RECT 1424.460 2593.020 1424.780 2593.340 ;
        RECT 1471.380 2593.020 1471.700 2593.340 ;
        RECT 1494.380 2593.020 1494.700 2593.340 ;
        RECT 1509.100 2593.020 1509.420 2593.340 ;
        RECT 1510.940 2589.620 1511.260 2589.940 ;
      LAYER met4 ;
        RECT 1400.535 2596.415 1400.865 2596.745 ;
        RECT 1424.455 2596.415 1424.785 2596.745 ;
        RECT 1400.550 2595.385 1400.850 2596.415 ;
        RECT 1184.335 2595.055 1184.665 2595.385 ;
        RECT 1364.655 2595.055 1364.985 2595.385 ;
        RECT 1400.535 2595.055 1400.865 2595.385 ;
        RECT 1184.350 2593.345 1184.650 2595.055 ;
        RECT 1268.055 2594.375 1268.385 2594.705 ;
        RECT 1268.070 2593.345 1268.370 2594.375 ;
        RECT 1364.670 2593.345 1364.970 2595.055 ;
        RECT 1424.470 2593.345 1424.770 2596.415 ;
        RECT 1471.375 2594.375 1471.705 2594.705 ;
        RECT 1494.375 2594.375 1494.705 2594.705 ;
        RECT 1471.390 2593.345 1471.690 2594.375 ;
        RECT 1494.390 2593.345 1494.690 2594.375 ;
        RECT 1184.335 2593.015 1184.665 2593.345 ;
        RECT 1268.055 2593.015 1268.385 2593.345 ;
        RECT 1364.655 2593.015 1364.985 2593.345 ;
        RECT 1424.455 2593.015 1424.785 2593.345 ;
        RECT 1471.375 2593.015 1471.705 2593.345 ;
        RECT 1494.375 2593.015 1494.705 2593.345 ;
        RECT 1509.095 2593.015 1509.425 2593.345 ;
        RECT 1509.110 2589.250 1509.410 2593.015 ;
        RECT 1510.935 2589.615 1511.265 2589.945 ;
        RECT 1510.950 2589.250 1511.250 2589.615 ;
        RECT 1509.110 2588.950 1511.250 2589.250 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1158.810 2725.680 1159.130 2725.740 ;
        RECT 2900.370 2725.680 2900.690 2725.740 ;
        RECT 1158.810 2725.540 2900.690 2725.680 ;
        RECT 1158.810 2725.480 1159.130 2725.540 ;
        RECT 2900.370 2725.480 2900.690 2725.540 ;
        RECT 1152.370 2632.520 1152.690 2632.580 ;
        RECT 1158.810 2632.520 1159.130 2632.580 ;
        RECT 1152.370 2632.380 1159.130 2632.520 ;
        RECT 1152.370 2632.320 1152.690 2632.380 ;
        RECT 1158.810 2632.320 1159.130 2632.380 ;
      LAYER via ;
        RECT 1158.840 2725.480 1159.100 2725.740 ;
        RECT 2900.400 2725.480 2900.660 2725.740 ;
        RECT 1152.400 2632.320 1152.660 2632.580 ;
        RECT 1158.840 2632.320 1159.100 2632.580 ;
      LAYER met2 ;
        RECT 2900.390 2727.635 2900.670 2728.005 ;
        RECT 2900.460 2725.770 2900.600 2727.635 ;
        RECT 1158.840 2725.450 1159.100 2725.770 ;
        RECT 2900.400 2725.450 2900.660 2725.770 ;
        RECT 1158.900 2632.610 1159.040 2725.450 ;
        RECT 1152.400 2632.290 1152.660 2632.610 ;
        RECT 1158.840 2632.290 1159.100 2632.610 ;
        RECT 1152.460 2600.050 1152.600 2632.290 ;
        RECT 1152.460 2600.000 1153.450 2600.050 ;
        RECT 1152.460 2599.910 1153.510 2600.000 ;
        RECT 1153.230 2596.000 1153.510 2599.910 ;
      LAYER via2 ;
        RECT 2900.390 2727.680 2900.670 2727.960 ;
      LAYER met3 ;
        RECT 2900.365 2727.970 2900.695 2727.985 ;
        RECT 2918.000 2727.970 2924.000 2728.420 ;
        RECT 2900.365 2727.670 2924.000 2727.970 ;
        RECT 2900.365 2727.655 2900.695 2727.670 ;
        RECT 2918.000 2727.220 2924.000 2727.670 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1179.510 2960.280 1179.830 2960.340 ;
        RECT 2900.370 2960.280 2900.690 2960.340 ;
        RECT 1179.510 2960.140 2900.690 2960.280 ;
        RECT 1179.510 2960.080 1179.830 2960.140 ;
        RECT 2900.370 2960.080 2900.690 2960.140 ;
        RECT 1173.070 2632.520 1173.390 2632.580 ;
        RECT 1179.510 2632.520 1179.830 2632.580 ;
        RECT 1173.070 2632.380 1179.830 2632.520 ;
        RECT 1173.070 2632.320 1173.390 2632.380 ;
        RECT 1179.510 2632.320 1179.830 2632.380 ;
      LAYER via ;
        RECT 1179.540 2960.080 1179.800 2960.340 ;
        RECT 2900.400 2960.080 2900.660 2960.340 ;
        RECT 1173.100 2632.320 1173.360 2632.580 ;
        RECT 1179.540 2632.320 1179.800 2632.580 ;
      LAYER met2 ;
        RECT 2900.390 2962.235 2900.670 2962.605 ;
        RECT 2900.460 2960.370 2900.600 2962.235 ;
        RECT 1179.540 2960.050 1179.800 2960.370 ;
        RECT 2900.400 2960.050 2900.660 2960.370 ;
        RECT 1179.600 2632.610 1179.740 2960.050 ;
        RECT 1173.100 2632.290 1173.360 2632.610 ;
        RECT 1179.540 2632.290 1179.800 2632.610 ;
        RECT 1173.160 2601.410 1173.300 2632.290 ;
        RECT 1173.160 2601.270 1177.440 2601.410 ;
        RECT 1177.300 2600.050 1177.440 2601.270 ;
        RECT 1177.300 2600.000 1179.210 2600.050 ;
        RECT 1177.300 2599.910 1179.270 2600.000 ;
        RECT 1178.990 2596.000 1179.270 2599.910 ;
      LAYER via2 ;
        RECT 2900.390 2962.280 2900.670 2962.560 ;
      LAYER met3 ;
        RECT 2900.365 2962.570 2900.695 2962.585 ;
        RECT 2918.000 2962.570 2924.000 2963.020 ;
        RECT 2900.365 2962.270 2924.000 2962.570 ;
        RECT 2900.365 2962.255 2900.695 2962.270 ;
        RECT 2918.000 2961.820 2924.000 2962.270 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1207.110 3194.880 1207.430 3194.940 ;
        RECT 2900.370 3194.880 2900.690 3194.940 ;
        RECT 1207.110 3194.740 2900.690 3194.880 ;
        RECT 1207.110 3194.680 1207.430 3194.740 ;
        RECT 2900.370 3194.680 2900.690 3194.740 ;
      LAYER via ;
        RECT 1207.140 3194.680 1207.400 3194.940 ;
        RECT 2900.400 3194.680 2900.660 3194.940 ;
      LAYER met2 ;
        RECT 2900.390 3196.835 2900.670 3197.205 ;
        RECT 2900.460 3194.970 2900.600 3196.835 ;
        RECT 1207.140 3194.650 1207.400 3194.970 ;
        RECT 2900.400 3194.650 2900.660 3194.970 ;
        RECT 1207.200 2600.730 1207.340 3194.650 ;
        RECT 1206.280 2600.590 1207.340 2600.730 ;
        RECT 1204.290 2599.370 1204.570 2600.000 ;
        RECT 1206.280 2599.370 1206.420 2600.590 ;
        RECT 1204.290 2599.230 1206.420 2599.370 ;
        RECT 1204.290 2596.000 1204.570 2599.230 ;
      LAYER via2 ;
        RECT 2900.390 3196.880 2900.670 3197.160 ;
      LAYER met3 ;
        RECT 2900.365 3197.170 2900.695 3197.185 ;
        RECT 2918.000 3197.170 2924.000 3197.620 ;
        RECT 2900.365 3196.870 2924.000 3197.170 ;
        RECT 2900.365 3196.855 2900.695 3196.870 ;
        RECT 2918.000 3196.420 2924.000 3196.870 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1497.460 3429.680 1506.340 3429.820 ;
        RECT 1234.710 3429.480 1235.030 3429.540 ;
        RECT 1497.460 3429.480 1497.600 3429.680 ;
        RECT 1234.710 3429.340 1497.600 3429.480 ;
        RECT 1506.200 3429.480 1506.340 3429.680 ;
        RECT 2762.920 3429.680 2798.940 3429.820 ;
        RECT 2762.920 3429.480 2763.060 3429.680 ;
        RECT 1506.200 3429.340 2763.060 3429.480 ;
        RECT 2798.800 3429.480 2798.940 3429.680 ;
        RECT 2900.370 3429.480 2900.690 3429.540 ;
        RECT 2798.800 3429.340 2900.690 3429.480 ;
        RECT 1234.710 3429.280 1235.030 3429.340 ;
        RECT 2900.370 3429.280 2900.690 3429.340 ;
      LAYER via ;
        RECT 1234.740 3429.280 1235.000 3429.540 ;
        RECT 2900.400 3429.280 2900.660 3429.540 ;
      LAYER met2 ;
        RECT 2900.390 3431.435 2900.670 3431.805 ;
        RECT 2900.460 3429.570 2900.600 3431.435 ;
        RECT 1234.740 3429.250 1235.000 3429.570 ;
        RECT 2900.400 3429.250 2900.660 3429.570 ;
        RECT 1234.800 2600.730 1234.940 3429.250 ;
        RECT 1231.580 2600.590 1234.940 2600.730 ;
        RECT 1230.050 2599.370 1230.330 2600.000 ;
        RECT 1231.580 2599.370 1231.720 2600.590 ;
        RECT 1230.050 2599.230 1231.720 2599.370 ;
        RECT 1230.050 2596.000 1230.330 2599.230 ;
      LAYER via2 ;
        RECT 2900.390 3431.480 2900.670 3431.760 ;
      LAYER met3 ;
        RECT 2900.365 3431.770 2900.695 3431.785 ;
        RECT 2918.000 3431.770 2924.000 3432.220 ;
        RECT 2900.365 3431.470 2924.000 3431.770 ;
        RECT 2900.365 3431.455 2900.695 3431.470 ;
        RECT 2918.000 3431.020 2924.000 3431.470 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1261.925 3381.045 1262.095 3429.155 ;
        RECT 1261.925 3284.485 1262.095 3332.595 ;
        RECT 1261.925 3187.925 1262.095 3236.035 ;
      LAYER mcon ;
        RECT 1261.925 3428.985 1262.095 3429.155 ;
        RECT 1261.925 3332.425 1262.095 3332.595 ;
        RECT 1261.925 3235.865 1262.095 3236.035 ;
      LAYER met1 ;
        RECT 1261.390 3443.080 1261.710 3443.140 ;
        RECT 1262.310 3443.080 1262.630 3443.140 ;
        RECT 1261.390 3442.940 1262.630 3443.080 ;
        RECT 1261.390 3442.880 1261.710 3442.940 ;
        RECT 1262.310 3442.880 1262.630 3442.940 ;
        RECT 1261.865 3429.140 1262.155 3429.185 ;
        RECT 1262.310 3429.140 1262.630 3429.200 ;
        RECT 1261.865 3429.000 1262.630 3429.140 ;
        RECT 1261.865 3428.955 1262.155 3429.000 ;
        RECT 1262.310 3428.940 1262.630 3429.000 ;
        RECT 1261.850 3381.200 1262.170 3381.260 ;
        RECT 1261.655 3381.060 1262.170 3381.200 ;
        RECT 1261.850 3381.000 1262.170 3381.060 ;
        RECT 1261.390 3346.520 1261.710 3346.580 ;
        RECT 1262.310 3346.520 1262.630 3346.580 ;
        RECT 1261.390 3346.380 1262.630 3346.520 ;
        RECT 1261.390 3346.320 1261.710 3346.380 ;
        RECT 1262.310 3346.320 1262.630 3346.380 ;
        RECT 1261.865 3332.580 1262.155 3332.625 ;
        RECT 1262.310 3332.580 1262.630 3332.640 ;
        RECT 1261.865 3332.440 1262.630 3332.580 ;
        RECT 1261.865 3332.395 1262.155 3332.440 ;
        RECT 1262.310 3332.380 1262.630 3332.440 ;
        RECT 1261.850 3284.640 1262.170 3284.700 ;
        RECT 1261.655 3284.500 1262.170 3284.640 ;
        RECT 1261.850 3284.440 1262.170 3284.500 ;
        RECT 1261.390 3249.960 1261.710 3250.020 ;
        RECT 1262.310 3249.960 1262.630 3250.020 ;
        RECT 1261.390 3249.820 1262.630 3249.960 ;
        RECT 1261.390 3249.760 1261.710 3249.820 ;
        RECT 1262.310 3249.760 1262.630 3249.820 ;
        RECT 1261.865 3236.020 1262.155 3236.065 ;
        RECT 1262.310 3236.020 1262.630 3236.080 ;
        RECT 1261.865 3235.880 1262.630 3236.020 ;
        RECT 1261.865 3235.835 1262.155 3235.880 ;
        RECT 1262.310 3235.820 1262.630 3235.880 ;
        RECT 1261.850 3188.080 1262.170 3188.140 ;
        RECT 1261.655 3187.940 1262.170 3188.080 ;
        RECT 1261.850 3187.880 1262.170 3187.940 ;
        RECT 1259.090 2670.600 1259.410 2670.660 ;
        RECT 1261.850 2670.600 1262.170 2670.660 ;
        RECT 1259.090 2670.460 1262.170 2670.600 ;
        RECT 1259.090 2670.400 1259.410 2670.460 ;
        RECT 1261.850 2670.400 1262.170 2670.460 ;
      LAYER via ;
        RECT 1261.420 3442.880 1261.680 3443.140 ;
        RECT 1262.340 3442.880 1262.600 3443.140 ;
        RECT 1262.340 3428.940 1262.600 3429.200 ;
        RECT 1261.880 3381.000 1262.140 3381.260 ;
        RECT 1261.420 3346.320 1261.680 3346.580 ;
        RECT 1262.340 3346.320 1262.600 3346.580 ;
        RECT 1262.340 3332.380 1262.600 3332.640 ;
        RECT 1261.880 3284.440 1262.140 3284.700 ;
        RECT 1261.420 3249.760 1261.680 3250.020 ;
        RECT 1262.340 3249.760 1262.600 3250.020 ;
        RECT 1262.340 3235.820 1262.600 3236.080 ;
        RECT 1261.880 3187.880 1262.140 3188.140 ;
        RECT 1259.120 2670.400 1259.380 2670.660 ;
        RECT 1261.880 2670.400 1262.140 2670.660 ;
      LAYER met2 ;
        RECT 2717.170 3518.000 2717.730 3524.000 ;
        RECT 2717.380 3501.845 2717.520 3518.000 ;
        RECT 1261.870 3501.475 1262.150 3501.845 ;
        RECT 2717.310 3501.475 2717.590 3501.845 ;
        RECT 1261.940 3443.250 1262.080 3501.475 ;
        RECT 1261.480 3443.170 1262.080 3443.250 ;
        RECT 1261.420 3443.110 1262.080 3443.170 ;
        RECT 1261.420 3442.850 1261.680 3443.110 ;
        RECT 1262.340 3442.850 1262.600 3443.170 ;
        RECT 1261.480 3442.695 1261.620 3442.850 ;
        RECT 1262.400 3429.230 1262.540 3442.850 ;
        RECT 1262.340 3428.910 1262.600 3429.230 ;
        RECT 1261.880 3380.970 1262.140 3381.290 ;
        RECT 1261.940 3346.690 1262.080 3380.970 ;
        RECT 1261.480 3346.610 1262.080 3346.690 ;
        RECT 1261.420 3346.550 1262.080 3346.610 ;
        RECT 1261.420 3346.290 1261.680 3346.550 ;
        RECT 1262.340 3346.290 1262.600 3346.610 ;
        RECT 1261.480 3346.135 1261.620 3346.290 ;
        RECT 1262.400 3332.670 1262.540 3346.290 ;
        RECT 1262.340 3332.350 1262.600 3332.670 ;
        RECT 1261.880 3284.410 1262.140 3284.730 ;
        RECT 1261.940 3250.130 1262.080 3284.410 ;
        RECT 1261.480 3250.050 1262.080 3250.130 ;
        RECT 1261.420 3249.990 1262.080 3250.050 ;
        RECT 1261.420 3249.730 1261.680 3249.990 ;
        RECT 1262.340 3249.730 1262.600 3250.050 ;
        RECT 1261.480 3249.575 1261.620 3249.730 ;
        RECT 1262.400 3236.110 1262.540 3249.730 ;
        RECT 1262.340 3235.790 1262.600 3236.110 ;
        RECT 1261.880 3187.850 1262.140 3188.170 ;
        RECT 1261.940 3153.570 1262.080 3187.850 ;
        RECT 1261.480 3153.430 1262.080 3153.570 ;
        RECT 1261.480 3152.890 1261.620 3153.430 ;
        RECT 1261.480 3152.750 1262.080 3152.890 ;
        RECT 1261.940 3105.290 1262.080 3152.750 ;
        RECT 1261.940 3105.150 1262.540 3105.290 ;
        RECT 1262.400 3104.610 1262.540 3105.150 ;
        RECT 1261.940 3104.470 1262.540 3104.610 ;
        RECT 1261.940 3057.010 1262.080 3104.470 ;
        RECT 1261.480 3056.870 1262.080 3057.010 ;
        RECT 1261.480 3056.330 1261.620 3056.870 ;
        RECT 1261.480 3056.190 1262.080 3056.330 ;
        RECT 1261.940 3008.730 1262.080 3056.190 ;
        RECT 1261.940 3008.590 1262.540 3008.730 ;
        RECT 1262.400 3008.050 1262.540 3008.590 ;
        RECT 1261.940 3007.910 1262.540 3008.050 ;
        RECT 1261.940 2960.450 1262.080 3007.910 ;
        RECT 1261.480 2960.310 1262.080 2960.450 ;
        RECT 1261.480 2959.770 1261.620 2960.310 ;
        RECT 1261.480 2959.630 1262.080 2959.770 ;
        RECT 1261.940 2912.170 1262.080 2959.630 ;
        RECT 1261.940 2912.030 1262.540 2912.170 ;
        RECT 1262.400 2911.490 1262.540 2912.030 ;
        RECT 1261.940 2911.350 1262.540 2911.490 ;
        RECT 1261.940 2863.890 1262.080 2911.350 ;
        RECT 1261.480 2863.750 1262.080 2863.890 ;
        RECT 1261.480 2863.210 1261.620 2863.750 ;
        RECT 1261.480 2863.070 1262.080 2863.210 ;
        RECT 1261.940 2815.610 1262.080 2863.070 ;
        RECT 1261.940 2815.470 1262.540 2815.610 ;
        RECT 1262.400 2814.930 1262.540 2815.470 ;
        RECT 1261.940 2814.790 1262.540 2814.930 ;
        RECT 1261.940 2767.330 1262.080 2814.790 ;
        RECT 1261.480 2767.190 1262.080 2767.330 ;
        RECT 1261.480 2766.650 1261.620 2767.190 ;
        RECT 1261.480 2766.510 1262.080 2766.650 ;
        RECT 1261.940 2719.050 1262.080 2766.510 ;
        RECT 1261.940 2718.910 1262.540 2719.050 ;
        RECT 1262.400 2718.370 1262.540 2718.910 ;
        RECT 1261.940 2718.230 1262.540 2718.370 ;
        RECT 1261.940 2670.690 1262.080 2718.230 ;
        RECT 1259.120 2670.370 1259.380 2670.690 ;
        RECT 1261.880 2670.370 1262.140 2670.690 ;
        RECT 1259.180 2642.890 1259.320 2670.370 ;
        RECT 1258.720 2642.750 1259.320 2642.890 ;
        RECT 1258.720 2600.730 1258.860 2642.750 ;
        RECT 1257.340 2600.590 1258.860 2600.730 ;
        RECT 1255.810 2599.370 1256.090 2600.000 ;
        RECT 1257.340 2599.370 1257.480 2600.590 ;
        RECT 1255.810 2599.230 1257.480 2599.370 ;
        RECT 1255.810 2596.000 1256.090 2599.230 ;
      LAYER via2 ;
        RECT 1261.870 3501.520 1262.150 3501.800 ;
        RECT 2717.310 3501.520 2717.590 3501.800 ;
      LAYER met3 ;
        RECT 1261.845 3501.810 1262.175 3501.825 ;
        RECT 2717.285 3501.810 2717.615 3501.825 ;
        RECT 1261.845 3501.510 2717.615 3501.810 ;
        RECT 1261.845 3501.495 1262.175 3501.510 ;
        RECT 2717.285 3501.495 2717.615 3501.510 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1283.010 3502.920 1283.330 3502.980 ;
        RECT 2392.530 3502.920 2392.850 3502.980 ;
        RECT 1283.010 3502.780 2392.850 3502.920 ;
        RECT 1283.010 3502.720 1283.330 3502.780 ;
        RECT 2392.530 3502.720 2392.850 3502.780 ;
      LAYER via ;
        RECT 1283.040 3502.720 1283.300 3502.980 ;
        RECT 2392.560 3502.720 2392.820 3502.980 ;
      LAYER met2 ;
        RECT 2392.410 3518.000 2392.970 3524.000 ;
        RECT 2392.620 3503.010 2392.760 3518.000 ;
        RECT 1283.040 3502.690 1283.300 3503.010 ;
        RECT 2392.560 3502.690 2392.820 3503.010 ;
        RECT 1281.570 2599.370 1281.850 2600.000 ;
        RECT 1283.100 2599.370 1283.240 3502.690 ;
        RECT 1281.570 2599.230 1283.240 2599.370 ;
        RECT 1281.570 2596.000 1281.850 2599.230 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1310.610 3504.620 1310.930 3504.680 ;
        RECT 2068.230 3504.620 2068.550 3504.680 ;
        RECT 1310.610 3504.480 2068.550 3504.620 ;
        RECT 1310.610 3504.420 1310.930 3504.480 ;
        RECT 2068.230 3504.420 2068.550 3504.480 ;
      LAYER via ;
        RECT 1310.640 3504.420 1310.900 3504.680 ;
        RECT 2068.260 3504.420 2068.520 3504.680 ;
      LAYER met2 ;
        RECT 2068.110 3518.000 2068.670 3524.000 ;
        RECT 2068.320 3504.710 2068.460 3518.000 ;
        RECT 1310.640 3504.390 1310.900 3504.710 ;
        RECT 2068.260 3504.390 2068.520 3504.710 ;
        RECT 1310.700 2600.730 1310.840 3504.390 ;
        RECT 1308.860 2600.590 1310.840 2600.730 ;
        RECT 1306.870 2599.370 1307.150 2600.000 ;
        RECT 1308.860 2599.370 1309.000 2600.590 ;
        RECT 1306.870 2599.230 1309.000 2599.370 ;
        RECT 1306.870 2596.000 1307.150 2599.230 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1347.025 3498.345 1347.195 3500.215 ;
        RECT 1337.825 3429.665 1337.995 3443.775 ;
        RECT 1337.825 3414.705 1337.995 3422.355 ;
        RECT 1336.905 3326.305 1337.075 3374.075 ;
        RECT 1337.825 3297.745 1337.995 3325.795 ;
        RECT 1337.365 3229.405 1337.535 3250.995 ;
        RECT 1337.365 3133.185 1337.535 3154.435 ;
        RECT 1336.445 2946.865 1336.615 2960.635 ;
      LAYER mcon ;
        RECT 1347.025 3500.045 1347.195 3500.215 ;
        RECT 1337.825 3443.605 1337.995 3443.775 ;
        RECT 1337.825 3422.185 1337.995 3422.355 ;
        RECT 1336.905 3373.905 1337.075 3374.075 ;
        RECT 1337.825 3325.625 1337.995 3325.795 ;
        RECT 1337.365 3250.825 1337.535 3250.995 ;
        RECT 1337.365 3154.265 1337.535 3154.435 ;
        RECT 1336.445 2960.465 1336.615 2960.635 ;
      LAYER met1 ;
        RECT 1346.965 3500.200 1347.255 3500.245 ;
        RECT 1743.930 3500.200 1744.250 3500.260 ;
        RECT 1346.965 3500.060 1744.250 3500.200 ;
        RECT 1346.965 3500.015 1347.255 3500.060 ;
        RECT 1743.930 3500.000 1744.250 3500.060 ;
        RECT 1338.210 3498.500 1338.530 3498.560 ;
        RECT 1346.965 3498.500 1347.255 3498.545 ;
        RECT 1338.210 3498.360 1347.255 3498.500 ;
        RECT 1338.210 3498.300 1338.530 3498.360 ;
        RECT 1346.965 3498.315 1347.255 3498.360 ;
        RECT 1337.765 3443.760 1338.055 3443.805 ;
        RECT 1338.210 3443.760 1338.530 3443.820 ;
        RECT 1337.765 3443.620 1338.530 3443.760 ;
        RECT 1337.765 3443.575 1338.055 3443.620 ;
        RECT 1338.210 3443.560 1338.530 3443.620 ;
        RECT 1337.750 3429.820 1338.070 3429.880 ;
        RECT 1337.555 3429.680 1338.070 3429.820 ;
        RECT 1337.750 3429.620 1338.070 3429.680 ;
        RECT 1337.750 3422.340 1338.070 3422.400 ;
        RECT 1337.555 3422.200 1338.070 3422.340 ;
        RECT 1337.750 3422.140 1338.070 3422.200 ;
        RECT 1337.765 3414.860 1338.055 3414.905 ;
        RECT 1338.210 3414.860 1338.530 3414.920 ;
        RECT 1337.765 3414.720 1338.530 3414.860 ;
        RECT 1337.765 3414.675 1338.055 3414.720 ;
        RECT 1338.210 3414.660 1338.530 3414.720 ;
        RECT 1336.845 3374.060 1337.135 3374.105 ;
        RECT 1338.210 3374.060 1338.530 3374.120 ;
        RECT 1336.845 3373.920 1338.530 3374.060 ;
        RECT 1336.845 3373.875 1337.135 3373.920 ;
        RECT 1338.210 3373.860 1338.530 3373.920 ;
        RECT 1336.830 3326.460 1337.150 3326.520 ;
        RECT 1336.635 3326.320 1337.150 3326.460 ;
        RECT 1336.830 3326.260 1337.150 3326.320 ;
        RECT 1336.830 3325.780 1337.150 3325.840 ;
        RECT 1337.765 3325.780 1338.055 3325.825 ;
        RECT 1336.830 3325.640 1338.055 3325.780 ;
        RECT 1336.830 3325.580 1337.150 3325.640 ;
        RECT 1337.765 3325.595 1338.055 3325.640 ;
        RECT 1337.750 3297.900 1338.070 3297.960 ;
        RECT 1337.555 3297.760 1338.070 3297.900 ;
        RECT 1337.750 3297.700 1338.070 3297.760 ;
        RECT 1337.305 3250.980 1337.595 3251.025 ;
        RECT 1337.750 3250.980 1338.070 3251.040 ;
        RECT 1337.305 3250.840 1338.070 3250.980 ;
        RECT 1337.305 3250.795 1337.595 3250.840 ;
        RECT 1337.750 3250.780 1338.070 3250.840 ;
        RECT 1337.290 3229.560 1337.610 3229.620 ;
        RECT 1337.095 3229.420 1337.610 3229.560 ;
        RECT 1337.290 3229.360 1337.610 3229.420 ;
        RECT 1337.305 3154.420 1337.595 3154.465 ;
        RECT 1337.750 3154.420 1338.070 3154.480 ;
        RECT 1337.305 3154.280 1338.070 3154.420 ;
        RECT 1337.305 3154.235 1337.595 3154.280 ;
        RECT 1337.750 3154.220 1338.070 3154.280 ;
        RECT 1337.290 3133.340 1337.610 3133.400 ;
        RECT 1337.095 3133.200 1337.610 3133.340 ;
        RECT 1337.290 3133.140 1337.610 3133.200 ;
        RECT 1337.290 3115.660 1337.610 3115.720 ;
        RECT 1337.750 3115.660 1338.070 3115.720 ;
        RECT 1337.290 3115.520 1338.070 3115.660 ;
        RECT 1337.290 3115.460 1337.610 3115.520 ;
        RECT 1337.750 3115.460 1338.070 3115.520 ;
        RECT 1336.385 2960.620 1336.675 2960.665 ;
        RECT 1336.830 2960.620 1337.150 2960.680 ;
        RECT 1336.385 2960.480 1337.150 2960.620 ;
        RECT 1336.385 2960.435 1336.675 2960.480 ;
        RECT 1336.830 2960.420 1337.150 2960.480 ;
        RECT 1336.370 2947.020 1336.690 2947.080 ;
        RECT 1336.175 2946.880 1336.690 2947.020 ;
        RECT 1336.370 2946.820 1336.690 2946.880 ;
        RECT 1336.370 2911.800 1336.690 2912.060 ;
        RECT 1336.460 2911.320 1336.600 2911.800 ;
        RECT 1336.830 2911.320 1337.150 2911.380 ;
        RECT 1336.460 2911.180 1337.150 2911.320 ;
        RECT 1336.830 2911.120 1337.150 2911.180 ;
        RECT 1336.830 2814.760 1337.150 2814.820 ;
        RECT 1337.750 2814.760 1338.070 2814.820 ;
        RECT 1336.830 2814.620 1338.070 2814.760 ;
        RECT 1336.830 2814.560 1337.150 2814.620 ;
        RECT 1337.750 2814.560 1338.070 2814.620 ;
        RECT 1335.910 2656.660 1336.230 2656.720 ;
        RECT 1337.750 2656.660 1338.070 2656.720 ;
        RECT 1335.910 2656.520 1338.070 2656.660 ;
        RECT 1335.910 2656.460 1336.230 2656.520 ;
        RECT 1337.750 2656.460 1338.070 2656.520 ;
      LAYER via ;
        RECT 1743.960 3500.000 1744.220 3500.260 ;
        RECT 1338.240 3498.300 1338.500 3498.560 ;
        RECT 1338.240 3443.560 1338.500 3443.820 ;
        RECT 1337.780 3429.620 1338.040 3429.880 ;
        RECT 1337.780 3422.140 1338.040 3422.400 ;
        RECT 1338.240 3414.660 1338.500 3414.920 ;
        RECT 1338.240 3373.860 1338.500 3374.120 ;
        RECT 1336.860 3326.260 1337.120 3326.520 ;
        RECT 1336.860 3325.580 1337.120 3325.840 ;
        RECT 1337.780 3297.700 1338.040 3297.960 ;
        RECT 1337.780 3250.780 1338.040 3251.040 ;
        RECT 1337.320 3229.360 1337.580 3229.620 ;
        RECT 1337.780 3154.220 1338.040 3154.480 ;
        RECT 1337.320 3133.140 1337.580 3133.400 ;
        RECT 1337.320 3115.460 1337.580 3115.720 ;
        RECT 1337.780 3115.460 1338.040 3115.720 ;
        RECT 1336.860 2960.420 1337.120 2960.680 ;
        RECT 1336.400 2946.820 1336.660 2947.080 ;
        RECT 1336.400 2911.800 1336.660 2912.060 ;
        RECT 1336.860 2911.120 1337.120 2911.380 ;
        RECT 1336.860 2814.560 1337.120 2814.820 ;
        RECT 1337.780 2814.560 1338.040 2814.820 ;
        RECT 1335.940 2656.460 1336.200 2656.720 ;
        RECT 1337.780 2656.460 1338.040 2656.720 ;
      LAYER met2 ;
        RECT 1743.810 3518.000 1744.370 3524.000 ;
        RECT 1744.020 3500.290 1744.160 3518.000 ;
        RECT 1743.960 3499.970 1744.220 3500.290 ;
        RECT 1338.240 3498.270 1338.500 3498.590 ;
        RECT 1338.300 3443.850 1338.440 3498.270 ;
        RECT 1338.240 3443.530 1338.500 3443.850 ;
        RECT 1337.780 3429.590 1338.040 3429.910 ;
        RECT 1337.840 3422.430 1337.980 3429.590 ;
        RECT 1337.780 3422.110 1338.040 3422.430 ;
        RECT 1338.240 3414.630 1338.500 3414.950 ;
        RECT 1338.300 3374.150 1338.440 3414.630 ;
        RECT 1338.240 3373.830 1338.500 3374.150 ;
        RECT 1336.860 3326.230 1337.120 3326.550 ;
        RECT 1336.920 3325.870 1337.060 3326.230 ;
        RECT 1336.860 3325.550 1337.120 3325.870 ;
        RECT 1337.780 3297.670 1338.040 3297.990 ;
        RECT 1337.840 3251.070 1337.980 3297.670 ;
        RECT 1337.780 3250.750 1338.040 3251.070 ;
        RECT 1337.320 3229.330 1337.580 3229.650 ;
        RECT 1337.380 3229.165 1337.520 3229.330 ;
        RECT 1337.310 3228.795 1337.590 3229.165 ;
        RECT 1337.770 3200.915 1338.050 3201.285 ;
        RECT 1337.840 3154.510 1337.980 3200.915 ;
        RECT 1337.780 3154.190 1338.040 3154.510 ;
        RECT 1337.320 3133.110 1337.580 3133.430 ;
        RECT 1337.380 3115.750 1337.520 3133.110 ;
        RECT 1337.320 3115.430 1337.580 3115.750 ;
        RECT 1337.780 3115.430 1338.040 3115.750 ;
        RECT 1337.840 3057.010 1337.980 3115.430 ;
        RECT 1337.840 3056.870 1338.440 3057.010 ;
        RECT 1338.300 3056.330 1338.440 3056.870 ;
        RECT 1337.380 3056.190 1338.440 3056.330 ;
        RECT 1337.380 3008.730 1337.520 3056.190 ;
        RECT 1336.920 3008.590 1337.520 3008.730 ;
        RECT 1336.920 2960.710 1337.060 3008.590 ;
        RECT 1336.860 2960.390 1337.120 2960.710 ;
        RECT 1336.400 2946.790 1336.660 2947.110 ;
        RECT 1336.460 2912.090 1336.600 2946.790 ;
        RECT 1336.400 2911.770 1336.660 2912.090 ;
        RECT 1336.860 2911.090 1337.120 2911.410 ;
        RECT 1336.920 2891.205 1337.060 2911.090 ;
        RECT 1336.850 2890.835 1337.130 2891.205 ;
        RECT 1337.770 2890.835 1338.050 2891.205 ;
        RECT 1337.840 2842.980 1337.980 2890.835 ;
        RECT 1336.920 2842.925 1337.980 2842.980 ;
        RECT 1336.850 2842.840 1338.050 2842.925 ;
        RECT 1336.850 2842.555 1337.130 2842.840 ;
        RECT 1337.770 2842.555 1338.050 2842.840 ;
        RECT 1337.840 2814.850 1337.980 2842.555 ;
        RECT 1336.860 2814.530 1337.120 2814.850 ;
        RECT 1337.780 2814.530 1338.040 2814.850 ;
        RECT 1336.920 2766.650 1337.060 2814.530 ;
        RECT 1336.920 2766.510 1337.520 2766.650 ;
        RECT 1337.380 2719.050 1337.520 2766.510 ;
        RECT 1337.380 2718.910 1337.980 2719.050 ;
        RECT 1337.840 2656.750 1337.980 2718.910 ;
        RECT 1335.940 2656.605 1336.200 2656.750 ;
        RECT 1335.010 2656.235 1335.290 2656.605 ;
        RECT 1335.930 2656.235 1336.210 2656.605 ;
        RECT 1337.780 2656.430 1338.040 2656.750 ;
        RECT 1332.630 2599.370 1332.910 2600.000 ;
        RECT 1335.080 2599.370 1335.220 2656.235 ;
        RECT 1332.630 2599.230 1335.220 2599.370 ;
        RECT 1332.630 2596.000 1332.910 2599.230 ;
      LAYER via2 ;
        RECT 1337.310 3228.840 1337.590 3229.120 ;
        RECT 1337.770 3200.960 1338.050 3201.240 ;
        RECT 1336.850 2890.880 1337.130 2891.160 ;
        RECT 1337.770 2890.880 1338.050 2891.160 ;
        RECT 1336.850 2842.600 1337.130 2842.880 ;
        RECT 1337.770 2842.600 1338.050 2842.880 ;
        RECT 1335.010 2656.280 1335.290 2656.560 ;
        RECT 1335.930 2656.280 1336.210 2656.560 ;
      LAYER met3 ;
        RECT 1337.285 3229.140 1337.615 3229.145 ;
        RECT 1337.030 3229.130 1337.615 3229.140 ;
        RECT 1337.030 3228.830 1337.840 3229.130 ;
        RECT 1337.030 3228.820 1337.615 3228.830 ;
        RECT 1337.285 3228.815 1337.615 3228.820 ;
        RECT 1337.030 3201.250 1337.410 3201.260 ;
        RECT 1337.745 3201.250 1338.075 3201.265 ;
        RECT 1337.030 3200.950 1338.075 3201.250 ;
        RECT 1337.030 3200.940 1337.410 3200.950 ;
        RECT 1337.745 3200.935 1338.075 3200.950 ;
        RECT 1336.825 2891.170 1337.155 2891.185 ;
        RECT 1337.745 2891.170 1338.075 2891.185 ;
        RECT 1336.825 2890.870 1338.075 2891.170 ;
        RECT 1336.825 2890.855 1337.155 2890.870 ;
        RECT 1337.745 2890.855 1338.075 2890.870 ;
        RECT 1336.825 2842.890 1337.155 2842.905 ;
        RECT 1337.745 2842.890 1338.075 2842.905 ;
        RECT 1336.825 2842.590 1338.075 2842.890 ;
        RECT 1336.825 2842.575 1337.155 2842.590 ;
        RECT 1337.745 2842.575 1338.075 2842.590 ;
        RECT 1334.985 2656.570 1335.315 2656.585 ;
        RECT 1335.905 2656.570 1336.235 2656.585 ;
        RECT 1334.985 2656.270 1336.235 2656.570 ;
        RECT 1334.985 2656.255 1335.315 2656.270 ;
        RECT 1335.905 2656.255 1336.235 2656.270 ;
      LAYER via3 ;
        RECT 1337.060 3228.820 1337.380 3229.140 ;
        RECT 1337.060 3200.940 1337.380 3201.260 ;
      LAYER met4 ;
        RECT 1337.055 3228.815 1337.385 3229.145 ;
        RECT 1337.070 3201.265 1337.370 3228.815 ;
        RECT 1337.055 3200.935 1337.385 3201.265 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1358.910 3498.500 1359.230 3498.560 ;
        RECT 1419.170 3498.500 1419.490 3498.560 ;
        RECT 1358.910 3498.360 1419.490 3498.500 ;
        RECT 1358.910 3498.300 1359.230 3498.360 ;
        RECT 1419.170 3498.300 1419.490 3498.360 ;
      LAYER via ;
        RECT 1358.940 3498.300 1359.200 3498.560 ;
        RECT 1419.200 3498.300 1419.460 3498.560 ;
      LAYER met2 ;
        RECT 1419.050 3518.000 1419.610 3524.000 ;
        RECT 1419.260 3498.590 1419.400 3518.000 ;
        RECT 1358.940 3498.270 1359.200 3498.590 ;
        RECT 1419.200 3498.270 1419.460 3498.590 ;
        RECT 1358.390 2599.370 1358.670 2600.000 ;
        RECT 1359.000 2599.370 1359.140 3498.270 ;
        RECT 1358.390 2599.230 1359.140 2599.370 ;
        RECT 1358.390 2596.000 1358.670 2599.230 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 897.145 2590.885 897.315 2597.855 ;
      LAYER mcon ;
        RECT 897.145 2597.685 897.315 2597.855 ;
      LAYER met1 ;
        RECT 897.070 2597.840 897.390 2597.900 ;
        RECT 896.875 2597.700 897.390 2597.840 ;
        RECT 897.070 2597.640 897.390 2597.700 ;
        RECT 897.085 2591.040 897.375 2591.085 ;
        RECT 2901.750 2591.040 2902.070 2591.100 ;
        RECT 897.085 2590.900 2902.070 2591.040 ;
        RECT 897.085 2590.855 897.375 2590.900 ;
        RECT 2901.750 2590.840 2902.070 2590.900 ;
      LAYER via ;
        RECT 897.100 2597.640 897.360 2597.900 ;
        RECT 2901.780 2590.840 2902.040 2591.100 ;
      LAYER met2 ;
        RECT 896.550 2598.010 896.830 2600.000 ;
        RECT 896.550 2597.930 897.300 2598.010 ;
        RECT 896.550 2597.870 897.360 2597.930 ;
        RECT 896.550 2596.000 896.830 2597.870 ;
        RECT 897.100 2597.610 897.360 2597.870 ;
        RECT 2901.780 2590.810 2902.040 2591.130 ;
        RECT 2901.840 381.325 2901.980 2590.810 ;
        RECT 2901.770 380.955 2902.050 381.325 ;
      LAYER via2 ;
        RECT 2901.770 381.000 2902.050 381.280 ;
      LAYER met3 ;
        RECT 2901.745 381.290 2902.075 381.305 ;
        RECT 2918.000 381.290 2924.000 381.740 ;
        RECT 2901.745 380.990 2924.000 381.290 ;
        RECT 2901.745 380.975 2902.075 380.990 ;
        RECT 2918.000 380.540 2924.000 380.990 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1380.605 3284.485 1380.775 3332.595 ;
        RECT 1381.065 2959.785 1381.235 2994.635 ;
        RECT 1381.065 2911.165 1381.235 2946.355 ;
      LAYER mcon ;
        RECT 1380.605 3332.425 1380.775 3332.595 ;
        RECT 1381.065 2994.465 1381.235 2994.635 ;
        RECT 1381.065 2946.185 1381.235 2946.355 ;
      LAYER met1 ;
        RECT 1094.870 3499.180 1095.190 3499.240 ;
        RECT 1380.070 3499.180 1380.390 3499.240 ;
        RECT 1094.870 3499.040 1380.390 3499.180 ;
        RECT 1094.870 3498.980 1095.190 3499.040 ;
        RECT 1380.070 3498.980 1380.390 3499.040 ;
        RECT 1380.070 3415.880 1380.390 3415.940 ;
        RECT 1380.990 3415.880 1381.310 3415.940 ;
        RECT 1380.070 3415.740 1381.310 3415.880 ;
        RECT 1380.070 3415.680 1380.390 3415.740 ;
        RECT 1380.990 3415.680 1381.310 3415.740 ;
        RECT 1380.070 3346.520 1380.390 3346.580 ;
        RECT 1380.990 3346.520 1381.310 3346.580 ;
        RECT 1380.070 3346.380 1381.310 3346.520 ;
        RECT 1380.070 3346.320 1380.390 3346.380 ;
        RECT 1380.990 3346.320 1381.310 3346.380 ;
        RECT 1380.545 3332.580 1380.835 3332.625 ;
        RECT 1380.990 3332.580 1381.310 3332.640 ;
        RECT 1380.545 3332.440 1381.310 3332.580 ;
        RECT 1380.545 3332.395 1380.835 3332.440 ;
        RECT 1380.990 3332.380 1381.310 3332.440 ;
        RECT 1380.530 3284.640 1380.850 3284.700 ;
        RECT 1380.335 3284.500 1380.850 3284.640 ;
        RECT 1380.530 3284.440 1380.850 3284.500 ;
        RECT 1380.070 3222.420 1380.390 3222.480 ;
        RECT 1380.990 3222.420 1381.310 3222.480 ;
        RECT 1380.070 3222.280 1381.310 3222.420 ;
        RECT 1380.070 3222.220 1380.390 3222.280 ;
        RECT 1380.990 3222.220 1381.310 3222.280 ;
        RECT 1380.070 3056.840 1380.390 3056.900 ;
        RECT 1380.990 3056.840 1381.310 3056.900 ;
        RECT 1380.070 3056.700 1381.310 3056.840 ;
        RECT 1380.070 3056.640 1380.390 3056.700 ;
        RECT 1380.990 3056.640 1381.310 3056.700 ;
        RECT 1380.530 3008.700 1380.850 3008.960 ;
        RECT 1380.620 3008.560 1380.760 3008.700 ;
        RECT 1380.990 3008.560 1381.310 3008.620 ;
        RECT 1380.620 3008.420 1381.310 3008.560 ;
        RECT 1380.990 3008.360 1381.310 3008.420 ;
        RECT 1380.990 2994.620 1381.310 2994.680 ;
        RECT 1380.795 2994.480 1381.310 2994.620 ;
        RECT 1380.990 2994.420 1381.310 2994.480 ;
        RECT 1380.990 2959.940 1381.310 2960.000 ;
        RECT 1380.795 2959.800 1381.310 2959.940 ;
        RECT 1380.990 2959.740 1381.310 2959.800 ;
        RECT 1380.990 2946.340 1381.310 2946.400 ;
        RECT 1380.795 2946.200 1381.310 2946.340 ;
        RECT 1380.990 2946.140 1381.310 2946.200 ;
        RECT 1380.990 2911.320 1381.310 2911.380 ;
        RECT 1380.795 2911.180 1381.310 2911.320 ;
        RECT 1380.990 2911.120 1381.310 2911.180 ;
        RECT 1380.070 2863.720 1380.390 2863.780 ;
        RECT 1380.990 2863.720 1381.310 2863.780 ;
        RECT 1380.070 2863.580 1381.310 2863.720 ;
        RECT 1380.070 2863.520 1380.390 2863.580 ;
        RECT 1380.990 2863.520 1381.310 2863.580 ;
        RECT 1380.070 2753.220 1380.390 2753.280 ;
        RECT 1380.530 2753.220 1380.850 2753.280 ;
        RECT 1380.070 2753.080 1380.850 2753.220 ;
        RECT 1380.070 2753.020 1380.390 2753.080 ;
        RECT 1380.530 2753.020 1380.850 2753.080 ;
        RECT 1381.450 2698.140 1381.770 2698.200 ;
        RECT 1381.910 2698.140 1382.230 2698.200 ;
        RECT 1381.450 2698.000 1382.230 2698.140 ;
        RECT 1381.450 2697.940 1381.770 2698.000 ;
        RECT 1381.910 2697.940 1382.230 2698.000 ;
        RECT 1381.450 2656.660 1381.770 2656.720 ;
        RECT 1382.830 2656.660 1383.150 2656.720 ;
        RECT 1381.450 2656.520 1383.150 2656.660 ;
        RECT 1381.450 2656.460 1381.770 2656.520 ;
        RECT 1382.830 2656.460 1383.150 2656.520 ;
        RECT 1381.910 2631.840 1382.230 2631.900 ;
        RECT 1382.830 2631.840 1383.150 2631.900 ;
        RECT 1381.910 2631.700 1383.150 2631.840 ;
        RECT 1381.910 2631.640 1382.230 2631.700 ;
        RECT 1382.830 2631.640 1383.150 2631.700 ;
      LAYER via ;
        RECT 1094.900 3498.980 1095.160 3499.240 ;
        RECT 1380.100 3498.980 1380.360 3499.240 ;
        RECT 1380.100 3415.680 1380.360 3415.940 ;
        RECT 1381.020 3415.680 1381.280 3415.940 ;
        RECT 1380.100 3346.320 1380.360 3346.580 ;
        RECT 1381.020 3346.320 1381.280 3346.580 ;
        RECT 1381.020 3332.380 1381.280 3332.640 ;
        RECT 1380.560 3284.440 1380.820 3284.700 ;
        RECT 1380.100 3222.220 1380.360 3222.480 ;
        RECT 1381.020 3222.220 1381.280 3222.480 ;
        RECT 1380.100 3056.640 1380.360 3056.900 ;
        RECT 1381.020 3056.640 1381.280 3056.900 ;
        RECT 1380.560 3008.700 1380.820 3008.960 ;
        RECT 1381.020 3008.360 1381.280 3008.620 ;
        RECT 1381.020 2994.420 1381.280 2994.680 ;
        RECT 1381.020 2959.740 1381.280 2960.000 ;
        RECT 1381.020 2946.140 1381.280 2946.400 ;
        RECT 1381.020 2911.120 1381.280 2911.380 ;
        RECT 1380.100 2863.520 1380.360 2863.780 ;
        RECT 1381.020 2863.520 1381.280 2863.780 ;
        RECT 1380.100 2753.020 1380.360 2753.280 ;
        RECT 1380.560 2753.020 1380.820 2753.280 ;
        RECT 1381.480 2697.940 1381.740 2698.200 ;
        RECT 1381.940 2697.940 1382.200 2698.200 ;
        RECT 1381.480 2656.460 1381.740 2656.720 ;
        RECT 1382.860 2656.460 1383.120 2656.720 ;
        RECT 1381.940 2631.640 1382.200 2631.900 ;
        RECT 1382.860 2631.640 1383.120 2631.900 ;
      LAYER met2 ;
        RECT 1094.750 3518.000 1095.310 3524.000 ;
        RECT 1094.960 3499.270 1095.100 3518.000 ;
        RECT 1094.900 3498.950 1095.160 3499.270 ;
        RECT 1380.100 3498.950 1380.360 3499.270 ;
        RECT 1380.160 3463.650 1380.300 3498.950 ;
        RECT 1380.160 3463.510 1381.220 3463.650 ;
        RECT 1381.080 3415.970 1381.220 3463.510 ;
        RECT 1380.100 3415.650 1380.360 3415.970 ;
        RECT 1381.020 3415.650 1381.280 3415.970 ;
        RECT 1380.160 3346.610 1380.300 3415.650 ;
        RECT 1380.100 3346.290 1380.360 3346.610 ;
        RECT 1381.020 3346.290 1381.280 3346.610 ;
        RECT 1381.080 3332.670 1381.220 3346.290 ;
        RECT 1381.020 3332.350 1381.280 3332.670 ;
        RECT 1380.560 3284.410 1380.820 3284.730 ;
        RECT 1380.620 3250.130 1380.760 3284.410 ;
        RECT 1380.620 3249.990 1381.220 3250.130 ;
        RECT 1381.080 3222.510 1381.220 3249.990 ;
        RECT 1380.100 3222.190 1380.360 3222.510 ;
        RECT 1381.020 3222.190 1381.280 3222.510 ;
        RECT 1380.160 3201.170 1380.300 3222.190 ;
        RECT 1380.160 3201.030 1380.760 3201.170 ;
        RECT 1380.620 3153.570 1380.760 3201.030 ;
        RECT 1380.620 3153.430 1381.220 3153.570 ;
        RECT 1381.080 3056.930 1381.220 3153.430 ;
        RECT 1380.100 3056.610 1380.360 3056.930 ;
        RECT 1381.020 3056.610 1381.280 3056.930 ;
        RECT 1380.160 3056.330 1380.300 3056.610 ;
        RECT 1380.160 3056.190 1380.760 3056.330 ;
        RECT 1380.620 3008.990 1380.760 3056.190 ;
        RECT 1380.560 3008.670 1380.820 3008.990 ;
        RECT 1381.020 3008.330 1381.280 3008.650 ;
        RECT 1381.080 2994.710 1381.220 3008.330 ;
        RECT 1381.020 2994.390 1381.280 2994.710 ;
        RECT 1381.020 2959.710 1381.280 2960.030 ;
        RECT 1381.080 2946.430 1381.220 2959.710 ;
        RECT 1381.020 2946.110 1381.280 2946.430 ;
        RECT 1381.020 2911.090 1381.280 2911.410 ;
        RECT 1381.080 2863.810 1381.220 2911.090 ;
        RECT 1380.100 2863.490 1380.360 2863.810 ;
        RECT 1381.020 2863.490 1381.280 2863.810 ;
        RECT 1380.160 2863.210 1380.300 2863.490 ;
        RECT 1380.160 2863.070 1380.760 2863.210 ;
        RECT 1380.620 2815.610 1380.760 2863.070 ;
        RECT 1380.620 2815.470 1381.220 2815.610 ;
        RECT 1381.080 2801.330 1381.220 2815.470 ;
        RECT 1380.620 2801.190 1381.220 2801.330 ;
        RECT 1380.620 2753.310 1380.760 2801.190 ;
        RECT 1380.100 2753.165 1380.360 2753.310 ;
        RECT 1380.090 2752.795 1380.370 2753.165 ;
        RECT 1380.560 2752.990 1380.820 2753.310 ;
        RECT 1382.390 2752.795 1382.670 2753.165 ;
        RECT 1382.460 2746.250 1382.600 2752.795 ;
        RECT 1382.000 2746.110 1382.600 2746.250 ;
        RECT 1382.000 2698.230 1382.140 2746.110 ;
        RECT 1381.480 2697.910 1381.740 2698.230 ;
        RECT 1381.940 2697.910 1382.200 2698.230 ;
        RECT 1381.540 2656.750 1381.680 2697.910 ;
        RECT 1381.480 2656.430 1381.740 2656.750 ;
        RECT 1382.860 2656.430 1383.120 2656.750 ;
        RECT 1382.920 2631.930 1383.060 2656.430 ;
        RECT 1381.940 2631.610 1382.200 2631.930 ;
        RECT 1382.860 2631.610 1383.120 2631.930 ;
        RECT 1382.000 2600.730 1382.140 2631.610 ;
        RECT 1382.000 2600.590 1383.060 2600.730 ;
        RECT 1382.920 2600.050 1383.060 2600.590 ;
        RECT 1382.920 2600.000 1384.370 2600.050 ;
        RECT 1382.920 2599.910 1384.430 2600.000 ;
        RECT 1384.150 2596.000 1384.430 2599.910 ;
      LAYER via2 ;
        RECT 1380.090 2752.840 1380.370 2753.120 ;
        RECT 1382.390 2752.840 1382.670 2753.120 ;
      LAYER met3 ;
        RECT 1380.065 2753.130 1380.395 2753.145 ;
        RECT 1382.365 2753.130 1382.695 2753.145 ;
        RECT 1380.065 2752.830 1382.695 2753.130 ;
        RECT 1380.065 2752.815 1380.395 2752.830 ;
        RECT 1382.365 2752.815 1382.695 2752.830 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 770.570 3500.880 770.890 3500.940 ;
        RECT 1407.670 3500.880 1407.990 3500.940 ;
        RECT 770.570 3500.740 1407.990 3500.880 ;
        RECT 770.570 3500.680 770.890 3500.740 ;
        RECT 1407.670 3500.680 1407.990 3500.740 ;
      LAYER via ;
        RECT 770.600 3500.680 770.860 3500.940 ;
        RECT 1407.700 3500.680 1407.960 3500.940 ;
      LAYER met2 ;
        RECT 770.450 3518.000 771.010 3524.000 ;
        RECT 770.660 3500.970 770.800 3518.000 ;
        RECT 770.600 3500.650 770.860 3500.970 ;
        RECT 1407.700 3500.650 1407.960 3500.970 ;
        RECT 1407.760 2600.050 1407.900 3500.650 ;
        RECT 1407.760 2600.000 1409.670 2600.050 ;
        RECT 1407.760 2599.910 1409.730 2600.000 ;
        RECT 1409.450 2596.000 1409.730 2599.910 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1435.805 3441.565 1435.975 3477.435 ;
        RECT 1435.805 3332.765 1435.975 3380.875 ;
        RECT 1435.805 2994.805 1435.975 3042.915 ;
        RECT 1435.805 2656.505 1435.975 2670.615 ;
      LAYER mcon ;
        RECT 1435.805 3477.265 1435.975 3477.435 ;
        RECT 1435.805 3380.705 1435.975 3380.875 ;
        RECT 1435.805 3042.745 1435.975 3042.915 ;
        RECT 1435.805 2670.445 1435.975 2670.615 ;
      LAYER met1 ;
        RECT 445.810 3503.940 446.130 3504.000 ;
        RECT 1436.190 3503.940 1436.510 3504.000 ;
        RECT 445.810 3503.800 1436.510 3503.940 ;
        RECT 445.810 3503.740 446.130 3503.800 ;
        RECT 1436.190 3503.740 1436.510 3503.800 ;
        RECT 1435.745 3477.420 1436.035 3477.465 ;
        RECT 1436.190 3477.420 1436.510 3477.480 ;
        RECT 1435.745 3477.280 1436.510 3477.420 ;
        RECT 1435.745 3477.235 1436.035 3477.280 ;
        RECT 1436.190 3477.220 1436.510 3477.280 ;
        RECT 1435.730 3441.720 1436.050 3441.780 ;
        RECT 1435.535 3441.580 1436.050 3441.720 ;
        RECT 1435.730 3441.520 1436.050 3441.580 ;
        RECT 1435.745 3380.860 1436.035 3380.905 ;
        RECT 1436.190 3380.860 1436.510 3380.920 ;
        RECT 1435.745 3380.720 1436.510 3380.860 ;
        RECT 1435.745 3380.675 1436.035 3380.720 ;
        RECT 1436.190 3380.660 1436.510 3380.720 ;
        RECT 1435.730 3332.920 1436.050 3332.980 ;
        RECT 1435.535 3332.780 1436.050 3332.920 ;
        RECT 1435.730 3332.720 1436.050 3332.780 ;
        RECT 1436.190 3249.420 1436.510 3249.680 ;
        RECT 1436.280 3249.000 1436.420 3249.420 ;
        RECT 1436.190 3248.740 1436.510 3249.000 ;
        RECT 1435.270 3153.400 1435.590 3153.460 ;
        RECT 1436.190 3153.400 1436.510 3153.460 ;
        RECT 1435.270 3153.260 1436.510 3153.400 ;
        RECT 1435.270 3153.200 1435.590 3153.260 ;
        RECT 1436.190 3153.200 1436.510 3153.260 ;
        RECT 1435.270 3056.840 1435.590 3056.900 ;
        RECT 1436.190 3056.840 1436.510 3056.900 ;
        RECT 1435.270 3056.700 1436.510 3056.840 ;
        RECT 1435.270 3056.640 1435.590 3056.700 ;
        RECT 1436.190 3056.640 1436.510 3056.700 ;
        RECT 1435.730 3042.900 1436.050 3042.960 ;
        RECT 1435.535 3042.760 1436.050 3042.900 ;
        RECT 1435.730 3042.700 1436.050 3042.760 ;
        RECT 1435.745 2994.960 1436.035 2995.005 ;
        RECT 1436.190 2994.960 1436.510 2995.020 ;
        RECT 1435.745 2994.820 1436.510 2994.960 ;
        RECT 1435.745 2994.775 1436.035 2994.820 ;
        RECT 1436.190 2994.760 1436.510 2994.820 ;
        RECT 1435.270 2863.720 1435.590 2863.780 ;
        RECT 1436.190 2863.720 1436.510 2863.780 ;
        RECT 1435.270 2863.580 1436.510 2863.720 ;
        RECT 1435.270 2863.520 1435.590 2863.580 ;
        RECT 1436.190 2863.520 1436.510 2863.580 ;
        RECT 1435.270 2753.220 1435.590 2753.280 ;
        RECT 1435.730 2753.220 1436.050 2753.280 ;
        RECT 1435.270 2753.080 1436.050 2753.220 ;
        RECT 1435.270 2753.020 1435.590 2753.080 ;
        RECT 1435.730 2753.020 1436.050 2753.080 ;
        RECT 1435.270 2704.600 1435.590 2704.660 ;
        RECT 1436.190 2704.600 1436.510 2704.660 ;
        RECT 1435.270 2704.460 1436.510 2704.600 ;
        RECT 1435.270 2704.400 1435.590 2704.460 ;
        RECT 1436.190 2704.400 1436.510 2704.460 ;
        RECT 1435.745 2670.600 1436.035 2670.645 ;
        RECT 1436.650 2670.600 1436.970 2670.660 ;
        RECT 1435.745 2670.460 1436.970 2670.600 ;
        RECT 1435.745 2670.415 1436.035 2670.460 ;
        RECT 1436.650 2670.400 1436.970 2670.460 ;
        RECT 1435.730 2656.660 1436.050 2656.720 ;
        RECT 1435.535 2656.520 1436.050 2656.660 ;
        RECT 1435.730 2656.460 1436.050 2656.520 ;
      LAYER via ;
        RECT 445.840 3503.740 446.100 3504.000 ;
        RECT 1436.220 3503.740 1436.480 3504.000 ;
        RECT 1436.220 3477.220 1436.480 3477.480 ;
        RECT 1435.760 3441.520 1436.020 3441.780 ;
        RECT 1436.220 3380.660 1436.480 3380.920 ;
        RECT 1435.760 3332.720 1436.020 3332.980 ;
        RECT 1436.220 3249.420 1436.480 3249.680 ;
        RECT 1436.220 3248.740 1436.480 3249.000 ;
        RECT 1435.300 3153.200 1435.560 3153.460 ;
        RECT 1436.220 3153.200 1436.480 3153.460 ;
        RECT 1435.300 3056.640 1435.560 3056.900 ;
        RECT 1436.220 3056.640 1436.480 3056.900 ;
        RECT 1435.760 3042.700 1436.020 3042.960 ;
        RECT 1436.220 2994.760 1436.480 2995.020 ;
        RECT 1435.300 2863.520 1435.560 2863.780 ;
        RECT 1436.220 2863.520 1436.480 2863.780 ;
        RECT 1435.300 2753.020 1435.560 2753.280 ;
        RECT 1435.760 2753.020 1436.020 2753.280 ;
        RECT 1435.300 2704.400 1435.560 2704.660 ;
        RECT 1436.220 2704.400 1436.480 2704.660 ;
        RECT 1436.680 2670.400 1436.940 2670.660 ;
        RECT 1435.760 2656.460 1436.020 2656.720 ;
      LAYER met2 ;
        RECT 445.690 3518.000 446.250 3524.000 ;
        RECT 445.900 3504.030 446.040 3518.000 ;
        RECT 445.840 3503.710 446.100 3504.030 ;
        RECT 1436.220 3503.710 1436.480 3504.030 ;
        RECT 1436.280 3477.510 1436.420 3503.710 ;
        RECT 1436.220 3477.190 1436.480 3477.510 ;
        RECT 1435.760 3441.490 1436.020 3441.810 ;
        RECT 1435.820 3394.970 1435.960 3441.490 ;
        RECT 1435.820 3394.830 1436.420 3394.970 ;
        RECT 1436.280 3380.950 1436.420 3394.830 ;
        RECT 1436.220 3380.630 1436.480 3380.950 ;
        RECT 1435.760 3332.690 1436.020 3333.010 ;
        RECT 1435.820 3298.410 1435.960 3332.690 ;
        RECT 1435.820 3298.270 1436.420 3298.410 ;
        RECT 1436.280 3249.710 1436.420 3298.270 ;
        RECT 1436.220 3249.390 1436.480 3249.710 ;
        RECT 1436.220 3248.710 1436.480 3249.030 ;
        RECT 1436.280 3153.490 1436.420 3248.710 ;
        RECT 1435.300 3153.170 1435.560 3153.490 ;
        RECT 1436.220 3153.170 1436.480 3153.490 ;
        RECT 1435.360 3152.890 1435.500 3153.170 ;
        RECT 1435.360 3152.750 1435.960 3152.890 ;
        RECT 1435.820 3105.290 1435.960 3152.750 ;
        RECT 1435.820 3105.150 1436.420 3105.290 ;
        RECT 1436.280 3056.930 1436.420 3105.150 ;
        RECT 1435.300 3056.610 1435.560 3056.930 ;
        RECT 1436.220 3056.610 1436.480 3056.930 ;
        RECT 1435.360 3056.330 1435.500 3056.610 ;
        RECT 1435.360 3056.190 1435.960 3056.330 ;
        RECT 1435.820 3042.990 1435.960 3056.190 ;
        RECT 1435.760 3042.670 1436.020 3042.990 ;
        RECT 1436.220 2994.730 1436.480 2995.050 ;
        RECT 1436.280 2863.810 1436.420 2994.730 ;
        RECT 1435.300 2863.490 1435.560 2863.810 ;
        RECT 1436.220 2863.490 1436.480 2863.810 ;
        RECT 1435.360 2863.210 1435.500 2863.490 ;
        RECT 1435.360 2863.070 1435.960 2863.210 ;
        RECT 1435.820 2815.610 1435.960 2863.070 ;
        RECT 1435.820 2815.470 1436.420 2815.610 ;
        RECT 1436.280 2801.330 1436.420 2815.470 ;
        RECT 1435.820 2801.190 1436.420 2801.330 ;
        RECT 1435.820 2753.310 1435.960 2801.190 ;
        RECT 1435.300 2753.165 1435.560 2753.310 ;
        RECT 1435.290 2752.795 1435.570 2753.165 ;
        RECT 1435.760 2752.990 1436.020 2753.310 ;
        RECT 1436.210 2752.795 1436.490 2753.165 ;
        RECT 1436.280 2746.365 1436.420 2752.795 ;
        RECT 1435.290 2745.995 1435.570 2746.365 ;
        RECT 1436.210 2745.995 1436.490 2746.365 ;
        RECT 1435.360 2704.690 1435.500 2745.995 ;
        RECT 1435.300 2704.370 1435.560 2704.690 ;
        RECT 1436.220 2704.370 1436.480 2704.690 ;
        RECT 1436.280 2697.970 1436.420 2704.370 ;
        RECT 1436.280 2697.830 1436.880 2697.970 ;
        RECT 1436.740 2670.690 1436.880 2697.830 ;
        RECT 1436.680 2670.370 1436.940 2670.690 ;
        RECT 1435.760 2656.430 1436.020 2656.750 ;
        RECT 1435.820 2622.490 1435.960 2656.430 ;
        RECT 1435.360 2622.350 1435.960 2622.490 ;
        RECT 1435.360 2621.810 1435.500 2622.350 ;
        RECT 1435.360 2621.670 1435.960 2621.810 ;
        RECT 1435.210 2599.370 1435.490 2600.000 ;
        RECT 1435.820 2599.370 1435.960 2621.670 ;
        RECT 1435.210 2599.230 1435.960 2599.370 ;
        RECT 1435.210 2596.000 1435.490 2599.230 ;
      LAYER via2 ;
        RECT 1435.290 2752.840 1435.570 2753.120 ;
        RECT 1436.210 2752.840 1436.490 2753.120 ;
        RECT 1435.290 2746.040 1435.570 2746.320 ;
        RECT 1436.210 2746.040 1436.490 2746.320 ;
      LAYER met3 ;
        RECT 1435.265 2753.130 1435.595 2753.145 ;
        RECT 1436.185 2753.130 1436.515 2753.145 ;
        RECT 1435.265 2752.830 1436.515 2753.130 ;
        RECT 1435.265 2752.815 1435.595 2752.830 ;
        RECT 1436.185 2752.815 1436.515 2752.830 ;
        RECT 1435.265 2746.330 1435.595 2746.345 ;
        RECT 1436.185 2746.330 1436.515 2746.345 ;
        RECT 1435.265 2746.030 1436.515 2746.330 ;
        RECT 1435.265 2746.015 1435.595 2746.030 ;
        RECT 1436.185 2746.015 1436.515 2746.030 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1456.965 3490.865 1457.135 3502.255 ;
        RECT 1456.965 3442.925 1457.135 3477.435 ;
        RECT 1456.505 3139.645 1456.675 3187.755 ;
        RECT 1456.505 3043.085 1456.675 3091.195 ;
        RECT 1456.505 2987.665 1456.675 3035.775 ;
        RECT 1456.965 2849.625 1457.135 2898.075 ;
      LAYER mcon ;
        RECT 1456.965 3502.085 1457.135 3502.255 ;
        RECT 1456.965 3477.265 1457.135 3477.435 ;
        RECT 1456.505 3187.585 1456.675 3187.755 ;
        RECT 1456.505 3091.025 1456.675 3091.195 ;
        RECT 1456.505 3035.605 1456.675 3035.775 ;
        RECT 1456.965 2897.905 1457.135 2898.075 ;
      LAYER met1 ;
        RECT 121.510 3502.240 121.830 3502.300 ;
        RECT 1456.905 3502.240 1457.195 3502.285 ;
        RECT 121.510 3502.100 1457.195 3502.240 ;
        RECT 121.510 3502.040 121.830 3502.100 ;
        RECT 1456.905 3502.055 1457.195 3502.100 ;
        RECT 1456.890 3491.020 1457.210 3491.080 ;
        RECT 1456.695 3490.880 1457.210 3491.020 ;
        RECT 1456.890 3490.820 1457.210 3490.880 ;
        RECT 1456.890 3477.420 1457.210 3477.480 ;
        RECT 1456.695 3477.280 1457.210 3477.420 ;
        RECT 1456.890 3477.220 1457.210 3477.280 ;
        RECT 1456.890 3443.080 1457.210 3443.140 ;
        RECT 1456.695 3442.940 1457.210 3443.080 ;
        RECT 1456.890 3442.880 1457.210 3442.940 ;
        RECT 1457.350 3395.140 1457.670 3395.200 ;
        RECT 1456.980 3395.000 1457.670 3395.140 ;
        RECT 1456.980 3394.860 1457.120 3395.000 ;
        RECT 1457.350 3394.940 1457.670 3395.000 ;
        RECT 1456.890 3394.600 1457.210 3394.860 ;
        RECT 1456.445 3187.740 1456.735 3187.785 ;
        RECT 1456.890 3187.740 1457.210 3187.800 ;
        RECT 1456.445 3187.600 1457.210 3187.740 ;
        RECT 1456.445 3187.555 1456.735 3187.600 ;
        RECT 1456.890 3187.540 1457.210 3187.600 ;
        RECT 1456.430 3139.800 1456.750 3139.860 ;
        RECT 1456.235 3139.660 1456.750 3139.800 ;
        RECT 1456.430 3139.600 1456.750 3139.660 ;
        RECT 1456.445 3091.180 1456.735 3091.225 ;
        RECT 1456.890 3091.180 1457.210 3091.240 ;
        RECT 1456.445 3091.040 1457.210 3091.180 ;
        RECT 1456.445 3090.995 1456.735 3091.040 ;
        RECT 1456.890 3090.980 1457.210 3091.040 ;
        RECT 1456.430 3043.240 1456.750 3043.300 ;
        RECT 1456.235 3043.100 1456.750 3043.240 ;
        RECT 1456.430 3043.040 1456.750 3043.100 ;
        RECT 1456.430 3035.760 1456.750 3035.820 ;
        RECT 1456.235 3035.620 1456.750 3035.760 ;
        RECT 1456.430 3035.560 1456.750 3035.620 ;
        RECT 1456.445 2987.820 1456.735 2987.865 ;
        RECT 1456.890 2987.820 1457.210 2987.880 ;
        RECT 1456.445 2987.680 1457.210 2987.820 ;
        RECT 1456.445 2987.635 1456.735 2987.680 ;
        RECT 1456.890 2987.620 1457.210 2987.680 ;
        RECT 1456.890 2898.060 1457.210 2898.120 ;
        RECT 1456.695 2897.920 1457.210 2898.060 ;
        RECT 1456.890 2897.860 1457.210 2897.920 ;
        RECT 1456.905 2849.780 1457.195 2849.825 ;
        RECT 1457.350 2849.780 1457.670 2849.840 ;
        RECT 1456.905 2849.640 1457.670 2849.780 ;
        RECT 1456.905 2849.595 1457.195 2849.640 ;
        RECT 1457.350 2849.580 1457.670 2849.640 ;
        RECT 1457.350 2815.780 1457.670 2815.840 ;
        RECT 1456.980 2815.640 1457.670 2815.780 ;
        RECT 1456.980 2815.160 1457.120 2815.640 ;
        RECT 1457.350 2815.580 1457.670 2815.640 ;
        RECT 1456.890 2814.900 1457.210 2815.160 ;
        RECT 1456.430 2766.620 1456.750 2766.880 ;
        RECT 1456.520 2766.200 1456.660 2766.620 ;
        RECT 1456.430 2765.940 1456.750 2766.200 ;
        RECT 1456.430 2656.660 1456.750 2656.720 ;
        RECT 1459.190 2656.660 1459.510 2656.720 ;
        RECT 1456.430 2656.520 1459.510 2656.660 ;
        RECT 1456.430 2656.460 1456.750 2656.520 ;
        RECT 1459.190 2656.460 1459.510 2656.520 ;
      LAYER via ;
        RECT 121.540 3502.040 121.800 3502.300 ;
        RECT 1456.920 3490.820 1457.180 3491.080 ;
        RECT 1456.920 3477.220 1457.180 3477.480 ;
        RECT 1456.920 3442.880 1457.180 3443.140 ;
        RECT 1457.380 3394.940 1457.640 3395.200 ;
        RECT 1456.920 3394.600 1457.180 3394.860 ;
        RECT 1456.920 3187.540 1457.180 3187.800 ;
        RECT 1456.460 3139.600 1456.720 3139.860 ;
        RECT 1456.920 3090.980 1457.180 3091.240 ;
        RECT 1456.460 3043.040 1456.720 3043.300 ;
        RECT 1456.460 3035.560 1456.720 3035.820 ;
        RECT 1456.920 2987.620 1457.180 2987.880 ;
        RECT 1456.920 2897.860 1457.180 2898.120 ;
        RECT 1457.380 2849.580 1457.640 2849.840 ;
        RECT 1457.380 2815.580 1457.640 2815.840 ;
        RECT 1456.920 2814.900 1457.180 2815.160 ;
        RECT 1456.460 2766.620 1456.720 2766.880 ;
        RECT 1456.460 2765.940 1456.720 2766.200 ;
        RECT 1456.460 2656.460 1456.720 2656.720 ;
        RECT 1459.220 2656.460 1459.480 2656.720 ;
      LAYER met2 ;
        RECT 121.390 3518.000 121.950 3524.000 ;
        RECT 121.600 3502.330 121.740 3518.000 ;
        RECT 121.540 3502.010 121.800 3502.330 ;
        RECT 1456.920 3490.790 1457.180 3491.110 ;
        RECT 1456.980 3477.510 1457.120 3490.790 ;
        RECT 1456.920 3477.190 1457.180 3477.510 ;
        RECT 1456.920 3442.850 1457.180 3443.170 ;
        RECT 1456.980 3429.650 1457.120 3442.850 ;
        RECT 1456.980 3429.510 1457.580 3429.650 ;
        RECT 1457.440 3395.230 1457.580 3429.510 ;
        RECT 1457.380 3394.910 1457.640 3395.230 ;
        RECT 1456.920 3394.570 1457.180 3394.890 ;
        RECT 1456.980 3187.830 1457.120 3394.570 ;
        RECT 1456.920 3187.510 1457.180 3187.830 ;
        RECT 1456.460 3139.570 1456.720 3139.890 ;
        RECT 1456.520 3139.290 1456.660 3139.570 ;
        RECT 1456.520 3139.150 1457.120 3139.290 ;
        RECT 1456.980 3091.270 1457.120 3139.150 ;
        RECT 1456.920 3090.950 1457.180 3091.270 ;
        RECT 1456.460 3043.010 1456.720 3043.330 ;
        RECT 1456.520 3035.850 1456.660 3043.010 ;
        RECT 1456.460 3035.530 1456.720 3035.850 ;
        RECT 1456.920 2987.590 1457.180 2987.910 ;
        RECT 1456.980 2898.150 1457.120 2987.590 ;
        RECT 1456.920 2897.830 1457.180 2898.150 ;
        RECT 1457.380 2849.550 1457.640 2849.870 ;
        RECT 1457.440 2815.870 1457.580 2849.550 ;
        RECT 1457.380 2815.550 1457.640 2815.870 ;
        RECT 1456.920 2814.870 1457.180 2815.190 ;
        RECT 1456.980 2801.330 1457.120 2814.870 ;
        RECT 1456.520 2801.190 1457.120 2801.330 ;
        RECT 1456.520 2766.910 1456.660 2801.190 ;
        RECT 1456.460 2766.590 1456.720 2766.910 ;
        RECT 1456.460 2765.910 1456.720 2766.230 ;
        RECT 1456.520 2746.365 1456.660 2765.910 ;
        RECT 1455.530 2745.995 1455.810 2746.365 ;
        RECT 1456.450 2745.995 1456.730 2746.365 ;
        RECT 1455.600 2703.410 1455.740 2745.995 ;
        RECT 1455.600 2703.270 1456.660 2703.410 ;
        RECT 1456.520 2656.750 1456.660 2703.270 ;
        RECT 1456.460 2656.430 1456.720 2656.750 ;
        RECT 1459.220 2656.430 1459.480 2656.750 ;
        RECT 1459.280 2632.010 1459.420 2656.430 ;
        RECT 1458.360 2631.870 1459.420 2632.010 ;
        RECT 1458.360 2600.050 1458.500 2631.870 ;
        RECT 1458.360 2600.000 1461.190 2600.050 ;
        RECT 1458.360 2599.910 1461.250 2600.000 ;
        RECT 1460.970 2596.000 1461.250 2599.910 ;
      LAYER via2 ;
        RECT 1455.530 2746.040 1455.810 2746.320 ;
        RECT 1456.450 2746.040 1456.730 2746.320 ;
      LAYER met3 ;
        RECT 1455.505 2746.330 1455.835 2746.345 ;
        RECT 1456.425 2746.330 1456.755 2746.345 ;
        RECT 1455.505 2746.030 1456.755 2746.330 ;
        RECT 1455.505 2746.015 1455.835 2746.030 ;
        RECT 1456.425 2746.015 1456.755 2746.030 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 3339.720 17.410 3339.780 ;
        RECT 1483.570 3339.720 1483.890 3339.780 ;
        RECT 17.090 3339.580 1483.890 3339.720 ;
        RECT 17.090 3339.520 17.410 3339.580 ;
        RECT 1483.570 3339.520 1483.890 3339.580 ;
      LAYER via ;
        RECT 17.120 3339.520 17.380 3339.780 ;
        RECT 1483.600 3339.520 1483.860 3339.780 ;
      LAYER met2 ;
        RECT 17.110 3339.635 17.390 3340.005 ;
        RECT 17.120 3339.490 17.380 3339.635 ;
        RECT 1483.600 3339.490 1483.860 3339.810 ;
        RECT 1483.660 2601.410 1483.800 3339.490 ;
        RECT 1483.660 2601.270 1484.720 2601.410 ;
        RECT 1484.580 2600.050 1484.720 2601.270 ;
        RECT 1484.580 2600.000 1486.950 2600.050 ;
        RECT 1484.580 2599.910 1487.010 2600.000 ;
        RECT 1486.730 2596.000 1487.010 2599.910 ;
      LAYER via2 ;
        RECT 17.110 3339.680 17.390 3339.960 ;
      LAYER met3 ;
        RECT -4.000 3339.970 2.000 3340.420 ;
        RECT 17.085 3339.970 17.415 3339.985 ;
        RECT -4.000 3339.670 17.415 3339.970 ;
        RECT -4.000 3339.220 2.000 3339.670 ;
        RECT 17.085 3339.655 17.415 3339.670 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 3050.040 17.410 3050.100 ;
        RECT 1511.170 3050.040 1511.490 3050.100 ;
        RECT 17.090 3049.900 1511.490 3050.040 ;
        RECT 17.090 3049.840 17.410 3049.900 ;
        RECT 1511.170 3049.840 1511.490 3049.900 ;
      LAYER via ;
        RECT 17.120 3049.840 17.380 3050.100 ;
        RECT 1511.200 3049.840 1511.460 3050.100 ;
      LAYER met2 ;
        RECT 17.110 3051.995 17.390 3052.365 ;
        RECT 17.180 3050.130 17.320 3051.995 ;
        RECT 17.120 3049.810 17.380 3050.130 ;
        RECT 1511.200 3049.810 1511.460 3050.130 ;
        RECT 1511.260 2600.050 1511.400 3049.810 ;
        RECT 1511.260 2600.000 1512.250 2600.050 ;
        RECT 1511.260 2599.910 1512.310 2600.000 ;
        RECT 1512.030 2596.000 1512.310 2599.910 ;
      LAYER via2 ;
        RECT 17.110 3052.040 17.390 3052.320 ;
      LAYER met3 ;
        RECT -4.000 3052.330 2.000 3052.780 ;
        RECT 17.085 3052.330 17.415 3052.345 ;
        RECT -4.000 3052.030 17.415 3052.330 ;
        RECT -4.000 3051.580 2.000 3052.030 ;
        RECT 17.085 3052.015 17.415 3052.030 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 2760.360 16.030 2760.420 ;
        RECT 1531.870 2760.360 1532.190 2760.420 ;
        RECT 15.710 2760.220 1532.190 2760.360 ;
        RECT 15.710 2760.160 16.030 2760.220 ;
        RECT 1531.870 2760.160 1532.190 2760.220 ;
      LAYER via ;
        RECT 15.740 2760.160 16.000 2760.420 ;
        RECT 1531.900 2760.160 1532.160 2760.420 ;
      LAYER met2 ;
        RECT 15.730 2765.035 16.010 2765.405 ;
        RECT 15.800 2760.450 15.940 2765.035 ;
        RECT 15.740 2760.130 16.000 2760.450 ;
        RECT 1531.900 2760.130 1532.160 2760.450 ;
        RECT 1531.960 2600.730 1532.100 2760.130 ;
        RECT 1531.960 2600.590 1535.320 2600.730 ;
        RECT 1535.180 2600.050 1535.320 2600.590 ;
        RECT 1535.180 2600.000 1538.010 2600.050 ;
        RECT 1535.180 2599.910 1538.070 2600.000 ;
        RECT 1537.790 2596.000 1538.070 2599.910 ;
      LAYER via2 ;
        RECT 15.730 2765.080 16.010 2765.360 ;
      LAYER met3 ;
        RECT -4.000 2765.370 2.000 2765.820 ;
        RECT 15.705 2765.370 16.035 2765.385 ;
        RECT -4.000 2765.070 16.035 2765.370 ;
        RECT -4.000 2764.620 2.000 2765.070 ;
        RECT 15.705 2765.055 16.035 2765.070 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 23.530 2613.480 23.850 2613.540 ;
        RECT 1562.230 2613.480 1562.550 2613.540 ;
        RECT 23.530 2613.340 1562.550 2613.480 ;
        RECT 23.530 2613.280 23.850 2613.340 ;
        RECT 1562.230 2613.280 1562.550 2613.340 ;
        RECT 13.870 2477.820 14.190 2477.880 ;
        RECT 23.530 2477.820 23.850 2477.880 ;
        RECT 13.870 2477.680 23.850 2477.820 ;
        RECT 13.870 2477.620 14.190 2477.680 ;
        RECT 23.530 2477.620 23.850 2477.680 ;
      LAYER via ;
        RECT 23.560 2613.280 23.820 2613.540 ;
        RECT 1562.260 2613.280 1562.520 2613.540 ;
        RECT 13.900 2477.620 14.160 2477.880 ;
        RECT 23.560 2477.620 23.820 2477.880 ;
      LAYER met2 ;
        RECT 23.560 2613.250 23.820 2613.570 ;
        RECT 1562.260 2613.250 1562.520 2613.570 ;
        RECT 23.620 2477.910 23.760 2613.250 ;
        RECT 1562.320 2600.050 1562.460 2613.250 ;
        RECT 1562.320 2600.000 1563.770 2600.050 ;
        RECT 1562.320 2599.910 1563.830 2600.000 ;
        RECT 1563.550 2596.000 1563.830 2599.910 ;
        RECT 13.900 2477.765 14.160 2477.910 ;
        RECT 13.890 2477.395 14.170 2477.765 ;
        RECT 23.560 2477.590 23.820 2477.910 ;
      LAYER via2 ;
        RECT 13.890 2477.440 14.170 2477.720 ;
      LAYER met3 ;
        RECT -4.000 2477.730 2.000 2478.180 ;
        RECT 13.865 2477.730 14.195 2477.745 ;
        RECT -4.000 2477.430 14.195 2477.730 ;
        RECT -4.000 2476.980 2.000 2477.430 ;
        RECT 13.865 2477.415 14.195 2477.430 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 2612.800 16.030 2612.860 ;
        RECT 1587.070 2612.800 1587.390 2612.860 ;
        RECT 15.710 2612.660 1587.390 2612.800 ;
        RECT 15.710 2612.600 16.030 2612.660 ;
        RECT 1587.070 2612.600 1587.390 2612.660 ;
      LAYER via ;
        RECT 15.740 2612.600 16.000 2612.860 ;
        RECT 1587.100 2612.600 1587.360 2612.860 ;
      LAYER met2 ;
        RECT 15.740 2612.570 16.000 2612.890 ;
        RECT 1587.100 2612.570 1587.360 2612.890 ;
        RECT 15.800 2190.125 15.940 2612.570 ;
        RECT 1587.160 2600.050 1587.300 2612.570 ;
        RECT 1587.160 2600.000 1589.070 2600.050 ;
        RECT 1587.160 2599.910 1589.130 2600.000 ;
        RECT 1588.850 2596.000 1589.130 2599.910 ;
        RECT 15.730 2189.755 16.010 2190.125 ;
      LAYER via2 ;
        RECT 15.730 2189.800 16.010 2190.080 ;
      LAYER met3 ;
        RECT -4.000 2190.090 2.000 2190.540 ;
        RECT 15.705 2190.090 16.035 2190.105 ;
        RECT -4.000 2189.790 16.035 2190.090 ;
        RECT -4.000 2189.340 2.000 2189.790 ;
        RECT 15.705 2189.775 16.035 2189.790 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 27.210 2612.120 27.530 2612.180 ;
        RECT 1615.130 2612.120 1615.450 2612.180 ;
        RECT 27.210 2611.980 1615.450 2612.120 ;
        RECT 27.210 2611.920 27.530 2611.980 ;
        RECT 1615.130 2611.920 1615.450 2611.980 ;
        RECT 13.870 1903.220 14.190 1903.280 ;
        RECT 27.210 1903.220 27.530 1903.280 ;
        RECT 13.870 1903.080 27.530 1903.220 ;
        RECT 13.870 1903.020 14.190 1903.080 ;
        RECT 27.210 1903.020 27.530 1903.080 ;
      LAYER via ;
        RECT 27.240 2611.920 27.500 2612.180 ;
        RECT 1615.160 2611.920 1615.420 2612.180 ;
        RECT 13.900 1903.020 14.160 1903.280 ;
        RECT 27.240 1903.020 27.500 1903.280 ;
      LAYER met2 ;
        RECT 27.240 2611.890 27.500 2612.210 ;
        RECT 1615.160 2611.890 1615.420 2612.210 ;
        RECT 27.300 1903.310 27.440 2611.890 ;
        RECT 1614.610 2599.370 1614.890 2600.000 ;
        RECT 1615.220 2599.370 1615.360 2611.890 ;
        RECT 1614.610 2599.230 1615.360 2599.370 ;
        RECT 1614.610 2596.000 1614.890 2599.230 ;
        RECT 13.900 1903.165 14.160 1903.310 ;
        RECT 13.890 1902.795 14.170 1903.165 ;
        RECT 27.240 1902.990 27.500 1903.310 ;
      LAYER via2 ;
        RECT 13.890 1902.840 14.170 1903.120 ;
      LAYER met3 ;
        RECT -4.000 1903.130 2.000 1903.580 ;
        RECT 13.865 1903.130 14.195 1903.145 ;
        RECT -4.000 1902.830 14.195 1903.130 ;
        RECT -4.000 1902.380 2.000 1902.830 ;
        RECT 13.865 1902.815 14.195 1902.830 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1628.470 2612.120 1628.790 2612.180 ;
        RECT 1676.310 2612.120 1676.630 2612.180 ;
        RECT 1628.470 2611.980 1676.630 2612.120 ;
        RECT 1628.470 2611.920 1628.790 2611.980 ;
        RECT 1676.310 2611.920 1676.630 2611.980 ;
        RECT 1725.070 2611.100 1725.390 2611.160 ;
        RECT 1772.910 2611.100 1773.230 2611.160 ;
        RECT 1725.070 2610.960 1773.230 2611.100 ;
        RECT 1725.070 2610.900 1725.390 2610.960 ;
        RECT 1772.910 2610.900 1773.230 2610.960 ;
        RECT 1559.010 2608.040 1559.330 2608.100 ;
        RECT 1559.930 2608.040 1560.250 2608.100 ;
        RECT 1559.010 2607.900 1560.250 2608.040 ;
        RECT 1559.010 2607.840 1559.330 2607.900 ;
        RECT 1559.930 2607.840 1560.250 2607.900 ;
      LAYER via ;
        RECT 1628.500 2611.920 1628.760 2612.180 ;
        RECT 1676.340 2611.920 1676.600 2612.180 ;
        RECT 1725.100 2610.900 1725.360 2611.160 ;
        RECT 1772.940 2610.900 1773.200 2611.160 ;
        RECT 1559.040 2607.840 1559.300 2608.100 ;
        RECT 1559.960 2607.840 1560.220 2608.100 ;
      LAYER met2 ;
        RECT 924.230 2613.395 924.510 2613.765 ;
        RECT 953.210 2613.395 953.490 2613.765 ;
        RECT 922.310 2599.370 922.590 2600.000 ;
        RECT 924.300 2599.370 924.440 2613.395 ;
        RECT 953.280 2611.045 953.420 2613.395 ;
        RECT 1628.500 2611.890 1628.760 2612.210 ;
        RECT 1676.340 2611.890 1676.600 2612.210 ;
        RECT 1628.560 2611.045 1628.700 2611.890 ;
        RECT 1676.400 2611.045 1676.540 2611.890 ;
        RECT 1725.100 2611.045 1725.360 2611.190 ;
        RECT 1772.940 2611.045 1773.200 2611.190 ;
        RECT 953.210 2610.675 953.490 2611.045 ;
        RECT 1559.030 2610.675 1559.310 2611.045 ;
        RECT 1559.950 2610.675 1560.230 2611.045 ;
        RECT 1628.490 2610.675 1628.770 2611.045 ;
        RECT 1676.330 2610.675 1676.610 2611.045 ;
        RECT 1725.090 2610.675 1725.370 2611.045 ;
        RECT 1772.930 2610.675 1773.210 2611.045 ;
        RECT 2904.070 2610.675 2904.350 2611.045 ;
        RECT 1559.100 2608.130 1559.240 2610.675 ;
        RECT 1560.020 2608.130 1560.160 2610.675 ;
        RECT 1559.040 2607.810 1559.300 2608.130 ;
        RECT 1559.960 2607.810 1560.220 2608.130 ;
        RECT 922.310 2599.230 924.440 2599.370 ;
        RECT 922.310 2596.000 922.590 2599.230 ;
        RECT 2904.140 615.925 2904.280 2610.675 ;
        RECT 2904.070 615.555 2904.350 615.925 ;
      LAYER via2 ;
        RECT 924.230 2613.440 924.510 2613.720 ;
        RECT 953.210 2613.440 953.490 2613.720 ;
        RECT 953.210 2610.720 953.490 2611.000 ;
        RECT 1559.030 2610.720 1559.310 2611.000 ;
        RECT 1559.950 2610.720 1560.230 2611.000 ;
        RECT 1628.490 2610.720 1628.770 2611.000 ;
        RECT 1676.330 2610.720 1676.610 2611.000 ;
        RECT 1725.090 2610.720 1725.370 2611.000 ;
        RECT 1772.930 2610.720 1773.210 2611.000 ;
        RECT 2904.070 2610.720 2904.350 2611.000 ;
        RECT 2904.070 615.600 2904.350 615.880 ;
      LAYER met3 ;
        RECT 924.205 2613.730 924.535 2613.745 ;
        RECT 953.185 2613.730 953.515 2613.745 ;
        RECT 924.205 2613.430 953.515 2613.730 ;
        RECT 924.205 2613.415 924.535 2613.430 ;
        RECT 953.185 2613.415 953.515 2613.430 ;
        RECT 953.185 2611.010 953.515 2611.025 ;
        RECT 1559.005 2611.010 1559.335 2611.025 ;
        RECT 953.185 2610.710 1559.335 2611.010 ;
        RECT 953.185 2610.695 953.515 2610.710 ;
        RECT 1559.005 2610.695 1559.335 2610.710 ;
        RECT 1559.925 2611.010 1560.255 2611.025 ;
        RECT 1628.465 2611.010 1628.795 2611.025 ;
        RECT 1559.925 2610.710 1628.795 2611.010 ;
        RECT 1559.925 2610.695 1560.255 2610.710 ;
        RECT 1628.465 2610.695 1628.795 2610.710 ;
        RECT 1676.305 2611.010 1676.635 2611.025 ;
        RECT 1725.065 2611.010 1725.395 2611.025 ;
        RECT 1676.305 2610.710 1725.395 2611.010 ;
        RECT 1676.305 2610.695 1676.635 2610.710 ;
        RECT 1725.065 2610.695 1725.395 2610.710 ;
        RECT 1772.905 2611.010 1773.235 2611.025 ;
        RECT 2904.045 2611.010 2904.375 2611.025 ;
        RECT 1772.905 2610.710 2904.375 2611.010 ;
        RECT 1772.905 2610.695 1773.235 2610.710 ;
        RECT 2904.045 2610.695 2904.375 2610.710 ;
        RECT 2904.045 615.890 2904.375 615.905 ;
        RECT 2918.000 615.890 2924.000 616.340 ;
        RECT 2904.045 615.590 2924.000 615.890 ;
        RECT 2904.045 615.575 2904.375 615.590 ;
        RECT 2918.000 615.140 2924.000 615.590 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 30.890 2611.780 31.210 2611.840 ;
        RECT 1638.590 2611.780 1638.910 2611.840 ;
        RECT 30.890 2611.640 1638.910 2611.780 ;
        RECT 30.890 2611.580 31.210 2611.640 ;
        RECT 1638.590 2611.580 1638.910 2611.640 ;
        RECT 15.710 1621.020 16.030 1621.080 ;
        RECT 30.890 1621.020 31.210 1621.080 ;
        RECT 15.710 1620.880 31.210 1621.020 ;
        RECT 15.710 1620.820 16.030 1620.880 ;
        RECT 30.890 1620.820 31.210 1620.880 ;
      LAYER via ;
        RECT 30.920 2611.580 31.180 2611.840 ;
        RECT 1638.620 2611.580 1638.880 2611.840 ;
        RECT 15.740 1620.820 16.000 1621.080 ;
        RECT 30.920 1620.820 31.180 1621.080 ;
      LAYER met2 ;
        RECT 30.920 2611.550 31.180 2611.870 ;
        RECT 1638.620 2611.550 1638.880 2611.870 ;
        RECT 30.980 1621.110 31.120 2611.550 ;
        RECT 1638.680 2600.050 1638.820 2611.550 ;
        RECT 1638.680 2600.000 1640.590 2600.050 ;
        RECT 1638.680 2599.910 1640.650 2600.000 ;
        RECT 1640.370 2596.000 1640.650 2599.910 ;
        RECT 15.740 1620.790 16.000 1621.110 ;
        RECT 30.920 1620.790 31.180 1621.110 ;
        RECT 15.800 1615.525 15.940 1620.790 ;
        RECT 15.730 1615.155 16.010 1615.525 ;
      LAYER via2 ;
        RECT 15.730 1615.200 16.010 1615.480 ;
      LAYER met3 ;
        RECT -4.000 1615.490 2.000 1615.940 ;
        RECT 15.705 1615.490 16.035 1615.505 ;
        RECT -4.000 1615.190 16.035 1615.490 ;
        RECT -4.000 1614.740 2.000 1615.190 ;
        RECT 15.705 1615.175 16.035 1615.190 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 51.590 2610.760 51.910 2610.820 ;
        RECT 1664.350 2610.760 1664.670 2610.820 ;
        RECT 51.590 2610.620 1664.670 2610.760 ;
        RECT 51.590 2610.560 51.910 2610.620 ;
        RECT 1664.350 2610.560 1664.670 2610.620 ;
        RECT 16.630 1400.700 16.950 1400.760 ;
        RECT 51.590 1400.700 51.910 1400.760 ;
        RECT 16.630 1400.560 51.910 1400.700 ;
        RECT 16.630 1400.500 16.950 1400.560 ;
        RECT 51.590 1400.500 51.910 1400.560 ;
      LAYER via ;
        RECT 51.620 2610.560 51.880 2610.820 ;
        RECT 1664.380 2610.560 1664.640 2610.820 ;
        RECT 16.660 1400.500 16.920 1400.760 ;
        RECT 51.620 1400.500 51.880 1400.760 ;
      LAYER met2 ;
        RECT 51.620 2610.530 51.880 2610.850 ;
        RECT 1664.380 2610.530 1664.640 2610.850 ;
        RECT 51.680 1400.790 51.820 2610.530 ;
        RECT 1664.440 2600.050 1664.580 2610.530 ;
        RECT 1664.440 2600.000 1666.350 2600.050 ;
        RECT 1664.440 2599.910 1666.410 2600.000 ;
        RECT 1666.130 2596.000 1666.410 2599.910 ;
        RECT 16.660 1400.645 16.920 1400.790 ;
        RECT 16.650 1400.275 16.930 1400.645 ;
        RECT 51.620 1400.470 51.880 1400.790 ;
      LAYER via2 ;
        RECT 16.650 1400.320 16.930 1400.600 ;
      LAYER met3 ;
        RECT -4.000 1400.610 2.000 1401.060 ;
        RECT 16.625 1400.610 16.955 1400.625 ;
        RECT -4.000 1400.310 16.955 1400.610 ;
        RECT -4.000 1399.860 2.000 1400.310 ;
        RECT 16.625 1400.295 16.955 1400.310 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 65.390 2610.420 65.710 2610.480 ;
        RECT 1690.570 2610.420 1690.890 2610.480 ;
        RECT 65.390 2610.280 1690.890 2610.420 ;
        RECT 65.390 2610.220 65.710 2610.280 ;
        RECT 1690.570 2610.220 1690.890 2610.280 ;
        RECT 16.630 1186.840 16.950 1186.900 ;
        RECT 65.390 1186.840 65.710 1186.900 ;
        RECT 16.630 1186.700 65.710 1186.840 ;
        RECT 16.630 1186.640 16.950 1186.700 ;
        RECT 65.390 1186.640 65.710 1186.700 ;
      LAYER via ;
        RECT 65.420 2610.220 65.680 2610.480 ;
        RECT 1690.600 2610.220 1690.860 2610.480 ;
        RECT 16.660 1186.640 16.920 1186.900 ;
        RECT 65.420 1186.640 65.680 1186.900 ;
      LAYER met2 ;
        RECT 65.420 2610.190 65.680 2610.510 ;
        RECT 1690.600 2610.190 1690.860 2610.510 ;
        RECT 65.480 1186.930 65.620 2610.190 ;
        RECT 1690.660 2600.050 1690.800 2610.190 ;
        RECT 1690.660 2600.000 1691.650 2600.050 ;
        RECT 1690.660 2599.910 1691.710 2600.000 ;
        RECT 1691.430 2596.000 1691.710 2599.910 ;
        RECT 16.660 1186.610 16.920 1186.930 ;
        RECT 65.420 1186.610 65.680 1186.930 ;
        RECT 16.720 1185.085 16.860 1186.610 ;
        RECT 16.650 1184.715 16.930 1185.085 ;
      LAYER via2 ;
        RECT 16.650 1184.760 16.930 1185.040 ;
      LAYER met3 ;
        RECT -4.000 1185.050 2.000 1185.500 ;
        RECT 16.625 1185.050 16.955 1185.065 ;
        RECT -4.000 1184.750 16.955 1185.050 ;
        RECT -4.000 1184.300 2.000 1184.750 ;
        RECT 16.625 1184.735 16.955 1184.750 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 99.890 2611.100 100.210 2611.160 ;
        RECT 1715.870 2611.100 1716.190 2611.160 ;
        RECT 99.890 2610.960 1716.190 2611.100 ;
        RECT 99.890 2610.900 100.210 2610.960 ;
        RECT 1715.870 2610.900 1716.190 2610.960 ;
        RECT 15.710 972.640 16.030 972.700 ;
        RECT 99.890 972.640 100.210 972.700 ;
        RECT 15.710 972.500 100.210 972.640 ;
        RECT 15.710 972.440 16.030 972.500 ;
        RECT 99.890 972.440 100.210 972.500 ;
      LAYER via ;
        RECT 99.920 2610.900 100.180 2611.160 ;
        RECT 1715.900 2610.900 1716.160 2611.160 ;
        RECT 15.740 972.440 16.000 972.700 ;
        RECT 99.920 972.440 100.180 972.700 ;
      LAYER met2 ;
        RECT 99.920 2610.870 100.180 2611.190 ;
        RECT 1715.900 2610.870 1716.160 2611.190 ;
        RECT 99.980 972.730 100.120 2610.870 ;
        RECT 1715.960 2600.050 1716.100 2610.870 ;
        RECT 1715.960 2600.000 1717.410 2600.050 ;
        RECT 1715.960 2599.910 1717.470 2600.000 ;
        RECT 1717.190 2596.000 1717.470 2599.910 ;
        RECT 15.740 972.410 16.000 972.730 ;
        RECT 99.920 972.410 100.180 972.730 ;
        RECT 15.800 969.525 15.940 972.410 ;
        RECT 15.730 969.155 16.010 969.525 ;
      LAYER via2 ;
        RECT 15.730 969.200 16.010 969.480 ;
      LAYER met3 ;
        RECT -4.000 969.490 2.000 969.940 ;
        RECT 15.705 969.490 16.035 969.505 ;
        RECT -4.000 969.190 16.035 969.490 ;
        RECT -4.000 968.740 2.000 969.190 ;
        RECT 15.705 969.175 16.035 969.190 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 106.790 2609.740 107.110 2609.800 ;
        RECT 1741.630 2609.740 1741.950 2609.800 ;
        RECT 106.790 2609.600 1741.950 2609.740 ;
        RECT 106.790 2609.540 107.110 2609.600 ;
        RECT 1741.630 2609.540 1741.950 2609.600 ;
        RECT 16.630 758.780 16.950 758.840 ;
        RECT 106.790 758.780 107.110 758.840 ;
        RECT 16.630 758.640 107.110 758.780 ;
        RECT 16.630 758.580 16.950 758.640 ;
        RECT 106.790 758.580 107.110 758.640 ;
      LAYER via ;
        RECT 106.820 2609.540 107.080 2609.800 ;
        RECT 1741.660 2609.540 1741.920 2609.800 ;
        RECT 16.660 758.580 16.920 758.840 ;
        RECT 106.820 758.580 107.080 758.840 ;
      LAYER met2 ;
        RECT 106.820 2609.510 107.080 2609.830 ;
        RECT 1741.660 2609.510 1741.920 2609.830 ;
        RECT 106.880 758.870 107.020 2609.510 ;
        RECT 1741.720 2600.050 1741.860 2609.510 ;
        RECT 1741.720 2600.000 1743.170 2600.050 ;
        RECT 1741.720 2599.910 1743.230 2600.000 ;
        RECT 1742.950 2596.000 1743.230 2599.910 ;
        RECT 16.660 758.550 16.920 758.870 ;
        RECT 106.820 758.550 107.080 758.870 ;
        RECT 16.720 753.965 16.860 758.550 ;
        RECT 16.650 753.595 16.930 753.965 ;
      LAYER via2 ;
        RECT 16.650 753.640 16.930 753.920 ;
      LAYER met3 ;
        RECT -4.000 753.930 2.000 754.380 ;
        RECT 16.625 753.930 16.955 753.945 ;
        RECT -4.000 753.630 16.955 753.930 ;
        RECT -4.000 753.180 2.000 753.630 ;
        RECT 16.625 753.615 16.955 753.630 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 544.920 16.950 544.980 ;
        RECT 141.290 544.920 141.610 544.980 ;
        RECT 16.630 544.780 141.610 544.920 ;
        RECT 16.630 544.720 16.950 544.780 ;
        RECT 141.290 544.720 141.610 544.780 ;
      LAYER via ;
        RECT 16.660 544.720 16.920 544.980 ;
        RECT 141.320 544.720 141.580 544.980 ;
      LAYER met2 ;
        RECT 141.310 2612.035 141.590 2612.405 ;
        RECT 1767.410 2612.035 1767.690 2612.405 ;
        RECT 141.380 545.010 141.520 2612.035 ;
        RECT 1767.480 2600.050 1767.620 2612.035 ;
        RECT 1767.480 2600.000 1768.930 2600.050 ;
        RECT 1767.480 2599.910 1768.990 2600.000 ;
        RECT 1768.710 2596.000 1768.990 2599.910 ;
        RECT 16.660 544.690 16.920 545.010 ;
        RECT 141.320 544.690 141.580 545.010 ;
        RECT 16.720 538.405 16.860 544.690 ;
        RECT 16.650 538.035 16.930 538.405 ;
      LAYER via2 ;
        RECT 141.310 2612.080 141.590 2612.360 ;
        RECT 1767.410 2612.080 1767.690 2612.360 ;
        RECT 16.650 538.080 16.930 538.360 ;
      LAYER met3 ;
        RECT 141.285 2612.370 141.615 2612.385 ;
        RECT 1767.385 2612.370 1767.715 2612.385 ;
        RECT 141.285 2612.070 1767.715 2612.370 ;
        RECT 141.285 2612.055 141.615 2612.070 ;
        RECT 1767.385 2612.055 1767.715 2612.070 ;
        RECT -4.000 538.370 2.000 538.820 ;
        RECT 16.625 538.370 16.955 538.385 ;
        RECT -4.000 538.070 16.955 538.370 ;
        RECT -4.000 537.620 2.000 538.070 ;
        RECT 16.625 538.055 16.955 538.070 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1794.010 2596.650 1794.290 2600.000 ;
        RECT 1795.010 2596.650 1795.290 2596.765 ;
        RECT 1794.010 2596.510 1795.290 2596.650 ;
        RECT 1794.010 2596.000 1794.290 2596.510 ;
        RECT 1795.010 2596.395 1795.290 2596.510 ;
        RECT 3.770 323.835 4.050 324.205 ;
        RECT 3.840 322.845 3.980 323.835 ;
        RECT 3.770 322.475 4.050 322.845 ;
      LAYER via2 ;
        RECT 1795.010 2596.440 1795.290 2596.720 ;
        RECT 3.770 323.880 4.050 324.160 ;
        RECT 3.770 322.520 4.050 322.800 ;
      LAYER met3 ;
        RECT 1794.985 2596.740 1795.315 2596.745 ;
        RECT 1794.985 2596.730 1795.570 2596.740 ;
        RECT 1794.985 2596.430 1795.770 2596.730 ;
        RECT 1794.985 2596.420 1795.570 2596.430 ;
        RECT 1794.985 2596.415 1795.315 2596.420 ;
        RECT 3.745 324.170 4.075 324.185 ;
        RECT 1795.190 324.170 1795.570 324.180 ;
        RECT 3.745 323.870 1795.570 324.170 ;
        RECT 3.745 323.855 4.075 323.870 ;
        RECT 1795.190 323.860 1795.570 323.870 ;
        RECT -4.000 322.810 2.000 323.260 ;
        RECT 3.745 322.810 4.075 322.825 ;
        RECT -4.000 322.510 4.075 322.810 ;
        RECT -4.000 322.060 2.000 322.510 ;
        RECT 3.745 322.495 4.075 322.510 ;
      LAYER via3 ;
        RECT 1795.220 2596.420 1795.540 2596.740 ;
        RECT 1795.220 323.860 1795.540 324.180 ;
      LAYER met4 ;
        RECT 1795.215 2596.415 1795.545 2596.745 ;
        RECT 1795.230 324.185 1795.530 2596.415 ;
        RECT 1795.215 323.855 1795.545 324.185 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1818.010 2596.650 1818.290 2596.765 ;
        RECT 1819.770 2596.650 1820.050 2600.000 ;
        RECT 1818.010 2596.510 1820.050 2596.650 ;
        RECT 1818.010 2596.395 1818.290 2596.510 ;
        RECT 1819.770 2596.000 1820.050 2596.510 ;
        RECT 2.390 109.635 2.670 110.005 ;
        RECT 2.460 107.285 2.600 109.635 ;
        RECT 2.390 106.915 2.670 107.285 ;
      LAYER via2 ;
        RECT 1818.010 2596.440 1818.290 2596.720 ;
        RECT 2.390 109.680 2.670 109.960 ;
        RECT 2.390 106.960 2.670 107.240 ;
      LAYER met3 ;
        RECT 1814.510 2596.730 1814.890 2596.740 ;
        RECT 1817.985 2596.730 1818.315 2596.745 ;
        RECT 1814.510 2596.430 1818.315 2596.730 ;
        RECT 1814.510 2596.420 1814.890 2596.430 ;
        RECT 1817.985 2596.415 1818.315 2596.430 ;
        RECT 2.365 109.970 2.695 109.985 ;
        RECT 1814.510 109.970 1814.890 109.980 ;
        RECT 2.365 109.670 1814.890 109.970 ;
        RECT 2.365 109.655 2.695 109.670 ;
        RECT 1814.510 109.660 1814.890 109.670 ;
        RECT -4.000 107.250 2.000 107.700 ;
        RECT 2.365 107.250 2.695 107.265 ;
        RECT -4.000 106.950 2.695 107.250 ;
        RECT -4.000 106.500 2.000 106.950 ;
        RECT 2.365 106.935 2.695 106.950 ;
      LAYER via3 ;
        RECT 1814.540 2596.420 1814.860 2596.740 ;
        RECT 1814.540 109.660 1814.860 109.980 ;
      LAYER met4 ;
        RECT 1814.535 2596.415 1814.865 2596.745 ;
        RECT 1814.550 109.985 1814.850 2596.415 ;
        RECT 1814.535 109.655 1814.865 109.985 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 949.970 2614.160 950.290 2614.220 ;
        RECT 1880.090 2614.160 1880.410 2614.220 ;
        RECT 949.970 2614.020 1880.410 2614.160 ;
        RECT 949.970 2613.960 950.290 2614.020 ;
        RECT 1880.090 2613.960 1880.410 2614.020 ;
        RECT 1880.090 855.340 1880.410 855.400 ;
        RECT 2900.830 855.340 2901.150 855.400 ;
        RECT 1880.090 855.200 2901.150 855.340 ;
        RECT 1880.090 855.140 1880.410 855.200 ;
        RECT 2900.830 855.140 2901.150 855.200 ;
      LAYER via ;
        RECT 950.000 2613.960 950.260 2614.220 ;
        RECT 1880.120 2613.960 1880.380 2614.220 ;
        RECT 1880.120 855.140 1880.380 855.400 ;
        RECT 2900.860 855.140 2901.120 855.400 ;
      LAYER met2 ;
        RECT 950.000 2613.930 950.260 2614.250 ;
        RECT 1880.120 2613.930 1880.380 2614.250 ;
        RECT 948.070 2599.370 948.350 2600.000 ;
        RECT 950.060 2599.370 950.200 2613.930 ;
        RECT 948.070 2599.230 950.200 2599.370 ;
        RECT 948.070 2596.000 948.350 2599.230 ;
        RECT 1880.180 855.430 1880.320 2613.930 ;
        RECT 1880.120 855.110 1880.380 855.430 ;
        RECT 2900.860 855.110 2901.120 855.430 ;
        RECT 2900.920 850.525 2901.060 855.110 ;
        RECT 2900.850 850.155 2901.130 850.525 ;
      LAYER via2 ;
        RECT 2900.850 850.200 2901.130 850.480 ;
      LAYER met3 ;
        RECT 2900.825 850.490 2901.155 850.505 ;
        RECT 2918.000 850.490 2924.000 850.940 ;
        RECT 2900.825 850.190 2924.000 850.490 ;
        RECT 2900.825 850.175 2901.155 850.190 ;
        RECT 2918.000 849.740 2924.000 850.190 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 973.830 2596.650 974.110 2600.000 ;
        RECT 975.290 2596.650 975.570 2596.765 ;
        RECT 973.830 2596.510 975.570 2596.650 ;
        RECT 973.830 2596.000 974.110 2596.510 ;
        RECT 975.290 2596.395 975.570 2596.510 ;
        RECT 2900.850 2590.955 2901.130 2591.325 ;
        RECT 2900.920 1085.125 2901.060 2590.955 ;
        RECT 2900.850 1084.755 2901.130 1085.125 ;
      LAYER via2 ;
        RECT 975.290 2596.440 975.570 2596.720 ;
        RECT 2900.850 2591.000 2901.130 2591.280 ;
        RECT 2900.850 1084.800 2901.130 1085.080 ;
      LAYER met3 ;
        RECT 975.265 2596.740 975.595 2596.745 ;
        RECT 975.265 2596.730 975.850 2596.740 ;
        RECT 975.265 2596.430 976.050 2596.730 ;
        RECT 975.265 2596.420 975.850 2596.430 ;
        RECT 975.265 2596.415 975.595 2596.420 ;
        RECT 1472.270 2596.050 1472.650 2596.060 ;
        RECT 1496.190 2596.050 1496.570 2596.060 ;
        RECT 1472.270 2595.750 1496.570 2596.050 ;
        RECT 1472.270 2595.740 1472.650 2595.750 ;
        RECT 1496.190 2595.740 1496.570 2595.750 ;
        RECT 975.470 2591.290 975.850 2591.300 ;
        RECT 1472.270 2591.290 1472.650 2591.300 ;
        RECT 975.470 2590.990 1472.650 2591.290 ;
        RECT 975.470 2590.980 975.850 2590.990 ;
        RECT 1472.270 2590.980 1472.650 2590.990 ;
        RECT 1496.190 2591.290 1496.570 2591.300 ;
        RECT 2900.825 2591.290 2901.155 2591.305 ;
        RECT 1496.190 2590.990 2901.155 2591.290 ;
        RECT 1496.190 2590.980 1496.570 2590.990 ;
        RECT 2900.825 2590.975 2901.155 2590.990 ;
        RECT 2900.825 1085.090 2901.155 1085.105 ;
        RECT 2918.000 1085.090 2924.000 1085.540 ;
        RECT 2900.825 1084.790 2924.000 1085.090 ;
        RECT 2900.825 1084.775 2901.155 1084.790 ;
        RECT 2918.000 1084.340 2924.000 1084.790 ;
      LAYER via3 ;
        RECT 975.500 2596.420 975.820 2596.740 ;
        RECT 1472.300 2595.740 1472.620 2596.060 ;
        RECT 1496.220 2595.740 1496.540 2596.060 ;
        RECT 975.500 2590.980 975.820 2591.300 ;
        RECT 1472.300 2590.980 1472.620 2591.300 ;
        RECT 1496.220 2590.980 1496.540 2591.300 ;
      LAYER met4 ;
        RECT 975.495 2596.415 975.825 2596.745 ;
        RECT 975.510 2591.305 975.810 2596.415 ;
        RECT 1472.295 2595.735 1472.625 2596.065 ;
        RECT 1496.215 2595.735 1496.545 2596.065 ;
        RECT 1472.310 2591.305 1472.610 2595.735 ;
        RECT 1496.230 2591.305 1496.530 2595.735 ;
        RECT 975.495 2590.975 975.825 2591.305 ;
        RECT 1472.295 2590.975 1472.625 2591.305 ;
        RECT 1496.215 2590.975 1496.545 2591.305 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 999.130 2596.650 999.410 2600.000 ;
        RECT 999.670 2596.650 999.950 2596.765 ;
        RECT 999.130 2596.510 999.950 2596.650 ;
        RECT 999.130 2596.000 999.410 2596.510 ;
        RECT 999.670 2596.395 999.950 2596.510 ;
        RECT 2899.010 2592.315 2899.290 2592.685 ;
        RECT 2899.080 1319.725 2899.220 2592.315 ;
        RECT 2899.010 1319.355 2899.290 1319.725 ;
      LAYER via2 ;
        RECT 999.670 2596.440 999.950 2596.720 ;
        RECT 2899.010 2592.360 2899.290 2592.640 ;
        RECT 2899.010 1319.400 2899.290 1319.680 ;
      LAYER met3 ;
        RECT 999.645 2596.740 999.975 2596.745 ;
        RECT 999.390 2596.730 999.975 2596.740 ;
        RECT 999.190 2596.430 999.975 2596.730 ;
        RECT 999.390 2596.420 999.975 2596.430 ;
        RECT 999.645 2596.415 999.975 2596.420 ;
        RECT 1174.230 2593.030 1176.370 2593.330 ;
        RECT 999.390 2592.650 999.770 2592.660 ;
        RECT 1174.230 2592.650 1174.530 2593.030 ;
        RECT 999.390 2592.350 1174.530 2592.650 ;
        RECT 1176.070 2592.650 1176.370 2593.030 ;
        RECT 2898.985 2592.650 2899.315 2592.665 ;
        RECT 1176.070 2592.350 2899.315 2592.650 ;
        RECT 999.390 2592.340 999.770 2592.350 ;
        RECT 2898.985 2592.335 2899.315 2592.350 ;
        RECT 2898.985 1319.690 2899.315 1319.705 ;
        RECT 2918.000 1319.690 2924.000 1320.140 ;
        RECT 2898.985 1319.390 2924.000 1319.690 ;
        RECT 2898.985 1319.375 2899.315 1319.390 ;
        RECT 2918.000 1318.940 2924.000 1319.390 ;
      LAYER via3 ;
        RECT 999.420 2596.420 999.740 2596.740 ;
        RECT 999.420 2592.340 999.740 2592.660 ;
      LAYER met4 ;
        RECT 999.415 2596.415 999.745 2596.745 ;
        RECT 999.430 2592.665 999.730 2596.415 ;
        RECT 999.415 2592.335 999.745 2592.665 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1024.890 2596.650 1025.170 2600.000 ;
        RECT 1025.890 2596.650 1026.170 2596.765 ;
        RECT 1024.890 2596.510 1026.170 2596.650 ;
        RECT 1024.890 2596.000 1025.170 2596.510 ;
        RECT 1025.890 2596.395 1026.170 2596.510 ;
        RECT 2916.950 1553.955 2917.230 1554.325 ;
        RECT 2917.020 1553.645 2917.160 1553.955 ;
        RECT 2916.950 1553.275 2917.230 1553.645 ;
      LAYER via2 ;
        RECT 1025.890 2596.440 1026.170 2596.720 ;
        RECT 2916.950 1554.000 2917.230 1554.280 ;
        RECT 2916.950 1553.320 2917.230 1553.600 ;
      LAYER met3 ;
        RECT 1025.865 2596.740 1026.195 2596.745 ;
        RECT 1025.865 2596.730 1026.450 2596.740 ;
        RECT 1025.865 2596.430 1026.650 2596.730 ;
        RECT 1025.865 2596.420 1026.450 2596.430 ;
        RECT 1025.865 2596.415 1026.195 2596.420 ;
        RECT 1026.070 2589.250 1026.450 2589.260 ;
        RECT 1492.510 2589.250 1492.890 2589.260 ;
        RECT 1026.070 2588.950 1492.890 2589.250 ;
        RECT 1026.070 2588.940 1026.450 2588.950 ;
        RECT 1492.510 2588.940 1492.890 2588.950 ;
        RECT 1494.350 2589.250 1494.730 2589.260 ;
        RECT 1836.590 2589.250 1836.970 2589.260 ;
        RECT 1494.350 2588.950 1836.970 2589.250 ;
        RECT 1494.350 2588.940 1494.730 2588.950 ;
        RECT 1836.590 2588.940 1836.970 2588.950 ;
        RECT 1836.590 2588.570 1836.970 2588.580 ;
        RECT 1844.870 2588.570 1845.250 2588.580 ;
        RECT 1836.590 2588.270 1845.250 2588.570 ;
        RECT 1836.590 2588.260 1836.970 2588.270 ;
        RECT 1844.870 2588.260 1845.250 2588.270 ;
        RECT 1844.870 1554.290 1845.250 1554.300 ;
        RECT 2916.925 1554.290 2917.255 1554.305 ;
        RECT 2918.000 1554.290 2924.000 1554.740 ;
        RECT 1844.870 1553.990 1870.050 1554.290 ;
        RECT 1844.870 1553.980 1845.250 1553.990 ;
        RECT 1869.750 1553.610 1870.050 1553.990 ;
        RECT 1918.510 1553.990 1966.650 1554.290 ;
        RECT 1869.750 1553.310 1917.890 1553.610 ;
        RECT 1917.590 1552.930 1917.890 1553.310 ;
        RECT 1918.510 1552.930 1918.810 1553.990 ;
        RECT 1966.350 1553.610 1966.650 1553.990 ;
        RECT 2015.110 1553.990 2063.250 1554.290 ;
        RECT 1966.350 1553.310 2014.490 1553.610 ;
        RECT 1917.590 1552.630 1918.810 1552.930 ;
        RECT 2014.190 1552.930 2014.490 1553.310 ;
        RECT 2015.110 1552.930 2015.410 1553.990 ;
        RECT 2062.950 1553.610 2063.250 1553.990 ;
        RECT 2111.710 1553.990 2159.850 1554.290 ;
        RECT 2062.950 1553.310 2111.090 1553.610 ;
        RECT 2014.190 1552.630 2015.410 1552.930 ;
        RECT 2110.790 1552.930 2111.090 1553.310 ;
        RECT 2111.710 1552.930 2112.010 1553.990 ;
        RECT 2159.550 1553.610 2159.850 1553.990 ;
        RECT 2208.310 1553.990 2256.450 1554.290 ;
        RECT 2159.550 1553.310 2207.690 1553.610 ;
        RECT 2110.790 1552.630 2112.010 1552.930 ;
        RECT 2207.390 1552.930 2207.690 1553.310 ;
        RECT 2208.310 1552.930 2208.610 1553.990 ;
        RECT 2256.150 1553.610 2256.450 1553.990 ;
        RECT 2304.910 1553.990 2353.050 1554.290 ;
        RECT 2256.150 1553.310 2304.290 1553.610 ;
        RECT 2207.390 1552.630 2208.610 1552.930 ;
        RECT 2303.990 1552.930 2304.290 1553.310 ;
        RECT 2304.910 1552.930 2305.210 1553.990 ;
        RECT 2352.750 1553.610 2353.050 1553.990 ;
        RECT 2401.510 1553.990 2449.650 1554.290 ;
        RECT 2352.750 1553.310 2400.890 1553.610 ;
        RECT 2303.990 1552.630 2305.210 1552.930 ;
        RECT 2400.590 1552.930 2400.890 1553.310 ;
        RECT 2401.510 1552.930 2401.810 1553.990 ;
        RECT 2449.350 1553.610 2449.650 1553.990 ;
        RECT 2498.110 1553.990 2546.250 1554.290 ;
        RECT 2449.350 1553.310 2497.490 1553.610 ;
        RECT 2400.590 1552.630 2401.810 1552.930 ;
        RECT 2497.190 1552.930 2497.490 1553.310 ;
        RECT 2498.110 1552.930 2498.410 1553.990 ;
        RECT 2545.950 1553.610 2546.250 1553.990 ;
        RECT 2594.710 1553.990 2642.850 1554.290 ;
        RECT 2545.950 1553.310 2594.090 1553.610 ;
        RECT 2497.190 1552.630 2498.410 1552.930 ;
        RECT 2593.790 1552.930 2594.090 1553.310 ;
        RECT 2594.710 1552.930 2595.010 1553.990 ;
        RECT 2642.550 1553.610 2642.850 1553.990 ;
        RECT 2691.310 1553.990 2739.450 1554.290 ;
        RECT 2642.550 1553.310 2690.690 1553.610 ;
        RECT 2593.790 1552.630 2595.010 1552.930 ;
        RECT 2690.390 1552.930 2690.690 1553.310 ;
        RECT 2691.310 1552.930 2691.610 1553.990 ;
        RECT 2739.150 1553.610 2739.450 1553.990 ;
        RECT 2787.910 1553.990 2836.050 1554.290 ;
        RECT 2739.150 1553.310 2787.290 1553.610 ;
        RECT 2690.390 1552.630 2691.610 1552.930 ;
        RECT 2786.990 1552.930 2787.290 1553.310 ;
        RECT 2787.910 1552.930 2788.210 1553.990 ;
        RECT 2835.750 1553.610 2836.050 1553.990 ;
        RECT 2916.925 1553.990 2924.000 1554.290 ;
        RECT 2916.925 1553.975 2917.255 1553.990 ;
        RECT 2916.925 1553.610 2917.255 1553.625 ;
        RECT 2835.750 1553.310 2883.890 1553.610 ;
        RECT 2786.990 1552.630 2788.210 1552.930 ;
        RECT 2883.590 1552.930 2883.890 1553.310 ;
        RECT 2884.510 1553.310 2917.255 1553.610 ;
        RECT 2918.000 1553.540 2924.000 1553.990 ;
        RECT 2884.510 1552.930 2884.810 1553.310 ;
        RECT 2916.925 1553.295 2917.255 1553.310 ;
        RECT 2883.590 1552.630 2884.810 1552.930 ;
      LAYER via3 ;
        RECT 1026.100 2596.420 1026.420 2596.740 ;
        RECT 1026.100 2588.940 1026.420 2589.260 ;
        RECT 1492.540 2588.940 1492.860 2589.260 ;
        RECT 1494.380 2588.940 1494.700 2589.260 ;
        RECT 1836.620 2588.940 1836.940 2589.260 ;
        RECT 1836.620 2588.260 1836.940 2588.580 ;
        RECT 1844.900 2588.260 1845.220 2588.580 ;
        RECT 1844.900 1553.980 1845.220 1554.300 ;
      LAYER met4 ;
        RECT 1026.095 2596.415 1026.425 2596.745 ;
        RECT 1026.110 2589.265 1026.410 2596.415 ;
        RECT 1026.095 2588.935 1026.425 2589.265 ;
        RECT 1492.535 2589.250 1492.865 2589.265 ;
        RECT 1494.375 2589.250 1494.705 2589.265 ;
        RECT 1492.535 2588.950 1494.705 2589.250 ;
        RECT 1492.535 2588.935 1492.865 2588.950 ;
        RECT 1494.375 2588.935 1494.705 2588.950 ;
        RECT 1836.615 2588.935 1836.945 2589.265 ;
        RECT 1836.630 2588.585 1836.930 2588.935 ;
        RECT 1836.615 2588.255 1836.945 2588.585 ;
        RECT 1844.895 2588.255 1845.225 2588.585 ;
        RECT 1844.910 1554.305 1845.210 2588.255 ;
        RECT 1844.895 1553.975 1845.225 1554.305 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1851.570 2593.420 1851.890 2593.480 ;
        RECT 1876.410 2593.420 1876.730 2593.480 ;
        RECT 1851.570 2593.280 1876.730 2593.420 ;
        RECT 1851.570 2593.220 1851.890 2593.280 ;
        RECT 1876.410 2593.220 1876.730 2593.280 ;
      LAYER via ;
        RECT 1851.600 2593.220 1851.860 2593.480 ;
        RECT 1876.440 2593.220 1876.700 2593.480 ;
      LAYER met2 ;
        RECT 1050.650 2596.650 1050.930 2600.000 ;
        RECT 1051.650 2596.650 1051.930 2596.765 ;
        RECT 1050.650 2596.510 1051.930 2596.650 ;
        RECT 1050.650 2596.000 1050.930 2596.510 ;
        RECT 1051.650 2596.395 1051.930 2596.510 ;
        RECT 1876.430 2593.675 1876.710 2594.045 ;
        RECT 1897.130 2593.675 1897.410 2594.045 ;
        RECT 2028.760 2593.790 2029.360 2593.930 ;
        RECT 1876.500 2593.510 1876.640 2593.675 ;
        RECT 1851.600 2593.365 1851.860 2593.510 ;
        RECT 1851.590 2592.995 1851.870 2593.365 ;
        RECT 1876.440 2593.190 1876.700 2593.510 ;
        RECT 1897.200 2593.250 1897.340 2593.675 ;
        RECT 2028.760 2593.365 2028.900 2593.790 ;
        RECT 1898.050 2593.250 1898.330 2593.365 ;
        RECT 1897.200 2593.110 1898.330 2593.250 ;
        RECT 1898.050 2592.995 1898.330 2593.110 ;
        RECT 1932.090 2592.995 1932.370 2593.365 ;
        RECT 1996.490 2592.995 1996.770 2593.365 ;
        RECT 2028.690 2592.995 2028.970 2593.365 ;
        RECT 1932.160 2589.285 1932.300 2592.995 ;
        RECT 1996.560 2589.285 1996.700 2592.995 ;
        RECT 2029.220 2589.965 2029.360 2593.790 ;
        RECT 2125.360 2593.790 2125.960 2593.930 ;
        RECT 2125.360 2593.365 2125.500 2593.790 ;
        RECT 2090.330 2592.995 2090.610 2593.365 ;
        RECT 2125.290 2592.995 2125.570 2593.365 ;
        RECT 2090.400 2589.965 2090.540 2592.995 ;
        RECT 2125.820 2589.965 2125.960 2593.790 ;
        RECT 2221.960 2593.790 2222.560 2593.930 ;
        RECT 2221.960 2593.365 2222.100 2593.790 ;
        RECT 2186.930 2592.995 2187.210 2593.365 ;
        RECT 2221.890 2592.995 2222.170 2593.365 ;
        RECT 2187.000 2589.965 2187.140 2592.995 ;
        RECT 2222.420 2589.965 2222.560 2593.790 ;
        RECT 2318.560 2593.790 2319.160 2593.930 ;
        RECT 2318.560 2593.365 2318.700 2593.790 ;
        RECT 2283.530 2592.995 2283.810 2593.365 ;
        RECT 2318.490 2592.995 2318.770 2593.365 ;
        RECT 2283.600 2589.965 2283.740 2592.995 ;
        RECT 2319.020 2589.965 2319.160 2593.790 ;
        RECT 2415.160 2593.790 2415.760 2593.930 ;
        RECT 2415.160 2593.365 2415.300 2593.790 ;
        RECT 2380.130 2592.995 2380.410 2593.365 ;
        RECT 2415.090 2592.995 2415.370 2593.365 ;
        RECT 2380.200 2589.965 2380.340 2592.995 ;
        RECT 2415.620 2589.965 2415.760 2593.790 ;
        RECT 2511.760 2593.790 2512.360 2593.930 ;
        RECT 2511.760 2593.365 2511.900 2593.790 ;
        RECT 2476.730 2592.995 2477.010 2593.365 ;
        RECT 2511.690 2592.995 2511.970 2593.365 ;
        RECT 2476.800 2589.965 2476.940 2592.995 ;
        RECT 2512.220 2589.965 2512.360 2593.790 ;
        RECT 2573.330 2592.995 2573.610 2593.365 ;
        RECT 2766.990 2592.995 2767.270 2593.365 ;
        RECT 2814.830 2592.995 2815.110 2593.365 ;
        RECT 2900.390 2592.995 2900.670 2593.365 ;
        RECT 2573.400 2589.965 2573.540 2592.995 ;
        RECT 2767.060 2589.965 2767.200 2592.995 ;
        RECT 2814.900 2589.965 2815.040 2592.995 ;
        RECT 2029.150 2589.595 2029.430 2589.965 ;
        RECT 2090.330 2589.595 2090.610 2589.965 ;
        RECT 2125.750 2589.595 2126.030 2589.965 ;
        RECT 2186.930 2589.595 2187.210 2589.965 ;
        RECT 2222.350 2589.595 2222.630 2589.965 ;
        RECT 2283.530 2589.595 2283.810 2589.965 ;
        RECT 2318.950 2589.595 2319.230 2589.965 ;
        RECT 2380.130 2589.595 2380.410 2589.965 ;
        RECT 2415.550 2589.595 2415.830 2589.965 ;
        RECT 2476.730 2589.595 2477.010 2589.965 ;
        RECT 2512.150 2589.595 2512.430 2589.965 ;
        RECT 2573.330 2589.595 2573.610 2589.965 ;
        RECT 2766.990 2589.595 2767.270 2589.965 ;
        RECT 2814.830 2589.595 2815.110 2589.965 ;
        RECT 1932.090 2588.915 1932.370 2589.285 ;
        RECT 1996.490 2588.915 1996.770 2589.285 ;
        RECT 2900.460 1789.605 2900.600 2592.995 ;
        RECT 2900.390 1789.235 2900.670 1789.605 ;
      LAYER via2 ;
        RECT 1051.650 2596.440 1051.930 2596.720 ;
        RECT 1876.430 2593.720 1876.710 2594.000 ;
        RECT 1897.130 2593.720 1897.410 2594.000 ;
        RECT 1851.590 2593.040 1851.870 2593.320 ;
        RECT 1898.050 2593.040 1898.330 2593.320 ;
        RECT 1932.090 2593.040 1932.370 2593.320 ;
        RECT 1996.490 2593.040 1996.770 2593.320 ;
        RECT 2028.690 2593.040 2028.970 2593.320 ;
        RECT 2090.330 2593.040 2090.610 2593.320 ;
        RECT 2125.290 2593.040 2125.570 2593.320 ;
        RECT 2186.930 2593.040 2187.210 2593.320 ;
        RECT 2221.890 2593.040 2222.170 2593.320 ;
        RECT 2283.530 2593.040 2283.810 2593.320 ;
        RECT 2318.490 2593.040 2318.770 2593.320 ;
        RECT 2380.130 2593.040 2380.410 2593.320 ;
        RECT 2415.090 2593.040 2415.370 2593.320 ;
        RECT 2476.730 2593.040 2477.010 2593.320 ;
        RECT 2511.690 2593.040 2511.970 2593.320 ;
        RECT 2573.330 2593.040 2573.610 2593.320 ;
        RECT 2766.990 2593.040 2767.270 2593.320 ;
        RECT 2814.830 2593.040 2815.110 2593.320 ;
        RECT 2900.390 2593.040 2900.670 2593.320 ;
        RECT 2029.150 2589.640 2029.430 2589.920 ;
        RECT 2090.330 2589.640 2090.610 2589.920 ;
        RECT 2125.750 2589.640 2126.030 2589.920 ;
        RECT 2186.930 2589.640 2187.210 2589.920 ;
        RECT 2222.350 2589.640 2222.630 2589.920 ;
        RECT 2283.530 2589.640 2283.810 2589.920 ;
        RECT 2318.950 2589.640 2319.230 2589.920 ;
        RECT 2380.130 2589.640 2380.410 2589.920 ;
        RECT 2415.550 2589.640 2415.830 2589.920 ;
        RECT 2476.730 2589.640 2477.010 2589.920 ;
        RECT 2512.150 2589.640 2512.430 2589.920 ;
        RECT 2573.330 2589.640 2573.610 2589.920 ;
        RECT 2766.990 2589.640 2767.270 2589.920 ;
        RECT 2814.830 2589.640 2815.110 2589.920 ;
        RECT 1932.090 2588.960 1932.370 2589.240 ;
        RECT 1996.490 2588.960 1996.770 2589.240 ;
        RECT 2900.390 1789.280 2900.670 1789.560 ;
      LAYER met3 ;
        RECT 1546.790 2597.410 1547.170 2597.420 ;
        RECT 1566.110 2597.410 1566.490 2597.420 ;
        RECT 1546.790 2597.110 1566.490 2597.410 ;
        RECT 1546.790 2597.100 1547.170 2597.110 ;
        RECT 1566.110 2597.100 1566.490 2597.110 ;
        RECT 1051.625 2596.740 1051.955 2596.745 ;
        RECT 1051.625 2596.730 1052.210 2596.740 ;
        RECT 1051.625 2596.430 1052.410 2596.730 ;
        RECT 1051.625 2596.420 1052.210 2596.430 ;
        RECT 1051.625 2596.415 1051.955 2596.420 ;
        RECT 1172.350 2596.050 1172.730 2596.060 ;
        RECT 1183.390 2596.050 1183.770 2596.060 ;
        RECT 1172.350 2595.750 1183.770 2596.050 ;
        RECT 1172.350 2595.740 1172.730 2595.750 ;
        RECT 1183.390 2595.740 1183.770 2595.750 ;
        RECT 1315.870 2596.050 1316.250 2596.060 ;
        RECT 1327.830 2596.050 1328.210 2596.060 ;
        RECT 1315.870 2595.750 1328.210 2596.050 ;
        RECT 1315.870 2595.740 1316.250 2595.750 ;
        RECT 1327.830 2595.740 1328.210 2595.750 ;
        RECT 1566.110 2596.050 1566.490 2596.060 ;
        RECT 1613.950 2596.050 1614.330 2596.060 ;
        RECT 1566.110 2595.750 1614.330 2596.050 ;
        RECT 1566.110 2595.740 1566.490 2595.750 ;
        RECT 1613.950 2595.740 1614.330 2595.750 ;
        RECT 1876.405 2594.010 1876.735 2594.025 ;
        RECT 1897.105 2594.010 1897.435 2594.025 ;
        RECT 1677.470 2593.710 1679.610 2594.010 ;
        RECT 1051.830 2593.330 1052.210 2593.340 ;
        RECT 1172.350 2593.330 1172.730 2593.340 ;
        RECT 1051.830 2593.030 1172.730 2593.330 ;
        RECT 1051.830 2593.020 1052.210 2593.030 ;
        RECT 1172.350 2593.020 1172.730 2593.030 ;
        RECT 1219.270 2593.330 1219.650 2593.340 ;
        RECT 1221.110 2593.330 1221.490 2593.340 ;
        RECT 1219.270 2593.030 1221.490 2593.330 ;
        RECT 1219.270 2593.020 1219.650 2593.030 ;
        RECT 1221.110 2593.020 1221.490 2593.030 ;
        RECT 1268.950 2593.330 1269.330 2593.340 ;
        RECT 1315.870 2593.330 1316.250 2593.340 ;
        RECT 1268.950 2593.030 1316.250 2593.330 ;
        RECT 1268.950 2593.020 1269.330 2593.030 ;
        RECT 1315.870 2593.020 1316.250 2593.030 ;
        RECT 1365.550 2593.330 1365.930 2593.340 ;
        RECT 1415.230 2593.330 1415.610 2593.340 ;
        RECT 1365.550 2593.030 1415.610 2593.330 ;
        RECT 1365.550 2593.020 1365.930 2593.030 ;
        RECT 1415.230 2593.020 1415.610 2593.030 ;
        RECT 1473.190 2593.330 1473.570 2593.340 ;
        RECT 1493.430 2593.330 1493.810 2593.340 ;
        RECT 1473.190 2593.030 1493.810 2593.330 ;
        RECT 1473.190 2593.020 1473.570 2593.030 ;
        RECT 1493.430 2593.020 1493.810 2593.030 ;
        RECT 1509.990 2593.330 1510.370 2593.340 ;
        RECT 1545.870 2593.330 1546.250 2593.340 ;
        RECT 1509.990 2593.030 1546.250 2593.330 ;
        RECT 1509.990 2593.020 1510.370 2593.030 ;
        RECT 1545.870 2593.020 1546.250 2593.030 ;
        RECT 1613.950 2593.330 1614.330 2593.340 ;
        RECT 1677.470 2593.330 1677.770 2593.710 ;
        RECT 1613.950 2593.030 1677.770 2593.330 ;
        RECT 1679.310 2593.330 1679.610 2593.710 ;
        RECT 1876.405 2593.710 1897.435 2594.010 ;
        RECT 1876.405 2593.695 1876.735 2593.710 ;
        RECT 1897.105 2593.695 1897.435 2593.710 ;
        RECT 1851.565 2593.330 1851.895 2593.345 ;
        RECT 1679.310 2593.030 1851.895 2593.330 ;
        RECT 1613.950 2593.020 1614.330 2593.030 ;
        RECT 1851.565 2593.015 1851.895 2593.030 ;
        RECT 1898.025 2593.330 1898.355 2593.345 ;
        RECT 1932.065 2593.330 1932.395 2593.345 ;
        RECT 1898.025 2593.030 1932.395 2593.330 ;
        RECT 1898.025 2593.015 1898.355 2593.030 ;
        RECT 1932.065 2593.015 1932.395 2593.030 ;
        RECT 1996.465 2593.330 1996.795 2593.345 ;
        RECT 2028.665 2593.330 2028.995 2593.345 ;
        RECT 1996.465 2593.030 2028.995 2593.330 ;
        RECT 1996.465 2593.015 1996.795 2593.030 ;
        RECT 2028.665 2593.015 2028.995 2593.030 ;
        RECT 2090.305 2593.330 2090.635 2593.345 ;
        RECT 2125.265 2593.330 2125.595 2593.345 ;
        RECT 2090.305 2593.030 2125.595 2593.330 ;
        RECT 2090.305 2593.015 2090.635 2593.030 ;
        RECT 2125.265 2593.015 2125.595 2593.030 ;
        RECT 2186.905 2593.330 2187.235 2593.345 ;
        RECT 2221.865 2593.330 2222.195 2593.345 ;
        RECT 2186.905 2593.030 2222.195 2593.330 ;
        RECT 2186.905 2593.015 2187.235 2593.030 ;
        RECT 2221.865 2593.015 2222.195 2593.030 ;
        RECT 2283.505 2593.330 2283.835 2593.345 ;
        RECT 2318.465 2593.330 2318.795 2593.345 ;
        RECT 2283.505 2593.030 2318.795 2593.330 ;
        RECT 2283.505 2593.015 2283.835 2593.030 ;
        RECT 2318.465 2593.015 2318.795 2593.030 ;
        RECT 2380.105 2593.330 2380.435 2593.345 ;
        RECT 2415.065 2593.330 2415.395 2593.345 ;
        RECT 2380.105 2593.030 2415.395 2593.330 ;
        RECT 2380.105 2593.015 2380.435 2593.030 ;
        RECT 2415.065 2593.015 2415.395 2593.030 ;
        RECT 2476.705 2593.330 2477.035 2593.345 ;
        RECT 2511.665 2593.330 2511.995 2593.345 ;
        RECT 2476.705 2593.030 2511.995 2593.330 ;
        RECT 2476.705 2593.015 2477.035 2593.030 ;
        RECT 2511.665 2593.015 2511.995 2593.030 ;
        RECT 2573.305 2593.330 2573.635 2593.345 ;
        RECT 2766.965 2593.330 2767.295 2593.345 ;
        RECT 2573.305 2593.030 2767.295 2593.330 ;
        RECT 2573.305 2593.015 2573.635 2593.030 ;
        RECT 2766.965 2593.015 2767.295 2593.030 ;
        RECT 2814.805 2593.330 2815.135 2593.345 ;
        RECT 2900.365 2593.330 2900.695 2593.345 ;
        RECT 2814.805 2593.030 2900.695 2593.330 ;
        RECT 2814.805 2593.015 2815.135 2593.030 ;
        RECT 2900.365 2593.015 2900.695 2593.030 ;
        RECT 1183.390 2589.930 1183.770 2589.940 ;
        RECT 1216.510 2589.930 1216.890 2589.940 ;
        RECT 1183.390 2589.630 1216.890 2589.930 ;
        RECT 1183.390 2589.620 1183.770 2589.630 ;
        RECT 1216.510 2589.620 1216.890 2589.630 ;
        RECT 1222.030 2589.930 1222.410 2589.940 ;
        RECT 1268.950 2589.930 1269.330 2589.940 ;
        RECT 1222.030 2589.630 1269.330 2589.930 ;
        RECT 1222.030 2589.620 1222.410 2589.630 ;
        RECT 1268.950 2589.620 1269.330 2589.630 ;
        RECT 1327.830 2589.930 1328.210 2589.940 ;
        RECT 1365.550 2589.930 1365.930 2589.940 ;
        RECT 1327.830 2589.630 1365.930 2589.930 ;
        RECT 1327.830 2589.620 1328.210 2589.630 ;
        RECT 1365.550 2589.620 1365.930 2589.630 ;
        RECT 1415.230 2589.930 1415.610 2589.940 ;
        RECT 1473.190 2589.930 1473.570 2589.940 ;
        RECT 1415.230 2589.630 1473.570 2589.930 ;
        RECT 1415.230 2589.620 1415.610 2589.630 ;
        RECT 1473.190 2589.620 1473.570 2589.630 ;
        RECT 1494.350 2589.930 1494.730 2589.940 ;
        RECT 1509.990 2589.930 1510.370 2589.940 ;
        RECT 1494.350 2589.630 1510.370 2589.930 ;
        RECT 1494.350 2589.620 1494.730 2589.630 ;
        RECT 1509.990 2589.620 1510.370 2589.630 ;
        RECT 2029.125 2589.930 2029.455 2589.945 ;
        RECT 2090.305 2589.930 2090.635 2589.945 ;
        RECT 2029.125 2589.630 2090.635 2589.930 ;
        RECT 2029.125 2589.615 2029.455 2589.630 ;
        RECT 2090.305 2589.615 2090.635 2589.630 ;
        RECT 2125.725 2589.930 2126.055 2589.945 ;
        RECT 2186.905 2589.930 2187.235 2589.945 ;
        RECT 2125.725 2589.630 2187.235 2589.930 ;
        RECT 2125.725 2589.615 2126.055 2589.630 ;
        RECT 2186.905 2589.615 2187.235 2589.630 ;
        RECT 2222.325 2589.930 2222.655 2589.945 ;
        RECT 2283.505 2589.930 2283.835 2589.945 ;
        RECT 2222.325 2589.630 2283.835 2589.930 ;
        RECT 2222.325 2589.615 2222.655 2589.630 ;
        RECT 2283.505 2589.615 2283.835 2589.630 ;
        RECT 2318.925 2589.930 2319.255 2589.945 ;
        RECT 2380.105 2589.930 2380.435 2589.945 ;
        RECT 2318.925 2589.630 2380.435 2589.930 ;
        RECT 2318.925 2589.615 2319.255 2589.630 ;
        RECT 2380.105 2589.615 2380.435 2589.630 ;
        RECT 2415.525 2589.930 2415.855 2589.945 ;
        RECT 2476.705 2589.930 2477.035 2589.945 ;
        RECT 2415.525 2589.630 2477.035 2589.930 ;
        RECT 2415.525 2589.615 2415.855 2589.630 ;
        RECT 2476.705 2589.615 2477.035 2589.630 ;
        RECT 2512.125 2589.930 2512.455 2589.945 ;
        RECT 2573.305 2589.930 2573.635 2589.945 ;
        RECT 2512.125 2589.630 2573.635 2589.930 ;
        RECT 2512.125 2589.615 2512.455 2589.630 ;
        RECT 2573.305 2589.615 2573.635 2589.630 ;
        RECT 2766.965 2589.930 2767.295 2589.945 ;
        RECT 2814.805 2589.930 2815.135 2589.945 ;
        RECT 2766.965 2589.630 2815.135 2589.930 ;
        RECT 2766.965 2589.615 2767.295 2589.630 ;
        RECT 2814.805 2589.615 2815.135 2589.630 ;
        RECT 1932.065 2589.250 1932.395 2589.265 ;
        RECT 1996.465 2589.250 1996.795 2589.265 ;
        RECT 1932.065 2588.950 1996.795 2589.250 ;
        RECT 1932.065 2588.935 1932.395 2588.950 ;
        RECT 1996.465 2588.935 1996.795 2588.950 ;
        RECT 2900.365 1789.570 2900.695 1789.585 ;
        RECT 2918.000 1789.570 2924.000 1790.020 ;
        RECT 2900.365 1789.270 2924.000 1789.570 ;
        RECT 2900.365 1789.255 2900.695 1789.270 ;
        RECT 2918.000 1788.820 2924.000 1789.270 ;
      LAYER via3 ;
        RECT 1546.820 2597.100 1547.140 2597.420 ;
        RECT 1566.140 2597.100 1566.460 2597.420 ;
        RECT 1051.860 2596.420 1052.180 2596.740 ;
        RECT 1172.380 2595.740 1172.700 2596.060 ;
        RECT 1183.420 2595.740 1183.740 2596.060 ;
        RECT 1315.900 2595.740 1316.220 2596.060 ;
        RECT 1327.860 2595.740 1328.180 2596.060 ;
        RECT 1566.140 2595.740 1566.460 2596.060 ;
        RECT 1613.980 2595.740 1614.300 2596.060 ;
        RECT 1051.860 2593.020 1052.180 2593.340 ;
        RECT 1172.380 2593.020 1172.700 2593.340 ;
        RECT 1219.300 2593.020 1219.620 2593.340 ;
        RECT 1221.140 2593.020 1221.460 2593.340 ;
        RECT 1268.980 2593.020 1269.300 2593.340 ;
        RECT 1315.900 2593.020 1316.220 2593.340 ;
        RECT 1365.580 2593.020 1365.900 2593.340 ;
        RECT 1415.260 2593.020 1415.580 2593.340 ;
        RECT 1473.220 2593.020 1473.540 2593.340 ;
        RECT 1493.460 2593.020 1493.780 2593.340 ;
        RECT 1510.020 2593.020 1510.340 2593.340 ;
        RECT 1545.900 2593.020 1546.220 2593.340 ;
        RECT 1613.980 2593.020 1614.300 2593.340 ;
        RECT 1183.420 2589.620 1183.740 2589.940 ;
        RECT 1216.540 2589.620 1216.860 2589.940 ;
        RECT 1222.060 2589.620 1222.380 2589.940 ;
        RECT 1268.980 2589.620 1269.300 2589.940 ;
        RECT 1327.860 2589.620 1328.180 2589.940 ;
        RECT 1365.580 2589.620 1365.900 2589.940 ;
        RECT 1415.260 2589.620 1415.580 2589.940 ;
        RECT 1473.220 2589.620 1473.540 2589.940 ;
        RECT 1494.380 2589.620 1494.700 2589.940 ;
        RECT 1510.020 2589.620 1510.340 2589.940 ;
      LAYER met4 ;
        RECT 1546.815 2597.095 1547.145 2597.425 ;
        RECT 1566.135 2597.095 1566.465 2597.425 ;
        RECT 1051.855 2596.415 1052.185 2596.745 ;
        RECT 1051.870 2593.345 1052.170 2596.415 ;
        RECT 1172.375 2595.735 1172.705 2596.065 ;
        RECT 1183.415 2595.735 1183.745 2596.065 ;
        RECT 1315.895 2595.735 1316.225 2596.065 ;
        RECT 1327.855 2595.735 1328.185 2596.065 ;
        RECT 1172.390 2593.345 1172.690 2595.735 ;
        RECT 1051.855 2593.015 1052.185 2593.345 ;
        RECT 1172.375 2593.015 1172.705 2593.345 ;
        RECT 1183.430 2589.945 1183.730 2595.735 ;
        RECT 1315.910 2593.345 1316.210 2595.735 ;
        RECT 1219.295 2593.330 1219.625 2593.345 ;
        RECT 1216.550 2593.030 1219.625 2593.330 ;
        RECT 1216.550 2589.945 1216.850 2593.030 ;
        RECT 1219.295 2593.015 1219.625 2593.030 ;
        RECT 1221.135 2593.015 1221.465 2593.345 ;
        RECT 1268.975 2593.015 1269.305 2593.345 ;
        RECT 1315.895 2593.015 1316.225 2593.345 ;
        RECT 1221.150 2592.650 1221.450 2593.015 ;
        RECT 1221.150 2592.350 1222.370 2592.650 ;
        RECT 1222.070 2589.945 1222.370 2592.350 ;
        RECT 1268.990 2589.945 1269.290 2593.015 ;
        RECT 1327.870 2589.945 1328.170 2595.735 ;
        RECT 1365.575 2593.015 1365.905 2593.345 ;
        RECT 1415.255 2593.015 1415.585 2593.345 ;
        RECT 1473.215 2593.015 1473.545 2593.345 ;
        RECT 1493.455 2593.015 1493.785 2593.345 ;
        RECT 1510.015 2593.015 1510.345 2593.345 ;
        RECT 1545.895 2593.015 1546.225 2593.345 ;
        RECT 1365.590 2589.945 1365.890 2593.015 ;
        RECT 1415.270 2589.945 1415.570 2593.015 ;
        RECT 1473.230 2589.945 1473.530 2593.015 ;
        RECT 1493.470 2592.650 1493.770 2593.015 ;
        RECT 1493.470 2592.350 1494.690 2592.650 ;
        RECT 1494.390 2589.945 1494.690 2592.350 ;
        RECT 1510.030 2589.945 1510.330 2593.015 ;
        RECT 1545.910 2592.650 1546.210 2593.015 ;
        RECT 1546.830 2592.650 1547.130 2597.095 ;
        RECT 1566.150 2596.065 1566.450 2597.095 ;
        RECT 1566.135 2595.735 1566.465 2596.065 ;
        RECT 1613.975 2595.735 1614.305 2596.065 ;
        RECT 1613.990 2593.345 1614.290 2595.735 ;
        RECT 1613.975 2593.015 1614.305 2593.345 ;
        RECT 1545.910 2592.350 1547.130 2592.650 ;
        RECT 1183.415 2589.615 1183.745 2589.945 ;
        RECT 1216.535 2589.615 1216.865 2589.945 ;
        RECT 1222.055 2589.615 1222.385 2589.945 ;
        RECT 1268.975 2589.615 1269.305 2589.945 ;
        RECT 1327.855 2589.615 1328.185 2589.945 ;
        RECT 1365.575 2589.615 1365.905 2589.945 ;
        RECT 1415.255 2589.615 1415.585 2589.945 ;
        RECT 1473.215 2589.615 1473.545 2589.945 ;
        RECT 1494.375 2589.615 1494.705 2589.945 ;
        RECT 1510.015 2589.615 1510.345 2589.945 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1077.850 2597.840 1078.170 2597.900 ;
        RECT 1853.410 2597.840 1853.730 2597.900 ;
        RECT 1077.850 2597.700 1853.730 2597.840 ;
        RECT 1077.850 2597.640 1078.170 2597.700 ;
        RECT 1853.410 2597.640 1853.730 2597.700 ;
        RECT 1853.410 2028.340 1853.730 2028.400 ;
        RECT 2899.450 2028.340 2899.770 2028.400 ;
        RECT 1853.410 2028.200 2899.770 2028.340 ;
        RECT 1853.410 2028.140 1853.730 2028.200 ;
        RECT 2899.450 2028.140 2899.770 2028.200 ;
      LAYER via ;
        RECT 1077.880 2597.640 1078.140 2597.900 ;
        RECT 1853.440 2597.640 1853.700 2597.900 ;
        RECT 1853.440 2028.140 1853.700 2028.400 ;
        RECT 2899.480 2028.140 2899.740 2028.400 ;
      LAYER met2 ;
        RECT 1076.410 2598.010 1076.690 2600.000 ;
        RECT 1076.410 2597.930 1078.080 2598.010 ;
        RECT 1076.410 2597.870 1078.140 2597.930 ;
        RECT 1076.410 2596.000 1076.690 2597.870 ;
        RECT 1077.880 2597.610 1078.140 2597.870 ;
        RECT 1853.440 2597.610 1853.700 2597.930 ;
        RECT 1853.500 2028.430 1853.640 2597.610 ;
        RECT 1853.440 2028.110 1853.700 2028.430 ;
        RECT 2899.480 2028.110 2899.740 2028.430 ;
        RECT 2899.540 2024.205 2899.680 2028.110 ;
        RECT 2899.470 2023.835 2899.750 2024.205 ;
      LAYER via2 ;
        RECT 2899.470 2023.880 2899.750 2024.160 ;
      LAYER met3 ;
        RECT 2899.445 2024.170 2899.775 2024.185 ;
        RECT 2918.000 2024.170 2924.000 2024.620 ;
        RECT 2899.445 2023.870 2924.000 2024.170 ;
        RECT 2899.445 2023.855 2899.775 2023.870 ;
        RECT 2918.000 2023.420 2924.000 2023.870 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1103.610 2603.960 1103.930 2604.020 ;
        RECT 1854.790 2603.960 1855.110 2604.020 ;
        RECT 1103.610 2603.820 1855.110 2603.960 ;
        RECT 1103.610 2603.760 1103.930 2603.820 ;
        RECT 1854.790 2603.760 1855.110 2603.820 ;
        RECT 1854.790 2262.940 1855.110 2263.000 ;
        RECT 2899.450 2262.940 2899.770 2263.000 ;
        RECT 1854.790 2262.800 2899.770 2262.940 ;
        RECT 1854.790 2262.740 1855.110 2262.800 ;
        RECT 2899.450 2262.740 2899.770 2262.800 ;
      LAYER via ;
        RECT 1103.640 2603.760 1103.900 2604.020 ;
        RECT 1854.820 2603.760 1855.080 2604.020 ;
        RECT 1854.820 2262.740 1855.080 2263.000 ;
        RECT 2899.480 2262.740 2899.740 2263.000 ;
      LAYER met2 ;
        RECT 1103.640 2603.730 1103.900 2604.050 ;
        RECT 1854.820 2603.730 1855.080 2604.050 ;
        RECT 1101.710 2599.370 1101.990 2600.000 ;
        RECT 1103.700 2599.370 1103.840 2603.730 ;
        RECT 1101.710 2599.230 1103.840 2599.370 ;
        RECT 1101.710 2596.000 1101.990 2599.230 ;
        RECT 1854.880 2263.030 1855.020 2603.730 ;
        RECT 1854.820 2262.710 1855.080 2263.030 ;
        RECT 2899.480 2262.710 2899.740 2263.030 ;
        RECT 2899.540 2258.805 2899.680 2262.710 ;
        RECT 2899.470 2258.435 2899.750 2258.805 ;
      LAYER via2 ;
        RECT 2899.470 2258.480 2899.750 2258.760 ;
      LAYER met3 ;
        RECT 2899.445 2258.770 2899.775 2258.785 ;
        RECT 2918.000 2258.770 2924.000 2259.220 ;
        RECT 2899.445 2258.470 2924.000 2258.770 ;
        RECT 2899.445 2258.455 2899.775 2258.470 ;
        RECT 2918.000 2258.020 2924.000 2258.470 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 633.030 46.140 633.350 46.200 ;
        RECT 1064.510 46.140 1064.830 46.200 ;
        RECT 633.030 46.000 1064.830 46.140 ;
        RECT 633.030 45.940 633.350 46.000 ;
        RECT 1064.510 45.940 1064.830 46.000 ;
      LAYER via ;
        RECT 633.060 45.940 633.320 46.200 ;
        RECT 1064.540 45.940 1064.800 46.200 ;
      LAYER met2 ;
        RECT 1067.210 1100.650 1067.490 1104.000 ;
        RECT 1065.980 1100.510 1067.490 1100.650 ;
        RECT 1065.980 1072.770 1066.120 1100.510 ;
        RECT 1067.210 1100.000 1067.490 1100.510 ;
        RECT 1064.600 1072.630 1066.120 1072.770 ;
        RECT 1064.600 46.230 1064.740 1072.630 ;
        RECT 633.060 45.910 633.320 46.230 ;
        RECT 1064.540 45.910 1064.800 46.230 ;
        RECT 633.120 2.000 633.260 45.910 ;
        RECT 632.910 -4.000 633.470 2.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1679.530 1088.580 1679.850 1088.640 ;
        RECT 1682.750 1088.580 1683.070 1088.640 ;
        RECT 1679.530 1088.440 1683.070 1088.580 ;
        RECT 1679.530 1088.380 1679.850 1088.440 ;
        RECT 1682.750 1088.380 1683.070 1088.440 ;
        RECT 1682.750 54.300 1683.070 54.360 ;
        RECT 2415.070 54.300 2415.390 54.360 ;
        RECT 1682.750 54.160 2415.390 54.300 ;
        RECT 1682.750 54.100 1683.070 54.160 ;
        RECT 2415.070 54.100 2415.390 54.160 ;
      LAYER via ;
        RECT 1679.560 1088.380 1679.820 1088.640 ;
        RECT 1682.780 1088.380 1683.040 1088.640 ;
        RECT 1682.780 54.100 1683.040 54.360 ;
        RECT 2415.100 54.100 2415.360 54.360 ;
      LAYER met2 ;
        RECT 1679.470 1100.580 1679.750 1104.000 ;
        RECT 1679.470 1100.000 1679.760 1100.580 ;
        RECT 1679.620 1088.670 1679.760 1100.000 ;
        RECT 1679.560 1088.350 1679.820 1088.670 ;
        RECT 1682.780 1088.350 1683.040 1088.670 ;
        RECT 1682.840 54.390 1682.980 1088.350 ;
        RECT 1682.780 54.070 1683.040 54.390 ;
        RECT 2415.100 54.070 2415.360 54.390 ;
        RECT 2415.160 2.450 2415.300 54.070 ;
        RECT 2415.160 2.310 2417.600 2.450 ;
        RECT 2417.460 2.000 2417.600 2.310 ;
        RECT 2417.250 -4.000 2417.810 2.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1685.510 1087.220 1685.830 1087.280 ;
        RECT 1690.110 1087.220 1690.430 1087.280 ;
        RECT 1685.510 1087.080 1690.430 1087.220 ;
        RECT 1685.510 1087.020 1685.830 1087.080 ;
        RECT 1690.110 1087.020 1690.430 1087.080 ;
        RECT 1690.110 53.960 1690.430 54.020 ;
        RECT 2429.330 53.960 2429.650 54.020 ;
        RECT 1690.110 53.820 2429.650 53.960 ;
        RECT 1690.110 53.760 1690.430 53.820 ;
        RECT 2429.330 53.760 2429.650 53.820 ;
        RECT 2429.330 2.620 2429.650 2.680 ;
        RECT 2434.850 2.620 2435.170 2.680 ;
        RECT 2429.330 2.480 2435.170 2.620 ;
        RECT 2429.330 2.420 2429.650 2.480 ;
        RECT 2434.850 2.420 2435.170 2.480 ;
      LAYER via ;
        RECT 1685.540 1087.020 1685.800 1087.280 ;
        RECT 1690.140 1087.020 1690.400 1087.280 ;
        RECT 1690.140 53.760 1690.400 54.020 ;
        RECT 2429.360 53.760 2429.620 54.020 ;
        RECT 2429.360 2.420 2429.620 2.680 ;
        RECT 2434.880 2.420 2435.140 2.680 ;
      LAYER met2 ;
        RECT 1685.450 1100.580 1685.730 1104.000 ;
        RECT 1685.450 1100.000 1685.740 1100.580 ;
        RECT 1685.600 1087.310 1685.740 1100.000 ;
        RECT 1685.540 1086.990 1685.800 1087.310 ;
        RECT 1690.140 1086.990 1690.400 1087.310 ;
        RECT 1690.200 54.050 1690.340 1086.990 ;
        RECT 1690.140 53.730 1690.400 54.050 ;
        RECT 2429.360 53.730 2429.620 54.050 ;
        RECT 2429.420 2.710 2429.560 53.730 ;
        RECT 2429.360 2.390 2429.620 2.710 ;
        RECT 2434.880 2.390 2435.140 2.710 ;
        RECT 2434.940 2.000 2435.080 2.390 ;
        RECT 2434.730 -4.000 2435.290 2.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1691.490 1088.580 1691.810 1088.640 ;
        RECT 1697.010 1088.580 1697.330 1088.640 ;
        RECT 1691.490 1088.440 1697.330 1088.580 ;
        RECT 1691.490 1088.380 1691.810 1088.440 ;
        RECT 1697.010 1088.380 1697.330 1088.440 ;
        RECT 1697.010 53.620 1697.330 53.680 ;
        RECT 2449.570 53.620 2449.890 53.680 ;
        RECT 1697.010 53.480 2449.890 53.620 ;
        RECT 1697.010 53.420 1697.330 53.480 ;
        RECT 2449.570 53.420 2449.890 53.480 ;
        RECT 2449.570 2.620 2449.890 2.680 ;
        RECT 2452.790 2.620 2453.110 2.680 ;
        RECT 2449.570 2.480 2453.110 2.620 ;
        RECT 2449.570 2.420 2449.890 2.480 ;
        RECT 2452.790 2.420 2453.110 2.480 ;
      LAYER via ;
        RECT 1691.520 1088.380 1691.780 1088.640 ;
        RECT 1697.040 1088.380 1697.300 1088.640 ;
        RECT 1697.040 53.420 1697.300 53.680 ;
        RECT 2449.600 53.420 2449.860 53.680 ;
        RECT 2449.600 2.420 2449.860 2.680 ;
        RECT 2452.820 2.420 2453.080 2.680 ;
      LAYER met2 ;
        RECT 1691.430 1100.580 1691.710 1104.000 ;
        RECT 1691.430 1100.000 1691.720 1100.580 ;
        RECT 1691.580 1088.670 1691.720 1100.000 ;
        RECT 1691.520 1088.350 1691.780 1088.670 ;
        RECT 1697.040 1088.350 1697.300 1088.670 ;
        RECT 1697.100 53.710 1697.240 1088.350 ;
        RECT 1697.040 53.390 1697.300 53.710 ;
        RECT 2449.600 53.390 2449.860 53.710 ;
        RECT 2449.660 2.710 2449.800 53.390 ;
        RECT 2449.600 2.390 2449.860 2.710 ;
        RECT 2452.820 2.390 2453.080 2.710 ;
        RECT 2452.880 2.000 2453.020 2.390 ;
        RECT 2452.670 -4.000 2453.230 2.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1697.930 1083.820 1698.250 1083.880 ;
        RECT 1703.910 1083.820 1704.230 1083.880 ;
        RECT 1697.930 1083.680 1704.230 1083.820 ;
        RECT 1697.930 1083.620 1698.250 1083.680 ;
        RECT 1703.910 1083.620 1704.230 1083.680 ;
        RECT 1703.910 53.280 1704.230 53.340 ;
        RECT 2470.730 53.280 2471.050 53.340 ;
        RECT 1703.910 53.140 2471.050 53.280 ;
        RECT 1703.910 53.080 1704.230 53.140 ;
        RECT 2470.730 53.080 2471.050 53.140 ;
      LAYER via ;
        RECT 1697.960 1083.620 1698.220 1083.880 ;
        RECT 1703.940 1083.620 1704.200 1083.880 ;
        RECT 1703.940 53.080 1704.200 53.340 ;
        RECT 2470.760 53.080 2471.020 53.340 ;
      LAYER met2 ;
        RECT 1697.870 1100.580 1698.150 1104.000 ;
        RECT 1697.870 1100.000 1698.160 1100.580 ;
        RECT 1698.020 1083.910 1698.160 1100.000 ;
        RECT 1697.960 1083.590 1698.220 1083.910 ;
        RECT 1703.940 1083.590 1704.200 1083.910 ;
        RECT 1704.000 53.370 1704.140 1083.590 ;
        RECT 1703.940 53.050 1704.200 53.370 ;
        RECT 2470.760 53.050 2471.020 53.370 ;
        RECT 2470.820 2.000 2470.960 53.050 ;
        RECT 2470.610 -4.000 2471.170 2.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1703.450 52.940 1703.770 53.000 ;
        RECT 2484.070 52.940 2484.390 53.000 ;
        RECT 1703.450 52.800 2484.390 52.940 ;
        RECT 1703.450 52.740 1703.770 52.800 ;
        RECT 2484.070 52.740 2484.390 52.800 ;
        RECT 2484.070 2.620 2484.390 2.680 ;
        RECT 2488.670 2.620 2488.990 2.680 ;
        RECT 2484.070 2.480 2488.990 2.620 ;
        RECT 2484.070 2.420 2484.390 2.480 ;
        RECT 2488.670 2.420 2488.990 2.480 ;
      LAYER via ;
        RECT 1703.480 52.740 1703.740 53.000 ;
        RECT 2484.100 52.740 2484.360 53.000 ;
        RECT 2484.100 2.420 2484.360 2.680 ;
        RECT 2488.700 2.420 2488.960 2.680 ;
      LAYER met2 ;
        RECT 1703.850 1100.650 1704.130 1104.000 ;
        RECT 1703.540 1100.510 1704.130 1100.650 ;
        RECT 1703.540 53.030 1703.680 1100.510 ;
        RECT 1703.850 1100.000 1704.130 1100.510 ;
        RECT 1703.480 52.710 1703.740 53.030 ;
        RECT 2484.100 52.710 2484.360 53.030 ;
        RECT 2484.160 2.710 2484.300 52.710 ;
        RECT 2484.100 2.390 2484.360 2.710 ;
        RECT 2488.700 2.390 2488.960 2.710 ;
        RECT 2488.760 2.000 2488.900 2.390 ;
        RECT 2488.550 -4.000 2489.110 2.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1710.810 52.600 1711.130 52.660 ;
        RECT 2504.770 52.600 2505.090 52.660 ;
        RECT 1710.810 52.460 2505.090 52.600 ;
        RECT 1710.810 52.400 1711.130 52.460 ;
        RECT 2504.770 52.400 2505.090 52.460 ;
      LAYER via ;
        RECT 1710.840 52.400 1711.100 52.660 ;
        RECT 2504.800 52.400 2505.060 52.660 ;
      LAYER met2 ;
        RECT 1709.830 1100.650 1710.110 1104.000 ;
        RECT 1709.830 1100.510 1711.040 1100.650 ;
        RECT 1709.830 1100.000 1710.110 1100.510 ;
        RECT 1710.900 52.690 1711.040 1100.510 ;
        RECT 1710.840 52.370 1711.100 52.690 ;
        RECT 2504.800 52.370 2505.060 52.690 ;
        RECT 2504.860 16.730 2505.000 52.370 ;
        RECT 2504.860 16.590 2506.380 16.730 ;
        RECT 2506.240 2.000 2506.380 16.590 ;
        RECT 2506.030 -4.000 2506.590 2.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1717.710 52.260 1718.030 52.320 ;
        RECT 2518.570 52.260 2518.890 52.320 ;
        RECT 1717.710 52.120 2518.890 52.260 ;
        RECT 1717.710 52.060 1718.030 52.120 ;
        RECT 2518.570 52.060 2518.890 52.120 ;
      LAYER via ;
        RECT 1717.740 52.060 1718.000 52.320 ;
        RECT 2518.600 52.060 2518.860 52.320 ;
      LAYER met2 ;
        RECT 1716.270 1100.650 1716.550 1104.000 ;
        RECT 1716.270 1100.510 1717.940 1100.650 ;
        RECT 1716.270 1100.000 1716.550 1100.510 ;
        RECT 1717.800 52.350 1717.940 1100.510 ;
        RECT 1717.740 52.030 1718.000 52.350 ;
        RECT 2518.600 52.030 2518.860 52.350 ;
        RECT 2518.660 16.730 2518.800 52.030 ;
        RECT 2518.660 16.590 2524.320 16.730 ;
        RECT 2524.180 2.000 2524.320 16.590 ;
        RECT 2523.970 -4.000 2524.530 2.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1724.150 51.920 1724.470 51.980 ;
        RECT 2539.270 51.920 2539.590 51.980 ;
        RECT 1724.150 51.780 2539.590 51.920 ;
        RECT 1724.150 51.720 1724.470 51.780 ;
        RECT 2539.270 51.720 2539.590 51.780 ;
      LAYER via ;
        RECT 1724.180 51.720 1724.440 51.980 ;
        RECT 2539.300 51.720 2539.560 51.980 ;
      LAYER met2 ;
        RECT 1722.250 1100.650 1722.530 1104.000 ;
        RECT 1722.250 1100.510 1723.920 1100.650 ;
        RECT 1722.250 1100.000 1722.530 1100.510 ;
        RECT 1723.780 1088.410 1723.920 1100.510 ;
        RECT 1723.780 1088.270 1724.380 1088.410 ;
        RECT 1724.240 52.010 1724.380 1088.270 ;
        RECT 1724.180 51.690 1724.440 52.010 ;
        RECT 2539.300 51.690 2539.560 52.010 ;
        RECT 2539.360 16.730 2539.500 51.690 ;
        RECT 2539.360 16.590 2542.260 16.730 ;
        RECT 2542.120 2.000 2542.260 16.590 ;
        RECT 2541.910 -4.000 2542.470 2.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1728.290 1089.260 1728.610 1089.320 ;
        RECT 1731.510 1089.260 1731.830 1089.320 ;
        RECT 1728.290 1089.120 1731.830 1089.260 ;
        RECT 1728.290 1089.060 1728.610 1089.120 ;
        RECT 1731.510 1089.060 1731.830 1089.120 ;
        RECT 1731.510 20.980 1731.830 21.040 ;
        RECT 2559.970 20.980 2560.290 21.040 ;
        RECT 1731.510 20.840 2560.290 20.980 ;
        RECT 1731.510 20.780 1731.830 20.840 ;
        RECT 2559.970 20.780 2560.290 20.840 ;
      LAYER via ;
        RECT 1728.320 1089.060 1728.580 1089.320 ;
        RECT 1731.540 1089.060 1731.800 1089.320 ;
        RECT 1731.540 20.780 1731.800 21.040 ;
        RECT 2560.000 20.780 2560.260 21.040 ;
      LAYER met2 ;
        RECT 1728.230 1100.580 1728.510 1104.000 ;
        RECT 1728.230 1100.000 1728.520 1100.580 ;
        RECT 1728.380 1089.350 1728.520 1100.000 ;
        RECT 1728.320 1089.030 1728.580 1089.350 ;
        RECT 1731.540 1089.030 1731.800 1089.350 ;
        RECT 1731.600 21.070 1731.740 1089.030 ;
        RECT 1731.540 20.750 1731.800 21.070 ;
        RECT 2560.000 20.750 2560.260 21.070 ;
        RECT 2560.060 2.000 2560.200 20.750 ;
        RECT 2559.850 -4.000 2560.410 2.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1734.730 1052.200 1735.050 1052.260 ;
        RECT 1738.410 1052.200 1738.730 1052.260 ;
        RECT 1734.730 1052.060 1738.730 1052.200 ;
        RECT 1734.730 1052.000 1735.050 1052.060 ;
        RECT 1738.410 1052.000 1738.730 1052.060 ;
        RECT 1738.410 21.320 1738.730 21.380 ;
        RECT 2577.910 21.320 2578.230 21.380 ;
        RECT 1738.410 21.180 2578.230 21.320 ;
        RECT 1738.410 21.120 1738.730 21.180 ;
        RECT 2577.910 21.120 2578.230 21.180 ;
      LAYER via ;
        RECT 1734.760 1052.000 1735.020 1052.260 ;
        RECT 1738.440 1052.000 1738.700 1052.260 ;
        RECT 1738.440 21.120 1738.700 21.380 ;
        RECT 2577.940 21.120 2578.200 21.380 ;
      LAYER met2 ;
        RECT 1734.670 1100.580 1734.950 1104.000 ;
        RECT 1734.670 1100.000 1734.960 1100.580 ;
        RECT 1734.820 1052.290 1734.960 1100.000 ;
        RECT 1734.760 1051.970 1735.020 1052.290 ;
        RECT 1738.440 1051.970 1738.700 1052.290 ;
        RECT 1738.500 21.410 1738.640 1051.970 ;
        RECT 1738.440 21.090 1738.700 21.410 ;
        RECT 2577.940 21.090 2578.200 21.410 ;
        RECT 2578.000 2.000 2578.140 21.090 ;
        RECT 2577.790 -4.000 2578.350 2.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1127.145 813.365 1127.315 862.495 ;
        RECT 1128.065 751.485 1128.235 793.475 ;
        RECT 1126.685 476.085 1126.855 498.355 ;
      LAYER mcon ;
        RECT 1127.145 862.325 1127.315 862.495 ;
        RECT 1128.065 793.305 1128.235 793.475 ;
        RECT 1126.685 498.185 1126.855 498.355 ;
      LAYER met1 ;
        RECT 1125.690 1048.800 1126.010 1048.860 ;
        RECT 1127.070 1048.800 1127.390 1048.860 ;
        RECT 1125.690 1048.660 1127.390 1048.800 ;
        RECT 1125.690 1048.600 1126.010 1048.660 ;
        RECT 1127.070 1048.600 1127.390 1048.660 ;
        RECT 1126.150 952.240 1126.470 952.300 ;
        RECT 1127.070 952.240 1127.390 952.300 ;
        RECT 1126.150 952.100 1127.390 952.240 ;
        RECT 1126.150 952.040 1126.470 952.100 ;
        RECT 1127.070 952.040 1127.390 952.100 ;
        RECT 1127.070 862.480 1127.390 862.540 ;
        RECT 1126.875 862.340 1127.390 862.480 ;
        RECT 1127.070 862.280 1127.390 862.340 ;
        RECT 1127.070 813.520 1127.390 813.580 ;
        RECT 1126.875 813.380 1127.390 813.520 ;
        RECT 1127.070 813.320 1127.390 813.380 ;
        RECT 1127.070 800.260 1127.390 800.320 ;
        RECT 1127.990 800.260 1128.310 800.320 ;
        RECT 1127.070 800.120 1128.310 800.260 ;
        RECT 1127.070 800.060 1127.390 800.120 ;
        RECT 1127.990 800.060 1128.310 800.120 ;
        RECT 1127.990 793.460 1128.310 793.520 ;
        RECT 1127.795 793.320 1128.310 793.460 ;
        RECT 1127.990 793.260 1128.310 793.320 ;
        RECT 1127.990 751.640 1128.310 751.700 ;
        RECT 1127.795 751.500 1128.310 751.640 ;
        RECT 1127.990 751.440 1128.310 751.500 ;
        RECT 1126.150 704.040 1126.470 704.100 ;
        RECT 1127.990 704.040 1128.310 704.100 ;
        RECT 1126.150 703.900 1128.310 704.040 ;
        RECT 1126.150 703.840 1126.470 703.900 ;
        RECT 1127.990 703.840 1128.310 703.900 ;
        RECT 1126.610 669.020 1126.930 669.080 ;
        RECT 1127.530 669.020 1127.850 669.080 ;
        RECT 1126.610 668.880 1127.850 669.020 ;
        RECT 1126.610 668.820 1126.930 668.880 ;
        RECT 1127.530 668.820 1127.850 668.880 ;
        RECT 1126.150 613.940 1126.470 614.000 ;
        RECT 1126.610 613.940 1126.930 614.000 ;
        RECT 1126.150 613.800 1126.930 613.940 ;
        RECT 1126.150 613.740 1126.470 613.800 ;
        RECT 1126.610 613.740 1126.930 613.800 ;
        RECT 1126.610 498.340 1126.930 498.400 ;
        RECT 1126.415 498.200 1126.930 498.340 ;
        RECT 1126.610 498.140 1126.930 498.200 ;
        RECT 1126.610 476.240 1126.930 476.300 ;
        RECT 1126.415 476.100 1126.930 476.240 ;
        RECT 1126.610 476.040 1126.930 476.100 ;
        RECT 1126.150 434.760 1126.470 434.820 ;
        RECT 1126.610 434.760 1126.930 434.820 ;
        RECT 1126.150 434.620 1126.930 434.760 ;
        RECT 1126.150 434.560 1126.470 434.620 ;
        RECT 1126.610 434.560 1126.930 434.620 ;
        RECT 1126.150 338.200 1126.470 338.260 ;
        RECT 1126.610 338.200 1126.930 338.260 ;
        RECT 1126.150 338.060 1126.930 338.200 ;
        RECT 1126.150 338.000 1126.470 338.060 ;
        RECT 1126.610 338.000 1126.930 338.060 ;
        RECT 1126.150 282.780 1126.470 282.840 ;
        RECT 1127.530 282.780 1127.850 282.840 ;
        RECT 1126.150 282.640 1127.850 282.780 ;
        RECT 1126.150 282.580 1126.470 282.640 ;
        RECT 1127.530 282.580 1127.850 282.640 ;
        RECT 1126.150 186.560 1126.470 186.620 ;
        RECT 1127.530 186.560 1127.850 186.620 ;
        RECT 1126.150 186.420 1127.850 186.560 ;
        RECT 1126.150 186.360 1126.470 186.420 ;
        RECT 1127.530 186.360 1127.850 186.420 ;
        RECT 811.510 43.080 811.830 43.140 ;
        RECT 1126.150 43.080 1126.470 43.140 ;
        RECT 811.510 42.940 1126.470 43.080 ;
        RECT 811.510 42.880 811.830 42.940 ;
        RECT 1126.150 42.880 1126.470 42.940 ;
      LAYER via ;
        RECT 1125.720 1048.600 1125.980 1048.860 ;
        RECT 1127.100 1048.600 1127.360 1048.860 ;
        RECT 1126.180 952.040 1126.440 952.300 ;
        RECT 1127.100 952.040 1127.360 952.300 ;
        RECT 1127.100 862.280 1127.360 862.540 ;
        RECT 1127.100 813.320 1127.360 813.580 ;
        RECT 1127.100 800.060 1127.360 800.320 ;
        RECT 1128.020 800.060 1128.280 800.320 ;
        RECT 1128.020 793.260 1128.280 793.520 ;
        RECT 1128.020 751.440 1128.280 751.700 ;
        RECT 1126.180 703.840 1126.440 704.100 ;
        RECT 1128.020 703.840 1128.280 704.100 ;
        RECT 1126.640 668.820 1126.900 669.080 ;
        RECT 1127.560 668.820 1127.820 669.080 ;
        RECT 1126.180 613.740 1126.440 614.000 ;
        RECT 1126.640 613.740 1126.900 614.000 ;
        RECT 1126.640 498.140 1126.900 498.400 ;
        RECT 1126.640 476.040 1126.900 476.300 ;
        RECT 1126.180 434.560 1126.440 434.820 ;
        RECT 1126.640 434.560 1126.900 434.820 ;
        RECT 1126.180 338.000 1126.440 338.260 ;
        RECT 1126.640 338.000 1126.900 338.260 ;
        RECT 1126.180 282.580 1126.440 282.840 ;
        RECT 1127.560 282.580 1127.820 282.840 ;
        RECT 1126.180 186.360 1126.440 186.620 ;
        RECT 1127.560 186.360 1127.820 186.620 ;
        RECT 811.540 42.880 811.800 43.140 ;
        RECT 1126.180 42.880 1126.440 43.140 ;
      LAYER met2 ;
        RECT 1128.390 1100.650 1128.670 1104.000 ;
        RECT 1127.620 1100.510 1128.670 1100.650 ;
        RECT 1127.620 1055.770 1127.760 1100.510 ;
        RECT 1128.390 1100.000 1128.670 1100.510 ;
        RECT 1127.160 1055.630 1127.760 1055.770 ;
        RECT 1127.160 1048.890 1127.300 1055.630 ;
        RECT 1125.720 1048.570 1125.980 1048.890 ;
        RECT 1127.100 1048.570 1127.360 1048.890 ;
        RECT 1125.780 1000.805 1125.920 1048.570 ;
        RECT 1125.710 1000.435 1125.990 1000.805 ;
        RECT 1126.630 1000.435 1126.910 1000.805 ;
        RECT 1126.700 952.410 1126.840 1000.435 ;
        RECT 1126.700 952.330 1127.300 952.410 ;
        RECT 1126.180 952.010 1126.440 952.330 ;
        RECT 1126.700 952.270 1127.360 952.330 ;
        RECT 1127.100 952.010 1127.360 952.270 ;
        RECT 1126.240 904.245 1126.380 952.010 ;
        RECT 1127.160 951.855 1127.300 952.010 ;
        RECT 1126.170 903.875 1126.450 904.245 ;
        RECT 1127.550 903.875 1127.830 904.245 ;
        RECT 1127.620 884.410 1127.760 903.875 ;
        RECT 1127.160 884.270 1127.760 884.410 ;
        RECT 1127.160 862.570 1127.300 884.270 ;
        RECT 1127.100 862.250 1127.360 862.570 ;
        RECT 1127.100 813.290 1127.360 813.610 ;
        RECT 1127.160 800.350 1127.300 813.290 ;
        RECT 1127.100 800.030 1127.360 800.350 ;
        RECT 1128.020 800.030 1128.280 800.350 ;
        RECT 1128.080 793.550 1128.220 800.030 ;
        RECT 1128.020 793.230 1128.280 793.550 ;
        RECT 1128.020 751.410 1128.280 751.730 ;
        RECT 1128.080 704.130 1128.220 751.410 ;
        RECT 1126.180 703.810 1126.440 704.130 ;
        RECT 1128.020 703.810 1128.280 704.130 ;
        RECT 1126.240 703.530 1126.380 703.810 ;
        RECT 1126.630 703.530 1126.910 703.645 ;
        RECT 1126.240 703.390 1126.910 703.530 ;
        RECT 1126.630 703.275 1126.910 703.390 ;
        RECT 1127.550 703.275 1127.830 703.645 ;
        RECT 1127.620 669.110 1127.760 703.275 ;
        RECT 1126.640 668.790 1126.900 669.110 ;
        RECT 1127.560 668.790 1127.820 669.110 ;
        RECT 1126.700 614.030 1126.840 668.790 ;
        RECT 1126.180 613.710 1126.440 614.030 ;
        RECT 1126.640 613.710 1126.900 614.030 ;
        RECT 1126.240 589.290 1126.380 613.710 ;
        RECT 1126.240 589.150 1126.840 589.290 ;
        RECT 1126.700 498.430 1126.840 589.150 ;
        RECT 1126.640 498.110 1126.900 498.430 ;
        RECT 1126.640 476.010 1126.900 476.330 ;
        RECT 1126.700 434.850 1126.840 476.010 ;
        RECT 1126.180 434.530 1126.440 434.850 ;
        RECT 1126.640 434.530 1126.900 434.850 ;
        RECT 1126.240 403.650 1126.380 434.530 ;
        RECT 1126.240 403.510 1127.300 403.650 ;
        RECT 1127.160 385.970 1127.300 403.510 ;
        RECT 1126.700 385.830 1127.300 385.970 ;
        RECT 1126.700 338.290 1126.840 385.830 ;
        RECT 1126.180 337.970 1126.440 338.290 ;
        RECT 1126.640 337.970 1126.900 338.290 ;
        RECT 1126.240 282.870 1126.380 337.970 ;
        RECT 1126.180 282.550 1126.440 282.870 ;
        RECT 1127.560 282.550 1127.820 282.870 ;
        RECT 1127.620 186.650 1127.760 282.550 ;
        RECT 1126.180 186.330 1126.440 186.650 ;
        RECT 1127.560 186.330 1127.820 186.650 ;
        RECT 1126.240 43.170 1126.380 186.330 ;
        RECT 811.540 42.850 811.800 43.170 ;
        RECT 1126.180 42.850 1126.440 43.170 ;
        RECT 811.600 2.000 811.740 42.850 ;
        RECT 811.390 -4.000 811.950 2.000 ;
      LAYER via2 ;
        RECT 1125.710 1000.480 1125.990 1000.760 ;
        RECT 1126.630 1000.480 1126.910 1000.760 ;
        RECT 1126.170 903.920 1126.450 904.200 ;
        RECT 1127.550 903.920 1127.830 904.200 ;
        RECT 1126.630 703.320 1126.910 703.600 ;
        RECT 1127.550 703.320 1127.830 703.600 ;
      LAYER met3 ;
        RECT 1125.685 1000.770 1126.015 1000.785 ;
        RECT 1126.605 1000.770 1126.935 1000.785 ;
        RECT 1125.685 1000.470 1126.935 1000.770 ;
        RECT 1125.685 1000.455 1126.015 1000.470 ;
        RECT 1126.605 1000.455 1126.935 1000.470 ;
        RECT 1126.145 904.210 1126.475 904.225 ;
        RECT 1127.525 904.210 1127.855 904.225 ;
        RECT 1126.145 903.910 1127.855 904.210 ;
        RECT 1126.145 903.895 1126.475 903.910 ;
        RECT 1127.525 903.895 1127.855 903.910 ;
        RECT 1126.605 703.610 1126.935 703.625 ;
        RECT 1127.525 703.610 1127.855 703.625 ;
        RECT 1126.605 703.310 1127.855 703.610 ;
        RECT 1126.605 703.295 1126.935 703.310 ;
        RECT 1127.525 703.295 1127.855 703.310 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1740.710 1089.260 1741.030 1089.320 ;
        RECT 1745.310 1089.260 1745.630 1089.320 ;
        RECT 1740.710 1089.120 1745.630 1089.260 ;
        RECT 1740.710 1089.060 1741.030 1089.120 ;
        RECT 1745.310 1089.060 1745.630 1089.120 ;
        RECT 1744.850 21.660 1745.170 21.720 ;
        RECT 2595.390 21.660 2595.710 21.720 ;
        RECT 1744.850 21.520 2595.710 21.660 ;
        RECT 1744.850 21.460 1745.170 21.520 ;
        RECT 2595.390 21.460 2595.710 21.520 ;
      LAYER via ;
        RECT 1740.740 1089.060 1741.000 1089.320 ;
        RECT 1745.340 1089.060 1745.600 1089.320 ;
        RECT 1744.880 21.460 1745.140 21.720 ;
        RECT 2595.420 21.460 2595.680 21.720 ;
      LAYER met2 ;
        RECT 1740.650 1100.580 1740.930 1104.000 ;
        RECT 1740.650 1100.000 1740.940 1100.580 ;
        RECT 1740.800 1089.350 1740.940 1100.000 ;
        RECT 1740.740 1089.030 1741.000 1089.350 ;
        RECT 1745.340 1089.030 1745.600 1089.350 ;
        RECT 1745.400 41.210 1745.540 1089.030 ;
        RECT 1744.940 41.070 1745.540 41.210 ;
        RECT 1744.940 21.750 1745.080 41.070 ;
        RECT 1744.880 21.430 1745.140 21.750 ;
        RECT 2595.420 21.430 2595.680 21.750 ;
        RECT 2595.480 2.000 2595.620 21.430 ;
        RECT 2595.270 -4.000 2595.830 2.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1746.690 1089.940 1747.010 1090.000 ;
        RECT 1752.210 1089.940 1752.530 1090.000 ;
        RECT 1746.690 1089.800 1752.530 1089.940 ;
        RECT 1746.690 1089.740 1747.010 1089.800 ;
        RECT 1752.210 1089.740 1752.530 1089.800 ;
        RECT 1752.210 22.000 1752.530 22.060 ;
        RECT 2613.330 22.000 2613.650 22.060 ;
        RECT 1752.210 21.860 2613.650 22.000 ;
        RECT 1752.210 21.800 1752.530 21.860 ;
        RECT 2613.330 21.800 2613.650 21.860 ;
      LAYER via ;
        RECT 1746.720 1089.740 1746.980 1090.000 ;
        RECT 1752.240 1089.740 1752.500 1090.000 ;
        RECT 1752.240 21.800 1752.500 22.060 ;
        RECT 2613.360 21.800 2613.620 22.060 ;
      LAYER met2 ;
        RECT 1746.630 1100.580 1746.910 1104.000 ;
        RECT 1746.630 1100.000 1746.920 1100.580 ;
        RECT 1746.780 1090.030 1746.920 1100.000 ;
        RECT 1746.720 1089.710 1746.980 1090.030 ;
        RECT 1752.240 1089.710 1752.500 1090.030 ;
        RECT 1752.300 22.090 1752.440 1089.710 ;
        RECT 1752.240 21.770 1752.500 22.090 ;
        RECT 2613.360 21.770 2613.620 22.090 ;
        RECT 2613.420 2.000 2613.560 21.770 ;
        RECT 2613.210 -4.000 2613.770 2.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1753.130 1088.920 1753.450 1088.980 ;
        RECT 1759.110 1088.920 1759.430 1088.980 ;
        RECT 1753.130 1088.780 1759.430 1088.920 ;
        RECT 1753.130 1088.720 1753.450 1088.780 ;
        RECT 1759.110 1088.720 1759.430 1088.780 ;
        RECT 1759.110 22.340 1759.430 22.400 ;
        RECT 2631.270 22.340 2631.590 22.400 ;
        RECT 1759.110 22.200 2631.590 22.340 ;
        RECT 1759.110 22.140 1759.430 22.200 ;
        RECT 2631.270 22.140 2631.590 22.200 ;
      LAYER via ;
        RECT 1753.160 1088.720 1753.420 1088.980 ;
        RECT 1759.140 1088.720 1759.400 1088.980 ;
        RECT 1759.140 22.140 1759.400 22.400 ;
        RECT 2631.300 22.140 2631.560 22.400 ;
      LAYER met2 ;
        RECT 1753.070 1100.580 1753.350 1104.000 ;
        RECT 1753.070 1100.000 1753.360 1100.580 ;
        RECT 1753.220 1089.010 1753.360 1100.000 ;
        RECT 1753.160 1088.690 1753.420 1089.010 ;
        RECT 1759.140 1088.690 1759.400 1089.010 ;
        RECT 1759.200 22.430 1759.340 1088.690 ;
        RECT 1759.140 22.110 1759.400 22.430 ;
        RECT 2631.300 22.110 2631.560 22.430 ;
        RECT 2631.360 2.000 2631.500 22.110 ;
        RECT 2631.150 -4.000 2631.710 2.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1758.650 22.680 1758.970 22.740 ;
        RECT 2649.210 22.680 2649.530 22.740 ;
        RECT 1758.650 22.540 2649.530 22.680 ;
        RECT 1758.650 22.480 1758.970 22.540 ;
        RECT 2649.210 22.480 2649.530 22.540 ;
      LAYER via ;
        RECT 1758.680 22.480 1758.940 22.740 ;
        RECT 2649.240 22.480 2649.500 22.740 ;
      LAYER met2 ;
        RECT 1759.050 1100.650 1759.330 1104.000 ;
        RECT 1758.740 1100.510 1759.330 1100.650 ;
        RECT 1758.740 22.770 1758.880 1100.510 ;
        RECT 1759.050 1100.000 1759.330 1100.510 ;
        RECT 1758.680 22.450 1758.940 22.770 ;
        RECT 2649.240 22.450 2649.500 22.770 ;
        RECT 2649.300 2.000 2649.440 22.450 ;
        RECT 2649.090 -4.000 2649.650 2.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1766.010 23.020 1766.330 23.080 ;
        RECT 2667.150 23.020 2667.470 23.080 ;
        RECT 1766.010 22.880 2667.470 23.020 ;
        RECT 1766.010 22.820 1766.330 22.880 ;
        RECT 2667.150 22.820 2667.470 22.880 ;
      LAYER via ;
        RECT 1766.040 22.820 1766.300 23.080 ;
        RECT 2667.180 22.820 2667.440 23.080 ;
      LAYER met2 ;
        RECT 1765.030 1100.650 1765.310 1104.000 ;
        RECT 1765.030 1100.510 1766.240 1100.650 ;
        RECT 1765.030 1100.000 1765.310 1100.510 ;
        RECT 1766.100 23.110 1766.240 1100.510 ;
        RECT 1766.040 22.790 1766.300 23.110 ;
        RECT 2667.180 22.790 2667.440 23.110 ;
        RECT 2667.240 2.000 2667.380 22.790 ;
        RECT 2667.030 -4.000 2667.590 2.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1772.910 23.360 1773.230 23.420 ;
        RECT 2684.630 23.360 2684.950 23.420 ;
        RECT 1772.910 23.220 2684.950 23.360 ;
        RECT 1772.910 23.160 1773.230 23.220 ;
        RECT 2684.630 23.160 2684.950 23.220 ;
      LAYER via ;
        RECT 1772.940 23.160 1773.200 23.420 ;
        RECT 2684.660 23.160 2684.920 23.420 ;
      LAYER met2 ;
        RECT 1771.010 1100.650 1771.290 1104.000 ;
        RECT 1771.010 1100.510 1773.140 1100.650 ;
        RECT 1771.010 1100.000 1771.290 1100.510 ;
        RECT 1773.000 23.450 1773.140 1100.510 ;
        RECT 1772.940 23.130 1773.200 23.450 ;
        RECT 2684.660 23.130 2684.920 23.450 ;
        RECT 2684.720 2.000 2684.860 23.130 ;
        RECT 2684.510 -4.000 2685.070 2.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1779.885 336.685 1780.055 379.355 ;
      LAYER mcon ;
        RECT 1779.885 379.185 1780.055 379.355 ;
      LAYER met1 ;
        RECT 1777.510 1088.580 1777.830 1088.640 ;
        RECT 1779.810 1088.580 1780.130 1088.640 ;
        RECT 1777.510 1088.440 1780.130 1088.580 ;
        RECT 1777.510 1088.380 1777.830 1088.440 ;
        RECT 1779.810 1088.380 1780.130 1088.440 ;
        RECT 1779.810 379.340 1780.130 379.400 ;
        RECT 1779.615 379.200 1780.130 379.340 ;
        RECT 1779.810 379.140 1780.130 379.200 ;
        RECT 1779.810 336.840 1780.130 336.900 ;
        RECT 1779.615 336.700 1780.130 336.840 ;
        RECT 1779.810 336.640 1780.130 336.700 ;
        RECT 1779.810 23.700 1780.130 23.760 ;
        RECT 2702.570 23.700 2702.890 23.760 ;
        RECT 1779.810 23.560 2702.890 23.700 ;
        RECT 1779.810 23.500 1780.130 23.560 ;
        RECT 2702.570 23.500 2702.890 23.560 ;
      LAYER via ;
        RECT 1777.540 1088.380 1777.800 1088.640 ;
        RECT 1779.840 1088.380 1780.100 1088.640 ;
        RECT 1779.840 379.140 1780.100 379.400 ;
        RECT 1779.840 336.640 1780.100 336.900 ;
        RECT 1779.840 23.500 1780.100 23.760 ;
        RECT 2702.600 23.500 2702.860 23.760 ;
      LAYER met2 ;
        RECT 1777.450 1100.580 1777.730 1104.000 ;
        RECT 1777.450 1100.000 1777.740 1100.580 ;
        RECT 1777.600 1088.670 1777.740 1100.000 ;
        RECT 1777.540 1088.350 1777.800 1088.670 ;
        RECT 1779.840 1088.350 1780.100 1088.670 ;
        RECT 1779.900 379.430 1780.040 1088.350 ;
        RECT 1779.840 379.110 1780.100 379.430 ;
        RECT 1779.840 336.610 1780.100 336.930 ;
        RECT 1779.900 23.790 1780.040 336.610 ;
        RECT 1779.840 23.470 1780.100 23.790 ;
        RECT 2702.600 23.470 2702.860 23.790 ;
        RECT 2702.660 2.000 2702.800 23.470 ;
        RECT 2702.450 -4.000 2703.010 2.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1783.490 1088.920 1783.810 1088.980 ;
        RECT 1786.710 1088.920 1787.030 1088.980 ;
        RECT 1783.490 1088.780 1787.030 1088.920 ;
        RECT 1783.490 1088.720 1783.810 1088.780 ;
        RECT 1786.710 1088.720 1787.030 1088.780 ;
        RECT 1786.710 27.440 1787.030 27.500 ;
        RECT 2720.510 27.440 2720.830 27.500 ;
        RECT 1786.710 27.300 2720.830 27.440 ;
        RECT 1786.710 27.240 1787.030 27.300 ;
        RECT 2720.510 27.240 2720.830 27.300 ;
      LAYER via ;
        RECT 1783.520 1088.720 1783.780 1088.980 ;
        RECT 1786.740 1088.720 1787.000 1088.980 ;
        RECT 1786.740 27.240 1787.000 27.500 ;
        RECT 2720.540 27.240 2720.800 27.500 ;
      LAYER met2 ;
        RECT 1783.430 1100.580 1783.710 1104.000 ;
        RECT 1783.430 1100.000 1783.720 1100.580 ;
        RECT 1783.580 1089.010 1783.720 1100.000 ;
        RECT 1783.520 1088.690 1783.780 1089.010 ;
        RECT 1786.740 1088.690 1787.000 1089.010 ;
        RECT 1786.800 27.530 1786.940 1088.690 ;
        RECT 1786.740 27.210 1787.000 27.530 ;
        RECT 2720.540 27.210 2720.800 27.530 ;
        RECT 2720.600 2.000 2720.740 27.210 ;
        RECT 2720.390 -4.000 2720.950 2.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1789.470 1088.920 1789.790 1088.980 ;
        RECT 1793.610 1088.920 1793.930 1088.980 ;
        RECT 1789.470 1088.780 1793.930 1088.920 ;
        RECT 1789.470 1088.720 1789.790 1088.780 ;
        RECT 1793.610 1088.720 1793.930 1088.780 ;
        RECT 1793.610 27.100 1793.930 27.160 ;
        RECT 2738.450 27.100 2738.770 27.160 ;
        RECT 1793.610 26.960 2738.770 27.100 ;
        RECT 1793.610 26.900 1793.930 26.960 ;
        RECT 2738.450 26.900 2738.770 26.960 ;
      LAYER via ;
        RECT 1789.500 1088.720 1789.760 1088.980 ;
        RECT 1793.640 1088.720 1793.900 1088.980 ;
        RECT 1793.640 26.900 1793.900 27.160 ;
        RECT 2738.480 26.900 2738.740 27.160 ;
      LAYER met2 ;
        RECT 1789.410 1100.580 1789.690 1104.000 ;
        RECT 1789.410 1100.000 1789.700 1100.580 ;
        RECT 1789.560 1089.010 1789.700 1100.000 ;
        RECT 1789.500 1088.690 1789.760 1089.010 ;
        RECT 1793.640 1088.690 1793.900 1089.010 ;
        RECT 1793.700 27.190 1793.840 1088.690 ;
        RECT 1793.640 26.870 1793.900 27.190 ;
        RECT 2738.480 26.870 2738.740 27.190 ;
        RECT 2738.540 2.000 2738.680 26.870 ;
        RECT 2738.330 -4.000 2738.890 2.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1795.910 1088.580 1796.230 1088.640 ;
        RECT 1800.050 1088.580 1800.370 1088.640 ;
        RECT 1795.910 1088.440 1800.370 1088.580 ;
        RECT 1795.910 1088.380 1796.230 1088.440 ;
        RECT 1800.050 1088.380 1800.370 1088.440 ;
        RECT 1800.050 26.760 1800.370 26.820 ;
        RECT 2755.930 26.760 2756.250 26.820 ;
        RECT 1800.050 26.620 2756.250 26.760 ;
        RECT 1800.050 26.560 1800.370 26.620 ;
        RECT 2755.930 26.560 2756.250 26.620 ;
      LAYER via ;
        RECT 1795.940 1088.380 1796.200 1088.640 ;
        RECT 1800.080 1088.380 1800.340 1088.640 ;
        RECT 1800.080 26.560 1800.340 26.820 ;
        RECT 2755.960 26.560 2756.220 26.820 ;
      LAYER met2 ;
        RECT 1795.850 1100.580 1796.130 1104.000 ;
        RECT 1795.850 1100.000 1796.140 1100.580 ;
        RECT 1796.000 1088.670 1796.140 1100.000 ;
        RECT 1795.940 1088.350 1796.200 1088.670 ;
        RECT 1800.080 1088.350 1800.340 1088.670 ;
        RECT 1800.140 26.850 1800.280 1088.350 ;
        RECT 1800.080 26.530 1800.340 26.850 ;
        RECT 2755.960 26.530 2756.220 26.850 ;
        RECT 2756.020 2.000 2756.160 26.530 ;
        RECT 2755.810 -4.000 2756.370 2.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 829.450 42.740 829.770 42.800 ;
        RECT 1133.050 42.740 1133.370 42.800 ;
        RECT 829.450 42.600 1133.370 42.740 ;
        RECT 829.450 42.540 829.770 42.600 ;
        RECT 1133.050 42.540 1133.370 42.600 ;
      LAYER via ;
        RECT 829.480 42.540 829.740 42.800 ;
        RECT 1133.080 42.540 1133.340 42.800 ;
      LAYER met2 ;
        RECT 1134.370 1100.650 1134.650 1104.000 ;
        RECT 1133.140 1100.510 1134.650 1100.650 ;
        RECT 1133.140 42.830 1133.280 1100.510 ;
        RECT 1134.370 1100.000 1134.650 1100.510 ;
        RECT 829.480 42.510 829.740 42.830 ;
        RECT 1133.080 42.510 1133.340 42.830 ;
        RECT 829.540 2.000 829.680 42.510 ;
        RECT 829.330 -4.000 829.890 2.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1801.890 1088.580 1802.210 1088.640 ;
        RECT 1807.410 1088.580 1807.730 1088.640 ;
        RECT 1801.890 1088.440 1807.730 1088.580 ;
        RECT 1801.890 1088.380 1802.210 1088.440 ;
        RECT 1807.410 1088.380 1807.730 1088.440 ;
        RECT 1807.410 26.420 1807.730 26.480 ;
        RECT 2773.870 26.420 2774.190 26.480 ;
        RECT 1807.410 26.280 2774.190 26.420 ;
        RECT 1807.410 26.220 1807.730 26.280 ;
        RECT 2773.870 26.220 2774.190 26.280 ;
      LAYER via ;
        RECT 1801.920 1088.380 1802.180 1088.640 ;
        RECT 1807.440 1088.380 1807.700 1088.640 ;
        RECT 1807.440 26.220 1807.700 26.480 ;
        RECT 2773.900 26.220 2774.160 26.480 ;
      LAYER met2 ;
        RECT 1801.830 1100.580 1802.110 1104.000 ;
        RECT 1801.830 1100.000 1802.120 1100.580 ;
        RECT 1801.980 1088.670 1802.120 1100.000 ;
        RECT 1801.920 1088.350 1802.180 1088.670 ;
        RECT 1807.440 1088.350 1807.700 1088.670 ;
        RECT 1807.500 26.510 1807.640 1088.350 ;
        RECT 1807.440 26.190 1807.700 26.510 ;
        RECT 2773.900 26.190 2774.160 26.510 ;
        RECT 2773.960 2.000 2774.100 26.190 ;
        RECT 2773.750 -4.000 2774.310 2.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1807.870 1088.920 1808.190 1088.980 ;
        RECT 1813.850 1088.920 1814.170 1088.980 ;
        RECT 1807.870 1088.780 1814.170 1088.920 ;
        RECT 1807.870 1088.720 1808.190 1088.780 ;
        RECT 1813.850 1088.720 1814.170 1088.780 ;
        RECT 1813.850 26.080 1814.170 26.140 ;
        RECT 2791.810 26.080 2792.130 26.140 ;
        RECT 1813.850 25.940 2792.130 26.080 ;
        RECT 1813.850 25.880 1814.170 25.940 ;
        RECT 2791.810 25.880 2792.130 25.940 ;
      LAYER via ;
        RECT 1807.900 1088.720 1808.160 1088.980 ;
        RECT 1813.880 1088.720 1814.140 1088.980 ;
        RECT 1813.880 25.880 1814.140 26.140 ;
        RECT 2791.840 25.880 2792.100 26.140 ;
      LAYER met2 ;
        RECT 1807.810 1100.580 1808.090 1104.000 ;
        RECT 1807.810 1100.000 1808.100 1100.580 ;
        RECT 1807.960 1089.010 1808.100 1100.000 ;
        RECT 1807.900 1088.690 1808.160 1089.010 ;
        RECT 1813.880 1088.690 1814.140 1089.010 ;
        RECT 1813.940 26.170 1814.080 1088.690 ;
        RECT 1813.880 25.850 1814.140 26.170 ;
        RECT 2791.840 25.850 2792.100 26.170 ;
        RECT 2791.900 2.000 2792.040 25.850 ;
        RECT 2791.690 -4.000 2792.250 2.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1813.390 25.740 1813.710 25.800 ;
        RECT 2809.750 25.740 2810.070 25.800 ;
        RECT 1813.390 25.600 2810.070 25.740 ;
        RECT 1813.390 25.540 1813.710 25.600 ;
        RECT 2809.750 25.540 2810.070 25.600 ;
      LAYER via ;
        RECT 1813.420 25.540 1813.680 25.800 ;
        RECT 2809.780 25.540 2810.040 25.800 ;
      LAYER met2 ;
        RECT 1814.250 1100.650 1814.530 1104.000 ;
        RECT 1813.480 1100.510 1814.530 1100.650 ;
        RECT 1813.480 25.830 1813.620 1100.510 ;
        RECT 1814.250 1100.000 1814.530 1100.510 ;
        RECT 1813.420 25.510 1813.680 25.830 ;
        RECT 2809.780 25.510 2810.040 25.830 ;
        RECT 2809.840 2.000 2809.980 25.510 ;
        RECT 2809.630 -4.000 2810.190 2.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1821.210 25.400 1821.530 25.460 ;
        RECT 2827.690 25.400 2828.010 25.460 ;
        RECT 1821.210 25.260 2828.010 25.400 ;
        RECT 1821.210 25.200 1821.530 25.260 ;
        RECT 2827.690 25.200 2828.010 25.260 ;
      LAYER via ;
        RECT 1821.240 25.200 1821.500 25.460 ;
        RECT 2827.720 25.200 2827.980 25.460 ;
      LAYER met2 ;
        RECT 1820.230 1100.650 1820.510 1104.000 ;
        RECT 1820.230 1100.510 1821.440 1100.650 ;
        RECT 1820.230 1100.000 1820.510 1100.510 ;
        RECT 1821.300 25.490 1821.440 1100.510 ;
        RECT 1821.240 25.170 1821.500 25.490 ;
        RECT 2827.720 25.170 2827.980 25.490 ;
        RECT 2827.780 2.000 2827.920 25.170 ;
        RECT 2827.570 -4.000 2828.130 2.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1827.650 25.060 1827.970 25.120 ;
        RECT 2845.170 25.060 2845.490 25.120 ;
        RECT 1827.650 24.920 2845.490 25.060 ;
        RECT 1827.650 24.860 1827.970 24.920 ;
        RECT 2845.170 24.860 2845.490 24.920 ;
      LAYER via ;
        RECT 1827.680 24.860 1827.940 25.120 ;
        RECT 2845.200 24.860 2845.460 25.120 ;
      LAYER met2 ;
        RECT 1826.210 1100.650 1826.490 1104.000 ;
        RECT 1826.210 1100.510 1827.880 1100.650 ;
        RECT 1826.210 1100.000 1826.490 1100.510 ;
        RECT 1827.740 25.150 1827.880 1100.510 ;
        RECT 1827.680 24.830 1827.940 25.150 ;
        RECT 2845.200 24.830 2845.460 25.150 ;
        RECT 2845.260 2.000 2845.400 24.830 ;
        RECT 2845.050 -4.000 2845.610 2.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1832.710 1088.580 1833.030 1088.640 ;
        RECT 1835.010 1088.580 1835.330 1088.640 ;
        RECT 1832.710 1088.440 1835.330 1088.580 ;
        RECT 1832.710 1088.380 1833.030 1088.440 ;
        RECT 1835.010 1088.380 1835.330 1088.440 ;
        RECT 1833.630 55.320 1833.950 55.380 ;
        RECT 1835.010 55.320 1835.330 55.380 ;
        RECT 1833.630 55.180 1835.330 55.320 ;
        RECT 1833.630 55.120 1833.950 55.180 ;
        RECT 1835.010 55.120 1835.330 55.180 ;
        RECT 1833.630 24.720 1833.950 24.780 ;
        RECT 2863.110 24.720 2863.430 24.780 ;
        RECT 1833.630 24.580 2863.430 24.720 ;
        RECT 1833.630 24.520 1833.950 24.580 ;
        RECT 2863.110 24.520 2863.430 24.580 ;
      LAYER via ;
        RECT 1832.740 1088.380 1833.000 1088.640 ;
        RECT 1835.040 1088.380 1835.300 1088.640 ;
        RECT 1833.660 55.120 1833.920 55.380 ;
        RECT 1835.040 55.120 1835.300 55.380 ;
        RECT 1833.660 24.520 1833.920 24.780 ;
        RECT 2863.140 24.520 2863.400 24.780 ;
      LAYER met2 ;
        RECT 1832.650 1100.580 1832.930 1104.000 ;
        RECT 1832.650 1100.000 1832.940 1100.580 ;
        RECT 1832.800 1088.670 1832.940 1100.000 ;
        RECT 1832.740 1088.350 1833.000 1088.670 ;
        RECT 1835.040 1088.350 1835.300 1088.670 ;
        RECT 1835.100 55.410 1835.240 1088.350 ;
        RECT 1833.660 55.090 1833.920 55.410 ;
        RECT 1835.040 55.090 1835.300 55.410 ;
        RECT 1833.720 24.810 1833.860 55.090 ;
        RECT 1833.660 24.490 1833.920 24.810 ;
        RECT 2863.140 24.490 2863.400 24.810 ;
        RECT 2863.200 2.000 2863.340 24.490 ;
        RECT 2862.990 -4.000 2863.550 2.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1838.690 1088.580 1839.010 1088.640 ;
        RECT 1841.450 1088.580 1841.770 1088.640 ;
        RECT 1838.690 1088.440 1841.770 1088.580 ;
        RECT 1838.690 1088.380 1839.010 1088.440 ;
        RECT 1841.450 1088.380 1841.770 1088.440 ;
        RECT 1841.450 24.380 1841.770 24.440 ;
        RECT 2881.050 24.380 2881.370 24.440 ;
        RECT 1841.450 24.240 2881.370 24.380 ;
        RECT 1841.450 24.180 1841.770 24.240 ;
        RECT 2881.050 24.180 2881.370 24.240 ;
      LAYER via ;
        RECT 1838.720 1088.380 1838.980 1088.640 ;
        RECT 1841.480 1088.380 1841.740 1088.640 ;
        RECT 1841.480 24.180 1841.740 24.440 ;
        RECT 2881.080 24.180 2881.340 24.440 ;
      LAYER met2 ;
        RECT 1838.630 1100.580 1838.910 1104.000 ;
        RECT 1838.630 1100.000 1838.920 1100.580 ;
        RECT 1838.780 1088.670 1838.920 1100.000 ;
        RECT 1838.720 1088.350 1838.980 1088.670 ;
        RECT 1841.480 1088.350 1841.740 1088.670 ;
        RECT 1841.540 24.470 1841.680 1088.350 ;
        RECT 1841.480 24.150 1841.740 24.470 ;
        RECT 2881.080 24.150 2881.340 24.470 ;
        RECT 2881.140 2.000 2881.280 24.150 ;
        RECT 2880.930 -4.000 2881.490 2.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1844.670 1088.580 1844.990 1088.640 ;
        RECT 1848.350 1088.580 1848.670 1088.640 ;
        RECT 1844.670 1088.440 1848.670 1088.580 ;
        RECT 1844.670 1088.380 1844.990 1088.440 ;
        RECT 1848.350 1088.380 1848.670 1088.440 ;
        RECT 1848.350 24.040 1848.670 24.100 ;
        RECT 2898.990 24.040 2899.310 24.100 ;
        RECT 1848.350 23.900 2899.310 24.040 ;
        RECT 1848.350 23.840 1848.670 23.900 ;
        RECT 2898.990 23.840 2899.310 23.900 ;
      LAYER via ;
        RECT 1844.700 1088.380 1844.960 1088.640 ;
        RECT 1848.380 1088.380 1848.640 1088.640 ;
        RECT 1848.380 23.840 1848.640 24.100 ;
        RECT 2899.020 23.840 2899.280 24.100 ;
      LAYER met2 ;
        RECT 1844.610 1100.580 1844.890 1104.000 ;
        RECT 1844.610 1100.000 1844.900 1100.580 ;
        RECT 1844.760 1088.670 1844.900 1100.000 ;
        RECT 1844.700 1088.350 1844.960 1088.670 ;
        RECT 1848.380 1088.350 1848.640 1088.670 ;
        RECT 1848.440 24.130 1848.580 1088.350 ;
        RECT 1848.380 23.810 1848.640 24.130 ;
        RECT 2899.020 23.810 2899.280 24.130 ;
        RECT 2899.080 2.000 2899.220 23.810 ;
        RECT 2898.870 -4.000 2899.430 2.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 846.930 42.400 847.250 42.460 ;
        RECT 1139.950 42.400 1140.270 42.460 ;
        RECT 846.930 42.260 1140.270 42.400 ;
        RECT 846.930 42.200 847.250 42.260 ;
        RECT 1139.950 42.200 1140.270 42.260 ;
      LAYER via ;
        RECT 846.960 42.200 847.220 42.460 ;
        RECT 1139.980 42.200 1140.240 42.460 ;
      LAYER met2 ;
        RECT 1140.810 1100.650 1141.090 1104.000 ;
        RECT 1140.040 1100.510 1141.090 1100.650 ;
        RECT 1140.040 42.490 1140.180 1100.510 ;
        RECT 1140.810 1100.000 1141.090 1100.510 ;
        RECT 846.960 42.170 847.220 42.490 ;
        RECT 1139.980 42.170 1140.240 42.490 ;
        RECT 847.020 2.000 847.160 42.170 ;
        RECT 846.810 -4.000 847.370 2.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1146.925 820.845 1147.095 862.495 ;
        RECT 1146.465 766.105 1146.635 814.215 ;
        RECT 1146.005 589.985 1146.175 613.955 ;
      LAYER mcon ;
        RECT 1146.925 862.325 1147.095 862.495 ;
        RECT 1146.465 814.045 1146.635 814.215 ;
        RECT 1146.005 613.785 1146.175 613.955 ;
      LAYER met1 ;
        RECT 1147.310 1000.520 1147.630 1000.580 ;
        RECT 1147.770 1000.520 1148.090 1000.580 ;
        RECT 1147.310 1000.380 1148.090 1000.520 ;
        RECT 1147.310 1000.320 1147.630 1000.380 ;
        RECT 1147.770 1000.320 1148.090 1000.380 ;
        RECT 1146.390 910.760 1146.710 910.820 ;
        RECT 1147.310 910.760 1147.630 910.820 ;
        RECT 1146.390 910.620 1147.630 910.760 ;
        RECT 1146.390 910.560 1146.710 910.620 ;
        RECT 1147.310 910.560 1147.630 910.620 ;
        RECT 1146.850 862.480 1147.170 862.540 ;
        RECT 1146.655 862.340 1147.170 862.480 ;
        RECT 1146.850 862.280 1147.170 862.340 ;
        RECT 1146.850 821.000 1147.170 821.060 ;
        RECT 1146.655 820.860 1147.170 821.000 ;
        RECT 1146.850 820.800 1147.170 820.860 ;
        RECT 1146.405 814.200 1146.695 814.245 ;
        RECT 1147.310 814.200 1147.630 814.260 ;
        RECT 1146.405 814.060 1147.630 814.200 ;
        RECT 1146.405 814.015 1146.695 814.060 ;
        RECT 1147.310 814.000 1147.630 814.060 ;
        RECT 1146.390 766.260 1146.710 766.320 ;
        RECT 1146.195 766.120 1146.710 766.260 ;
        RECT 1146.390 766.060 1146.710 766.120 ;
        RECT 1146.390 710.500 1146.710 710.560 ;
        RECT 1146.850 710.500 1147.170 710.560 ;
        RECT 1146.390 710.360 1147.170 710.500 ;
        RECT 1146.390 710.300 1146.710 710.360 ;
        RECT 1146.850 710.300 1147.170 710.360 ;
        RECT 1145.945 613.940 1146.235 613.985 ;
        RECT 1146.390 613.940 1146.710 614.000 ;
        RECT 1145.945 613.800 1146.710 613.940 ;
        RECT 1145.945 613.755 1146.235 613.800 ;
        RECT 1146.390 613.740 1146.710 613.800 ;
        RECT 1145.945 590.140 1146.235 590.185 ;
        RECT 1146.390 590.140 1146.710 590.200 ;
        RECT 1145.945 590.000 1146.710 590.140 ;
        RECT 1145.945 589.955 1146.235 590.000 ;
        RECT 1146.390 589.940 1146.710 590.000 ;
        RECT 1146.390 434.560 1146.710 434.820 ;
        RECT 1146.480 434.420 1146.620 434.560 ;
        RECT 1146.850 434.420 1147.170 434.480 ;
        RECT 1146.480 434.280 1147.170 434.420 ;
        RECT 1146.850 434.220 1147.170 434.280 ;
        RECT 1146.850 387.300 1147.170 387.560 ;
        RECT 1146.940 386.880 1147.080 387.300 ;
        RECT 1146.850 386.620 1147.170 386.880 ;
        RECT 1146.390 337.660 1146.710 337.920 ;
        RECT 1146.480 337.520 1146.620 337.660 ;
        RECT 1146.850 337.520 1147.170 337.580 ;
        RECT 1146.480 337.380 1147.170 337.520 ;
        RECT 1146.850 337.320 1147.170 337.380 ;
        RECT 1146.850 255.380 1147.170 255.640 ;
        RECT 1146.940 254.960 1147.080 255.380 ;
        RECT 1146.850 254.700 1147.170 254.960 ;
        RECT 1146.390 193.020 1146.710 193.080 ;
        RECT 1146.850 193.020 1147.170 193.080 ;
        RECT 1146.390 192.880 1147.170 193.020 ;
        RECT 1146.390 192.820 1146.710 192.880 ;
        RECT 1146.850 192.820 1147.170 192.880 ;
        RECT 1146.390 96.800 1146.710 96.860 ;
        RECT 1146.850 96.800 1147.170 96.860 ;
        RECT 1146.390 96.660 1147.170 96.800 ;
        RECT 1146.390 96.600 1146.710 96.660 ;
        RECT 1146.850 96.600 1147.170 96.660 ;
        RECT 864.870 42.060 865.190 42.120 ;
        RECT 1146.850 42.060 1147.170 42.120 ;
        RECT 864.870 41.920 1147.170 42.060 ;
        RECT 864.870 41.860 865.190 41.920 ;
        RECT 1146.850 41.860 1147.170 41.920 ;
      LAYER via ;
        RECT 1147.340 1000.320 1147.600 1000.580 ;
        RECT 1147.800 1000.320 1148.060 1000.580 ;
        RECT 1146.420 910.560 1146.680 910.820 ;
        RECT 1147.340 910.560 1147.600 910.820 ;
        RECT 1146.880 862.280 1147.140 862.540 ;
        RECT 1146.880 820.800 1147.140 821.060 ;
        RECT 1147.340 814.000 1147.600 814.260 ;
        RECT 1146.420 766.060 1146.680 766.320 ;
        RECT 1146.420 710.300 1146.680 710.560 ;
        RECT 1146.880 710.300 1147.140 710.560 ;
        RECT 1146.420 613.740 1146.680 614.000 ;
        RECT 1146.420 589.940 1146.680 590.200 ;
        RECT 1146.420 434.560 1146.680 434.820 ;
        RECT 1146.880 434.220 1147.140 434.480 ;
        RECT 1146.880 387.300 1147.140 387.560 ;
        RECT 1146.880 386.620 1147.140 386.880 ;
        RECT 1146.420 337.660 1146.680 337.920 ;
        RECT 1146.880 337.320 1147.140 337.580 ;
        RECT 1146.880 255.380 1147.140 255.640 ;
        RECT 1146.880 254.700 1147.140 254.960 ;
        RECT 1146.420 192.820 1146.680 193.080 ;
        RECT 1146.880 192.820 1147.140 193.080 ;
        RECT 1146.420 96.600 1146.680 96.860 ;
        RECT 1146.880 96.600 1147.140 96.860 ;
        RECT 864.900 41.860 865.160 42.120 ;
        RECT 1146.880 41.860 1147.140 42.120 ;
      LAYER met2 ;
        RECT 1146.790 1100.580 1147.070 1104.000 ;
        RECT 1146.790 1100.000 1147.080 1100.580 ;
        RECT 1146.940 1062.685 1147.080 1100.000 ;
        RECT 1146.870 1062.315 1147.150 1062.685 ;
        RECT 1147.790 1062.315 1148.070 1062.685 ;
        RECT 1147.860 1051.690 1148.000 1062.315 ;
        RECT 1147.400 1051.550 1148.000 1051.690 ;
        RECT 1147.400 1000.610 1147.540 1051.550 ;
        RECT 1147.340 1000.290 1147.600 1000.610 ;
        RECT 1147.800 1000.290 1148.060 1000.610 ;
        RECT 1147.860 911.045 1148.000 1000.290 ;
        RECT 1146.410 910.675 1146.690 911.045 ;
        RECT 1146.420 910.530 1146.680 910.675 ;
        RECT 1147.340 910.530 1147.600 910.850 ;
        RECT 1147.790 910.675 1148.070 911.045 ;
        RECT 1147.400 882.370 1147.540 910.530 ;
        RECT 1146.940 882.230 1147.540 882.370 ;
        RECT 1146.940 862.570 1147.080 882.230 ;
        RECT 1146.880 862.250 1147.140 862.570 ;
        RECT 1146.880 820.770 1147.140 821.090 ;
        RECT 1146.940 814.370 1147.080 820.770 ;
        RECT 1146.940 814.290 1147.540 814.370 ;
        RECT 1146.940 814.230 1147.600 814.290 ;
        RECT 1147.340 813.970 1147.600 814.230 ;
        RECT 1146.420 766.030 1146.680 766.350 ;
        RECT 1146.480 710.590 1146.620 766.030 ;
        RECT 1146.420 710.270 1146.680 710.590 ;
        RECT 1146.880 710.270 1147.140 710.590 ;
        RECT 1146.940 628.845 1147.080 710.270 ;
        RECT 1146.870 628.475 1147.150 628.845 ;
        RECT 1146.410 627.795 1146.690 628.165 ;
        RECT 1146.480 614.030 1146.620 627.795 ;
        RECT 1146.420 613.710 1146.680 614.030 ;
        RECT 1146.420 589.910 1146.680 590.230 ;
        RECT 1146.480 500.210 1146.620 589.910 ;
        RECT 1146.480 500.070 1147.540 500.210 ;
        RECT 1147.400 496.130 1147.540 500.070 ;
        RECT 1146.940 495.990 1147.540 496.130 ;
        RECT 1146.940 459.410 1147.080 495.990 ;
        RECT 1146.940 459.270 1147.540 459.410 ;
        RECT 1147.400 435.045 1147.540 459.270 ;
        RECT 1146.410 434.675 1146.690 435.045 ;
        RECT 1147.330 434.675 1147.610 435.045 ;
        RECT 1146.420 434.530 1146.680 434.675 ;
        RECT 1146.880 434.190 1147.140 434.510 ;
        RECT 1146.940 387.590 1147.080 434.190 ;
        RECT 1146.880 387.270 1147.140 387.590 ;
        RECT 1146.880 386.590 1147.140 386.910 ;
        RECT 1146.940 385.970 1147.080 386.590 ;
        RECT 1146.480 385.830 1147.080 385.970 ;
        RECT 1146.480 337.950 1146.620 385.830 ;
        RECT 1146.420 337.630 1146.680 337.950 ;
        RECT 1146.880 337.290 1147.140 337.610 ;
        RECT 1146.940 255.670 1147.080 337.290 ;
        RECT 1146.880 255.350 1147.140 255.670 ;
        RECT 1146.880 254.670 1147.140 254.990 ;
        RECT 1146.940 193.110 1147.080 254.670 ;
        RECT 1146.420 192.790 1146.680 193.110 ;
        RECT 1146.880 192.790 1147.140 193.110 ;
        RECT 1146.480 96.890 1146.620 192.790 ;
        RECT 1146.420 96.570 1146.680 96.890 ;
        RECT 1146.880 96.570 1147.140 96.890 ;
        RECT 1146.940 42.150 1147.080 96.570 ;
        RECT 864.900 41.830 865.160 42.150 ;
        RECT 1146.880 41.830 1147.140 42.150 ;
        RECT 864.960 2.000 865.100 41.830 ;
        RECT 864.750 -4.000 865.310 2.000 ;
      LAYER via2 ;
        RECT 1146.870 1062.360 1147.150 1062.640 ;
        RECT 1147.790 1062.360 1148.070 1062.640 ;
        RECT 1146.410 910.720 1146.690 911.000 ;
        RECT 1147.790 910.720 1148.070 911.000 ;
        RECT 1146.870 628.520 1147.150 628.800 ;
        RECT 1146.410 627.840 1146.690 628.120 ;
        RECT 1146.410 434.720 1146.690 435.000 ;
        RECT 1147.330 434.720 1147.610 435.000 ;
      LAYER met3 ;
        RECT 1146.845 1062.650 1147.175 1062.665 ;
        RECT 1147.765 1062.650 1148.095 1062.665 ;
        RECT 1146.845 1062.350 1148.095 1062.650 ;
        RECT 1146.845 1062.335 1147.175 1062.350 ;
        RECT 1147.765 1062.335 1148.095 1062.350 ;
        RECT 1146.385 911.010 1146.715 911.025 ;
        RECT 1147.765 911.010 1148.095 911.025 ;
        RECT 1146.385 910.710 1148.095 911.010 ;
        RECT 1146.385 910.695 1146.715 910.710 ;
        RECT 1147.765 910.695 1148.095 910.710 ;
        RECT 1146.845 628.810 1147.175 628.825 ;
        RECT 1146.630 628.495 1147.175 628.810 ;
        RECT 1146.630 628.145 1146.930 628.495 ;
        RECT 1146.385 627.830 1146.930 628.145 ;
        RECT 1146.385 627.815 1146.715 627.830 ;
        RECT 1146.385 435.010 1146.715 435.025 ;
        RECT 1147.305 435.010 1147.635 435.025 ;
        RECT 1146.385 434.710 1147.635 435.010 ;
        RECT 1146.385 434.695 1146.715 434.710 ;
        RECT 1147.305 434.695 1147.635 434.710 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1152.830 955.640 1153.150 955.700 ;
        RECT 1153.750 955.640 1154.070 955.700 ;
        RECT 1152.830 955.500 1154.070 955.640 ;
        RECT 1152.830 955.440 1153.150 955.500 ;
        RECT 1153.750 955.440 1154.070 955.500 ;
        RECT 1152.830 907.360 1153.150 907.420 ;
        RECT 1153.750 907.360 1154.070 907.420 ;
        RECT 1152.830 907.220 1154.070 907.360 ;
        RECT 1152.830 907.160 1153.150 907.220 ;
        RECT 1153.750 907.160 1154.070 907.220 ;
        RECT 1152.830 760.480 1153.150 760.540 ;
        RECT 1153.750 760.480 1154.070 760.540 ;
        RECT 1152.830 760.340 1154.070 760.480 ;
        RECT 1152.830 760.280 1153.150 760.340 ;
        RECT 1153.750 760.280 1154.070 760.340 ;
        RECT 1152.830 714.240 1153.150 714.300 ;
        RECT 1153.750 714.240 1154.070 714.300 ;
        RECT 1152.830 714.100 1154.070 714.240 ;
        RECT 1152.830 714.040 1153.150 714.100 ;
        RECT 1153.750 714.040 1154.070 714.100 ;
        RECT 1153.750 569.400 1154.070 569.460 ;
        RECT 1154.670 569.400 1154.990 569.460 ;
        RECT 1153.750 569.260 1154.990 569.400 ;
        RECT 1153.750 569.200 1154.070 569.260 ;
        RECT 1154.670 569.200 1154.990 569.260 ;
        RECT 1153.750 521.120 1154.070 521.180 ;
        RECT 1154.670 521.120 1154.990 521.180 ;
        RECT 1153.750 520.980 1154.990 521.120 ;
        RECT 1153.750 520.920 1154.070 520.980 ;
        RECT 1154.670 520.920 1154.990 520.980 ;
        RECT 1153.750 472.840 1154.070 472.900 ;
        RECT 1154.670 472.840 1154.990 472.900 ;
        RECT 1153.750 472.700 1154.990 472.840 ;
        RECT 1153.750 472.640 1154.070 472.700 ;
        RECT 1154.670 472.640 1154.990 472.700 ;
        RECT 1153.750 424.560 1154.070 424.620 ;
        RECT 1154.670 424.560 1154.990 424.620 ;
        RECT 1153.750 424.420 1154.990 424.560 ;
        RECT 1153.750 424.360 1154.070 424.420 ;
        RECT 1154.670 424.360 1154.990 424.420 ;
        RECT 1153.750 376.280 1154.070 376.340 ;
        RECT 1154.670 376.280 1154.990 376.340 ;
        RECT 1153.750 376.140 1154.990 376.280 ;
        RECT 1153.750 376.080 1154.070 376.140 ;
        RECT 1154.670 376.080 1154.990 376.140 ;
        RECT 1153.750 193.360 1154.070 193.420 ;
        RECT 1154.670 193.360 1154.990 193.420 ;
        RECT 1153.750 193.220 1154.990 193.360 ;
        RECT 1153.750 193.160 1154.070 193.220 ;
        RECT 1154.670 193.160 1154.990 193.220 ;
        RECT 1152.830 83.880 1153.150 83.940 ;
        RECT 1153.750 83.880 1154.070 83.940 ;
        RECT 1152.830 83.740 1154.070 83.880 ;
        RECT 1152.830 83.680 1153.150 83.740 ;
        RECT 1153.750 83.680 1154.070 83.740 ;
        RECT 882.810 44.780 883.130 44.840 ;
        RECT 1152.830 44.780 1153.150 44.840 ;
        RECT 882.810 44.640 1153.150 44.780 ;
        RECT 882.810 44.580 883.130 44.640 ;
        RECT 1152.830 44.580 1153.150 44.640 ;
      LAYER via ;
        RECT 1152.860 955.440 1153.120 955.700 ;
        RECT 1153.780 955.440 1154.040 955.700 ;
        RECT 1152.860 907.160 1153.120 907.420 ;
        RECT 1153.780 907.160 1154.040 907.420 ;
        RECT 1152.860 760.280 1153.120 760.540 ;
        RECT 1153.780 760.280 1154.040 760.540 ;
        RECT 1152.860 714.040 1153.120 714.300 ;
        RECT 1153.780 714.040 1154.040 714.300 ;
        RECT 1153.780 569.200 1154.040 569.460 ;
        RECT 1154.700 569.200 1154.960 569.460 ;
        RECT 1153.780 520.920 1154.040 521.180 ;
        RECT 1154.700 520.920 1154.960 521.180 ;
        RECT 1153.780 472.640 1154.040 472.900 ;
        RECT 1154.700 472.640 1154.960 472.900 ;
        RECT 1153.780 424.360 1154.040 424.620 ;
        RECT 1154.700 424.360 1154.960 424.620 ;
        RECT 1153.780 376.080 1154.040 376.340 ;
        RECT 1154.700 376.080 1154.960 376.340 ;
        RECT 1153.780 193.160 1154.040 193.420 ;
        RECT 1154.700 193.160 1154.960 193.420 ;
        RECT 1152.860 83.680 1153.120 83.940 ;
        RECT 1153.780 83.680 1154.040 83.940 ;
        RECT 882.840 44.580 883.100 44.840 ;
        RECT 1152.860 44.580 1153.120 44.840 ;
      LAYER met2 ;
        RECT 1152.770 1101.330 1153.050 1104.000 ;
        RECT 1152.770 1101.190 1153.980 1101.330 ;
        RECT 1152.770 1100.000 1153.050 1101.190 ;
        RECT 1153.840 955.730 1153.980 1101.190 ;
        RECT 1152.860 955.410 1153.120 955.730 ;
        RECT 1153.780 955.410 1154.040 955.730 ;
        RECT 1152.920 907.450 1153.060 955.410 ;
        RECT 1152.860 907.130 1153.120 907.450 ;
        RECT 1153.780 907.130 1154.040 907.450 ;
        RECT 1153.840 859.250 1153.980 907.130 ;
        RECT 1153.840 859.110 1154.900 859.250 ;
        RECT 1154.760 811.650 1154.900 859.110 ;
        RECT 1153.840 811.510 1154.900 811.650 ;
        RECT 1153.840 760.570 1153.980 811.510 ;
        RECT 1152.860 760.250 1153.120 760.570 ;
        RECT 1153.780 760.250 1154.040 760.570 ;
        RECT 1152.920 714.330 1153.060 760.250 ;
        RECT 1152.860 714.010 1153.120 714.330 ;
        RECT 1153.780 714.010 1154.040 714.330 ;
        RECT 1153.840 666.130 1153.980 714.010 ;
        RECT 1153.840 665.990 1154.900 666.130 ;
        RECT 1154.760 617.850 1154.900 665.990 ;
        RECT 1153.840 617.710 1154.900 617.850 ;
        RECT 1153.840 569.490 1153.980 617.710 ;
        RECT 1153.780 569.170 1154.040 569.490 ;
        RECT 1154.700 569.170 1154.960 569.490 ;
        RECT 1154.760 521.210 1154.900 569.170 ;
        RECT 1153.780 520.890 1154.040 521.210 ;
        RECT 1154.700 520.890 1154.960 521.210 ;
        RECT 1153.840 472.930 1153.980 520.890 ;
        RECT 1153.780 472.610 1154.040 472.930 ;
        RECT 1154.700 472.610 1154.960 472.930 ;
        RECT 1154.760 424.650 1154.900 472.610 ;
        RECT 1153.780 424.330 1154.040 424.650 ;
        RECT 1154.700 424.330 1154.960 424.650 ;
        RECT 1153.840 376.370 1153.980 424.330 ;
        RECT 1153.780 376.050 1154.040 376.370 ;
        RECT 1154.700 376.050 1154.960 376.370 ;
        RECT 1154.760 305.050 1154.900 376.050 ;
        RECT 1153.840 304.910 1154.900 305.050 ;
        RECT 1153.840 279.210 1153.980 304.910 ;
        RECT 1153.840 279.070 1154.900 279.210 ;
        RECT 1154.760 193.450 1154.900 279.070 ;
        RECT 1153.780 193.130 1154.040 193.450 ;
        RECT 1154.700 193.130 1154.960 193.450 ;
        RECT 1153.840 182.650 1153.980 193.130 ;
        RECT 1153.840 182.510 1154.900 182.650 ;
        RECT 1154.760 134.370 1154.900 182.510 ;
        RECT 1153.840 134.230 1154.900 134.370 ;
        RECT 1153.840 83.970 1153.980 134.230 ;
        RECT 1152.860 83.650 1153.120 83.970 ;
        RECT 1153.780 83.650 1154.040 83.970 ;
        RECT 1152.920 44.870 1153.060 83.650 ;
        RECT 882.840 44.550 883.100 44.870 ;
        RECT 1152.860 44.550 1153.120 44.870 ;
        RECT 882.900 2.000 883.040 44.550 ;
        RECT 882.690 -4.000 883.250 2.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1154.745 724.285 1154.915 765.935 ;
        RECT 1155.205 572.645 1155.375 620.755 ;
        RECT 1153.825 282.965 1153.995 329.715 ;
      LAYER mcon ;
        RECT 1154.745 765.765 1154.915 765.935 ;
        RECT 1155.205 620.585 1155.375 620.755 ;
        RECT 1153.825 329.545 1153.995 329.715 ;
      LAYER met1 ;
        RECT 1154.210 1000.520 1154.530 1000.580 ;
        RECT 1156.970 1000.520 1157.290 1000.580 ;
        RECT 1154.210 1000.380 1157.290 1000.520 ;
        RECT 1154.210 1000.320 1154.530 1000.380 ;
        RECT 1156.970 1000.320 1157.290 1000.380 ;
        RECT 1155.130 932.180 1155.450 932.240 ;
        RECT 1154.760 932.040 1155.450 932.180 ;
        RECT 1154.760 931.560 1154.900 932.040 ;
        RECT 1155.130 931.980 1155.450 932.040 ;
        RECT 1154.670 931.300 1154.990 931.560 ;
        RECT 1154.670 910.760 1154.990 910.820 ;
        RECT 1155.130 910.760 1155.450 910.820 ;
        RECT 1154.670 910.620 1155.450 910.760 ;
        RECT 1154.670 910.560 1154.990 910.620 ;
        RECT 1155.130 910.560 1155.450 910.620 ;
        RECT 1154.670 765.920 1154.990 765.980 ;
        RECT 1154.475 765.780 1154.990 765.920 ;
        RECT 1154.670 765.720 1154.990 765.780 ;
        RECT 1154.670 724.440 1154.990 724.500 ;
        RECT 1154.475 724.300 1154.990 724.440 ;
        RECT 1154.670 724.240 1154.990 724.300 ;
        RECT 1155.130 676.160 1155.450 676.220 ;
        RECT 1156.050 676.160 1156.370 676.220 ;
        RECT 1155.130 676.020 1156.370 676.160 ;
        RECT 1155.130 675.960 1155.450 676.020 ;
        RECT 1156.050 675.960 1156.370 676.020 ;
        RECT 1155.145 620.740 1155.435 620.785 ;
        RECT 1155.590 620.740 1155.910 620.800 ;
        RECT 1155.145 620.600 1155.910 620.740 ;
        RECT 1155.145 620.555 1155.435 620.600 ;
        RECT 1155.590 620.540 1155.910 620.600 ;
        RECT 1155.130 572.800 1155.450 572.860 ;
        RECT 1154.935 572.660 1155.450 572.800 ;
        RECT 1155.130 572.600 1155.450 572.660 ;
        RECT 1153.750 555.460 1154.070 555.520 ;
        RECT 1155.130 555.460 1155.450 555.520 ;
        RECT 1153.750 555.320 1155.450 555.460 ;
        RECT 1153.750 555.260 1154.070 555.320 ;
        RECT 1155.130 555.260 1155.450 555.320 ;
        RECT 1153.750 329.700 1154.070 329.760 ;
        RECT 1153.555 329.560 1154.070 329.700 ;
        RECT 1153.750 329.500 1154.070 329.560 ;
        RECT 1153.765 283.120 1154.055 283.165 ;
        RECT 1155.130 283.120 1155.450 283.180 ;
        RECT 1153.765 282.980 1155.450 283.120 ;
        RECT 1153.765 282.935 1154.055 282.980 ;
        RECT 1155.130 282.920 1155.450 282.980 ;
        RECT 1155.130 282.440 1155.450 282.500 ;
        RECT 1156.970 282.440 1157.290 282.500 ;
        RECT 1155.130 282.300 1157.290 282.440 ;
        RECT 1155.130 282.240 1155.450 282.300 ;
        RECT 1156.970 282.240 1157.290 282.300 ;
        RECT 1156.050 227.700 1156.370 227.760 ;
        RECT 1156.510 227.700 1156.830 227.760 ;
        RECT 1156.050 227.560 1156.830 227.700 ;
        RECT 1156.050 227.500 1156.370 227.560 ;
        RECT 1156.510 227.500 1156.830 227.560 ;
        RECT 1156.510 145.420 1156.830 145.480 ;
        RECT 1155.680 145.280 1156.830 145.420 ;
        RECT 1155.680 144.800 1155.820 145.280 ;
        RECT 1156.510 145.220 1156.830 145.280 ;
        RECT 1155.590 144.540 1155.910 144.800 ;
        RECT 1154.670 133.180 1154.990 133.240 ;
        RECT 1155.590 133.180 1155.910 133.240 ;
        RECT 1154.670 133.040 1155.910 133.180 ;
        RECT 1154.670 132.980 1154.990 133.040 ;
        RECT 1155.590 132.980 1155.910 133.040 ;
        RECT 900.750 45.460 901.070 45.520 ;
        RECT 1154.670 45.460 1154.990 45.520 ;
        RECT 900.750 45.320 1154.990 45.460 ;
        RECT 900.750 45.260 901.070 45.320 ;
        RECT 1154.670 45.260 1154.990 45.320 ;
      LAYER via ;
        RECT 1154.240 1000.320 1154.500 1000.580 ;
        RECT 1157.000 1000.320 1157.260 1000.580 ;
        RECT 1155.160 931.980 1155.420 932.240 ;
        RECT 1154.700 931.300 1154.960 931.560 ;
        RECT 1154.700 910.560 1154.960 910.820 ;
        RECT 1155.160 910.560 1155.420 910.820 ;
        RECT 1154.700 765.720 1154.960 765.980 ;
        RECT 1154.700 724.240 1154.960 724.500 ;
        RECT 1155.160 675.960 1155.420 676.220 ;
        RECT 1156.080 675.960 1156.340 676.220 ;
        RECT 1155.620 620.540 1155.880 620.800 ;
        RECT 1155.160 572.600 1155.420 572.860 ;
        RECT 1153.780 555.260 1154.040 555.520 ;
        RECT 1155.160 555.260 1155.420 555.520 ;
        RECT 1153.780 329.500 1154.040 329.760 ;
        RECT 1155.160 282.920 1155.420 283.180 ;
        RECT 1155.160 282.240 1155.420 282.500 ;
        RECT 1157.000 282.240 1157.260 282.500 ;
        RECT 1156.080 227.500 1156.340 227.760 ;
        RECT 1156.540 227.500 1156.800 227.760 ;
        RECT 1156.540 145.220 1156.800 145.480 ;
        RECT 1155.620 144.540 1155.880 144.800 ;
        RECT 1154.700 132.980 1154.960 133.240 ;
        RECT 1155.620 132.980 1155.880 133.240 ;
        RECT 900.780 45.260 901.040 45.520 ;
        RECT 1154.700 45.260 1154.960 45.520 ;
      LAYER met2 ;
        RECT 1158.750 1100.650 1159.030 1104.000 ;
        RECT 1158.440 1100.510 1159.030 1100.650 ;
        RECT 1158.440 1076.170 1158.580 1100.510 ;
        RECT 1158.750 1100.000 1159.030 1100.510 ;
        RECT 1157.060 1076.030 1158.580 1076.170 ;
        RECT 1157.060 1000.610 1157.200 1076.030 ;
        RECT 1154.240 1000.290 1154.500 1000.610 ;
        RECT 1157.000 1000.290 1157.260 1000.610 ;
        RECT 1154.300 952.525 1154.440 1000.290 ;
        RECT 1154.230 952.155 1154.510 952.525 ;
        RECT 1155.150 952.155 1155.430 952.525 ;
        RECT 1155.220 932.270 1155.360 952.155 ;
        RECT 1155.160 931.950 1155.420 932.270 ;
        RECT 1154.700 931.270 1154.960 931.590 ;
        RECT 1154.760 910.850 1154.900 931.270 ;
        RECT 1154.700 910.530 1154.960 910.850 ;
        RECT 1155.160 910.530 1155.420 910.850 ;
        RECT 1155.220 845.650 1155.360 910.530 ;
        RECT 1155.220 845.510 1156.280 845.650 ;
        RECT 1156.140 773.005 1156.280 845.510 ;
        RECT 1154.690 772.635 1154.970 773.005 ;
        RECT 1156.070 772.635 1156.350 773.005 ;
        RECT 1154.760 766.010 1154.900 772.635 ;
        RECT 1154.700 765.690 1154.960 766.010 ;
        RECT 1154.700 724.210 1154.960 724.530 ;
        RECT 1154.760 717.810 1154.900 724.210 ;
        RECT 1154.760 717.670 1155.360 717.810 ;
        RECT 1155.220 676.250 1155.360 717.670 ;
        RECT 1155.160 675.930 1155.420 676.250 ;
        RECT 1156.080 675.930 1156.340 676.250 ;
        RECT 1156.140 645.050 1156.280 675.930 ;
        RECT 1155.680 644.910 1156.280 645.050 ;
        RECT 1155.680 620.830 1155.820 644.910 ;
        RECT 1155.620 620.510 1155.880 620.830 ;
        RECT 1155.160 572.570 1155.420 572.890 ;
        RECT 1155.220 555.550 1155.360 572.570 ;
        RECT 1153.780 555.230 1154.040 555.550 ;
        RECT 1155.160 555.230 1155.420 555.550 ;
        RECT 1153.840 521.970 1153.980 555.230 ;
        RECT 1153.840 521.830 1154.440 521.970 ;
        RECT 1154.300 472.330 1154.440 521.830 ;
        RECT 1153.840 472.190 1154.440 472.330 ;
        RECT 1153.840 425.410 1153.980 472.190 ;
        RECT 1153.840 425.270 1154.440 425.410 ;
        RECT 1154.300 375.770 1154.440 425.270 ;
        RECT 1153.840 375.630 1154.440 375.770 ;
        RECT 1153.840 329.790 1153.980 375.630 ;
        RECT 1153.780 329.470 1154.040 329.790 ;
        RECT 1155.160 282.890 1155.420 283.210 ;
        RECT 1155.220 282.530 1155.360 282.890 ;
        RECT 1155.160 282.210 1155.420 282.530 ;
        RECT 1157.000 282.210 1157.260 282.530 ;
        RECT 1157.060 235.010 1157.200 282.210 ;
        RECT 1156.140 234.870 1157.200 235.010 ;
        RECT 1156.140 227.790 1156.280 234.870 ;
        RECT 1156.080 227.470 1156.340 227.790 ;
        RECT 1156.540 227.470 1156.800 227.790 ;
        RECT 1156.600 145.510 1156.740 227.470 ;
        RECT 1156.540 145.190 1156.800 145.510 ;
        RECT 1155.620 144.510 1155.880 144.830 ;
        RECT 1155.680 133.270 1155.820 144.510 ;
        RECT 1154.700 132.950 1154.960 133.270 ;
        RECT 1155.620 132.950 1155.880 133.270 ;
        RECT 1154.760 45.550 1154.900 132.950 ;
        RECT 900.780 45.230 901.040 45.550 ;
        RECT 1154.700 45.230 1154.960 45.550 ;
        RECT 900.840 2.000 900.980 45.230 ;
        RECT 900.630 -4.000 901.190 2.000 ;
      LAYER via2 ;
        RECT 1154.230 952.200 1154.510 952.480 ;
        RECT 1155.150 952.200 1155.430 952.480 ;
        RECT 1154.690 772.680 1154.970 772.960 ;
        RECT 1156.070 772.680 1156.350 772.960 ;
      LAYER met3 ;
        RECT 1154.205 952.490 1154.535 952.505 ;
        RECT 1155.125 952.490 1155.455 952.505 ;
        RECT 1154.205 952.190 1155.455 952.490 ;
        RECT 1154.205 952.175 1154.535 952.190 ;
        RECT 1155.125 952.175 1155.455 952.190 ;
        RECT 1154.665 772.970 1154.995 772.985 ;
        RECT 1156.045 772.970 1156.375 772.985 ;
        RECT 1154.665 772.670 1156.375 772.970 ;
        RECT 1154.665 772.655 1154.995 772.670 ;
        RECT 1156.045 772.655 1156.375 772.670 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1159.270 1052.200 1159.590 1052.260 ;
        RECT 1163.870 1052.200 1164.190 1052.260 ;
        RECT 1159.270 1052.060 1164.190 1052.200 ;
        RECT 1159.270 1052.000 1159.590 1052.060 ;
        RECT 1163.870 1052.000 1164.190 1052.060 ;
        RECT 918.690 17.920 919.010 17.980 ;
        RECT 1159.270 17.920 1159.590 17.980 ;
        RECT 918.690 17.780 1159.590 17.920 ;
        RECT 918.690 17.720 919.010 17.780 ;
        RECT 1159.270 17.720 1159.590 17.780 ;
      LAYER via ;
        RECT 1159.300 1052.000 1159.560 1052.260 ;
        RECT 1163.900 1052.000 1164.160 1052.260 ;
        RECT 918.720 17.720 918.980 17.980 ;
        RECT 1159.300 17.720 1159.560 17.980 ;
      LAYER met2 ;
        RECT 1165.190 1100.650 1165.470 1104.000 ;
        RECT 1163.960 1100.510 1165.470 1100.650 ;
        RECT 1163.960 1052.290 1164.100 1100.510 ;
        RECT 1165.190 1100.000 1165.470 1100.510 ;
        RECT 1159.300 1051.970 1159.560 1052.290 ;
        RECT 1163.900 1051.970 1164.160 1052.290 ;
        RECT 1159.360 18.010 1159.500 1051.970 ;
        RECT 918.720 17.690 918.980 18.010 ;
        RECT 1159.300 17.690 1159.560 18.010 ;
        RECT 918.780 2.000 918.920 17.690 ;
        RECT 918.570 -4.000 919.130 2.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1166.630 1052.200 1166.950 1052.260 ;
        RECT 1169.850 1052.200 1170.170 1052.260 ;
        RECT 1166.630 1052.060 1170.170 1052.200 ;
        RECT 1166.630 1052.000 1166.950 1052.060 ;
        RECT 1169.850 1052.000 1170.170 1052.060 ;
        RECT 936.170 24.720 936.490 24.780 ;
        RECT 1166.630 24.720 1166.950 24.780 ;
        RECT 936.170 24.580 1166.950 24.720 ;
        RECT 936.170 24.520 936.490 24.580 ;
        RECT 1166.630 24.520 1166.950 24.580 ;
      LAYER via ;
        RECT 1166.660 1052.000 1166.920 1052.260 ;
        RECT 1169.880 1052.000 1170.140 1052.260 ;
        RECT 936.200 24.520 936.460 24.780 ;
        RECT 1166.660 24.520 1166.920 24.780 ;
      LAYER met2 ;
        RECT 1171.170 1100.650 1171.450 1104.000 ;
        RECT 1169.940 1100.510 1171.450 1100.650 ;
        RECT 1169.940 1052.290 1170.080 1100.510 ;
        RECT 1171.170 1100.000 1171.450 1100.510 ;
        RECT 1166.660 1051.970 1166.920 1052.290 ;
        RECT 1169.880 1051.970 1170.140 1052.290 ;
        RECT 1166.720 24.810 1166.860 1051.970 ;
        RECT 936.200 24.490 936.460 24.810 ;
        RECT 1166.660 24.490 1166.920 24.810 ;
        RECT 936.260 2.000 936.400 24.490 ;
        RECT 936.050 -4.000 936.610 2.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 954.110 25.060 954.430 25.120 ;
        RECT 1174.450 25.060 1174.770 25.120 ;
        RECT 954.110 24.920 1174.770 25.060 ;
        RECT 954.110 24.860 954.430 24.920 ;
        RECT 1174.450 24.860 1174.770 24.920 ;
      LAYER via ;
        RECT 954.140 24.860 954.400 25.120 ;
        RECT 1174.480 24.860 1174.740 25.120 ;
      LAYER met2 ;
        RECT 1177.150 1100.650 1177.430 1104.000 ;
        RECT 1176.380 1100.510 1177.430 1100.650 ;
        RECT 1176.380 1088.410 1176.520 1100.510 ;
        RECT 1177.150 1100.000 1177.430 1100.510 ;
        RECT 1175.460 1088.270 1176.520 1088.410 ;
        RECT 1175.460 1051.010 1175.600 1088.270 ;
        RECT 1174.540 1050.870 1175.600 1051.010 ;
        RECT 1174.540 25.150 1174.680 1050.870 ;
        RECT 954.140 24.830 954.400 25.150 ;
        RECT 1174.480 24.830 1174.740 25.150 ;
        RECT 954.200 2.000 954.340 24.830 ;
        RECT 953.990 -4.000 954.550 2.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1181.885 800.785 1182.055 855.355 ;
        RECT 1181.425 603.245 1181.595 710.515 ;
        RECT 1181.425 483.225 1181.595 531.335 ;
        RECT 1181.425 379.525 1181.595 434.775 ;
        RECT 1181.885 96.645 1182.055 144.755 ;
      LAYER mcon ;
        RECT 1181.885 855.185 1182.055 855.355 ;
        RECT 1181.425 710.345 1181.595 710.515 ;
        RECT 1181.425 531.165 1181.595 531.335 ;
        RECT 1181.425 434.605 1181.595 434.775 ;
        RECT 1181.885 144.585 1182.055 144.755 ;
      LAYER met1 ;
        RECT 1181.350 1062.740 1181.670 1062.800 ;
        RECT 1183.650 1062.740 1183.970 1062.800 ;
        RECT 1181.350 1062.600 1183.970 1062.740 ;
        RECT 1181.350 1062.540 1181.670 1062.600 ;
        RECT 1183.650 1062.540 1183.970 1062.600 ;
        RECT 1181.350 1028.060 1181.670 1028.120 ;
        RECT 1182.270 1028.060 1182.590 1028.120 ;
        RECT 1181.350 1027.920 1182.590 1028.060 ;
        RECT 1181.350 1027.860 1181.670 1027.920 ;
        RECT 1182.270 1027.860 1182.590 1027.920 ;
        RECT 1181.350 910.760 1181.670 910.820 ;
        RECT 1182.270 910.760 1182.590 910.820 ;
        RECT 1181.350 910.620 1182.590 910.760 ;
        RECT 1181.350 910.560 1181.670 910.620 ;
        RECT 1182.270 910.560 1182.590 910.620 ;
        RECT 1181.810 855.340 1182.130 855.400 ;
        RECT 1181.615 855.200 1182.130 855.340 ;
        RECT 1181.810 855.140 1182.130 855.200 ;
        RECT 1181.825 800.940 1182.115 800.985 ;
        RECT 1181.440 800.800 1182.115 800.940 ;
        RECT 1181.440 800.660 1181.580 800.800 ;
        RECT 1181.825 800.755 1182.115 800.800 ;
        RECT 1181.350 800.400 1181.670 800.660 ;
        RECT 1180.890 711.180 1181.210 711.240 ;
        RECT 1181.350 711.180 1181.670 711.240 ;
        RECT 1180.890 711.040 1181.670 711.180 ;
        RECT 1180.890 710.980 1181.210 711.040 ;
        RECT 1181.350 710.980 1181.670 711.040 ;
        RECT 1180.890 710.500 1181.210 710.560 ;
        RECT 1181.365 710.500 1181.655 710.545 ;
        RECT 1180.890 710.360 1181.655 710.500 ;
        RECT 1180.890 710.300 1181.210 710.360 ;
        RECT 1181.365 710.315 1181.655 710.360 ;
        RECT 1181.350 603.400 1181.670 603.460 ;
        RECT 1181.155 603.260 1181.670 603.400 ;
        RECT 1181.350 603.200 1181.670 603.260 ;
        RECT 1181.810 545.600 1182.130 545.660 ;
        RECT 1181.440 545.460 1182.130 545.600 ;
        RECT 1181.440 544.980 1181.580 545.460 ;
        RECT 1181.810 545.400 1182.130 545.460 ;
        RECT 1181.350 544.720 1181.670 544.980 ;
        RECT 1181.350 531.320 1181.670 531.380 ;
        RECT 1181.155 531.180 1181.670 531.320 ;
        RECT 1181.350 531.120 1181.670 531.180 ;
        RECT 1181.365 483.380 1181.655 483.425 ;
        RECT 1181.810 483.380 1182.130 483.440 ;
        RECT 1181.365 483.240 1182.130 483.380 ;
        RECT 1181.365 483.195 1181.655 483.240 ;
        RECT 1181.810 483.180 1182.130 483.240 ;
        RECT 1181.810 448.840 1182.130 449.100 ;
        RECT 1181.900 448.420 1182.040 448.840 ;
        RECT 1181.810 448.160 1182.130 448.420 ;
        RECT 1181.350 434.760 1181.670 434.820 ;
        RECT 1181.155 434.620 1181.670 434.760 ;
        RECT 1181.350 434.560 1181.670 434.620 ;
        RECT 1181.365 379.680 1181.655 379.725 ;
        RECT 1182.270 379.680 1182.590 379.740 ;
        RECT 1181.365 379.540 1182.590 379.680 ;
        RECT 1181.365 379.495 1181.655 379.540 ;
        RECT 1182.270 379.480 1182.590 379.540 ;
        RECT 1181.350 338.200 1181.670 338.260 ;
        RECT 1182.270 338.200 1182.590 338.260 ;
        RECT 1181.350 338.060 1182.590 338.200 ;
        RECT 1181.350 338.000 1181.670 338.060 ;
        RECT 1182.270 338.000 1182.590 338.060 ;
        RECT 1181.350 207.100 1181.670 207.360 ;
        RECT 1181.440 206.680 1181.580 207.100 ;
        RECT 1181.350 206.420 1181.670 206.680 ;
        RECT 1181.810 144.740 1182.130 144.800 ;
        RECT 1181.615 144.600 1182.130 144.740 ;
        RECT 1181.810 144.540 1182.130 144.600 ;
        RECT 1181.810 96.800 1182.130 96.860 ;
        RECT 1181.615 96.660 1182.130 96.800 ;
        RECT 1181.810 96.600 1182.130 96.660 ;
        RECT 972.050 25.400 972.370 25.460 ;
        RECT 1181.810 25.400 1182.130 25.460 ;
        RECT 972.050 25.260 1182.130 25.400 ;
        RECT 972.050 25.200 972.370 25.260 ;
        RECT 1181.810 25.200 1182.130 25.260 ;
      LAYER via ;
        RECT 1181.380 1062.540 1181.640 1062.800 ;
        RECT 1183.680 1062.540 1183.940 1062.800 ;
        RECT 1181.380 1027.860 1181.640 1028.120 ;
        RECT 1182.300 1027.860 1182.560 1028.120 ;
        RECT 1181.380 910.560 1181.640 910.820 ;
        RECT 1182.300 910.560 1182.560 910.820 ;
        RECT 1181.840 855.140 1182.100 855.400 ;
        RECT 1181.380 800.400 1181.640 800.660 ;
        RECT 1180.920 710.980 1181.180 711.240 ;
        RECT 1181.380 710.980 1181.640 711.240 ;
        RECT 1180.920 710.300 1181.180 710.560 ;
        RECT 1181.380 603.200 1181.640 603.460 ;
        RECT 1181.840 545.400 1182.100 545.660 ;
        RECT 1181.380 544.720 1181.640 544.980 ;
        RECT 1181.380 531.120 1181.640 531.380 ;
        RECT 1181.840 483.180 1182.100 483.440 ;
        RECT 1181.840 448.840 1182.100 449.100 ;
        RECT 1181.840 448.160 1182.100 448.420 ;
        RECT 1181.380 434.560 1181.640 434.820 ;
        RECT 1182.300 379.480 1182.560 379.740 ;
        RECT 1181.380 338.000 1181.640 338.260 ;
        RECT 1182.300 338.000 1182.560 338.260 ;
        RECT 1181.380 207.100 1181.640 207.360 ;
        RECT 1181.380 206.420 1181.640 206.680 ;
        RECT 1181.840 144.540 1182.100 144.800 ;
        RECT 1181.840 96.600 1182.100 96.860 ;
        RECT 972.080 25.200 972.340 25.460 ;
        RECT 1181.840 25.200 1182.100 25.460 ;
      LAYER met2 ;
        RECT 1183.590 1100.580 1183.870 1104.000 ;
        RECT 1183.590 1100.000 1183.880 1100.580 ;
        RECT 1183.740 1062.830 1183.880 1100.000 ;
        RECT 1181.380 1062.510 1181.640 1062.830 ;
        RECT 1183.680 1062.510 1183.940 1062.830 ;
        RECT 1181.440 1028.150 1181.580 1062.510 ;
        RECT 1181.380 1027.830 1181.640 1028.150 ;
        RECT 1182.300 1027.830 1182.560 1028.150 ;
        RECT 1182.360 989.130 1182.500 1027.830 ;
        RECT 1181.900 988.990 1182.500 989.130 ;
        RECT 1181.900 931.330 1182.040 988.990 ;
        RECT 1181.440 931.190 1182.040 931.330 ;
        RECT 1181.440 910.850 1181.580 931.190 ;
        RECT 1181.380 910.530 1181.640 910.850 ;
        RECT 1182.300 910.530 1182.560 910.850 ;
        RECT 1182.360 862.650 1182.500 910.530 ;
        RECT 1181.900 862.510 1182.500 862.650 ;
        RECT 1181.900 855.430 1182.040 862.510 ;
        RECT 1181.840 855.110 1182.100 855.430 ;
        RECT 1181.380 800.370 1181.640 800.690 ;
        RECT 1181.440 711.270 1181.580 800.370 ;
        RECT 1180.920 710.950 1181.180 711.270 ;
        RECT 1181.380 710.950 1181.640 711.270 ;
        RECT 1180.980 710.590 1181.120 710.950 ;
        RECT 1180.920 710.270 1181.180 710.590 ;
        RECT 1181.380 603.170 1181.640 603.490 ;
        RECT 1181.440 579.770 1181.580 603.170 ;
        RECT 1181.440 579.630 1182.040 579.770 ;
        RECT 1181.900 545.690 1182.040 579.630 ;
        RECT 1181.840 545.370 1182.100 545.690 ;
        RECT 1181.380 544.690 1181.640 545.010 ;
        RECT 1181.440 531.410 1181.580 544.690 ;
        RECT 1181.380 531.090 1181.640 531.410 ;
        RECT 1181.840 483.150 1182.100 483.470 ;
        RECT 1181.900 449.130 1182.040 483.150 ;
        RECT 1181.840 448.810 1182.100 449.130 ;
        RECT 1181.840 448.130 1182.100 448.450 ;
        RECT 1181.900 434.930 1182.040 448.130 ;
        RECT 1181.440 434.850 1182.040 434.930 ;
        RECT 1181.380 434.790 1182.040 434.850 ;
        RECT 1181.380 434.530 1181.640 434.790 ;
        RECT 1182.300 379.450 1182.560 379.770 ;
        RECT 1182.360 338.290 1182.500 379.450 ;
        RECT 1181.380 337.970 1181.640 338.290 ;
        RECT 1182.300 337.970 1182.560 338.290 ;
        RECT 1181.440 307.770 1181.580 337.970 ;
        RECT 1181.440 307.630 1182.500 307.770 ;
        RECT 1182.360 303.520 1182.500 307.630 ;
        RECT 1181.900 303.380 1182.500 303.520 ;
        RECT 1181.900 242.605 1182.040 303.380 ;
        RECT 1181.830 242.235 1182.110 242.605 ;
        RECT 1181.370 241.555 1181.650 241.925 ;
        RECT 1181.440 207.390 1181.580 241.555 ;
        RECT 1181.380 207.070 1181.640 207.390 ;
        RECT 1181.380 206.390 1181.640 206.710 ;
        RECT 1181.440 158.170 1181.580 206.390 ;
        RECT 1181.440 158.030 1182.040 158.170 ;
        RECT 1181.900 144.830 1182.040 158.030 ;
        RECT 1181.840 144.510 1182.100 144.830 ;
        RECT 1181.840 96.570 1182.100 96.890 ;
        RECT 1181.900 25.490 1182.040 96.570 ;
        RECT 972.080 25.170 972.340 25.490 ;
        RECT 1181.840 25.170 1182.100 25.490 ;
        RECT 972.140 2.000 972.280 25.170 ;
        RECT 971.930 -4.000 972.490 2.000 ;
      LAYER via2 ;
        RECT 1181.830 242.280 1182.110 242.560 ;
        RECT 1181.370 241.600 1181.650 241.880 ;
      LAYER met3 ;
        RECT 1181.805 242.570 1182.135 242.585 ;
        RECT 1180.670 242.270 1182.135 242.570 ;
        RECT 1180.670 241.890 1180.970 242.270 ;
        RECT 1181.805 242.255 1182.135 242.270 ;
        RECT 1181.345 241.890 1181.675 241.905 ;
        RECT 1180.670 241.590 1181.675 241.890 ;
        RECT 1181.345 241.575 1181.675 241.590 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1071.485 48.365 1071.655 96.475 ;
      LAYER mcon ;
        RECT 1071.485 96.305 1071.655 96.475 ;
      LAYER met1 ;
        RECT 1070.490 110.400 1070.810 110.460 ;
        RECT 1071.410 110.400 1071.730 110.460 ;
        RECT 1070.490 110.260 1071.730 110.400 ;
        RECT 1070.490 110.200 1070.810 110.260 ;
        RECT 1071.410 110.200 1071.730 110.260 ;
        RECT 1071.410 96.460 1071.730 96.520 ;
        RECT 1071.215 96.320 1071.730 96.460 ;
        RECT 1071.410 96.260 1071.730 96.320 ;
        RECT 1071.410 48.520 1071.730 48.580 ;
        RECT 1071.215 48.380 1071.730 48.520 ;
        RECT 1071.410 48.320 1071.730 48.380 ;
        RECT 650.970 46.480 651.290 46.540 ;
        RECT 1071.410 46.480 1071.730 46.540 ;
        RECT 650.970 46.340 1071.730 46.480 ;
        RECT 650.970 46.280 651.290 46.340 ;
        RECT 1071.410 46.280 1071.730 46.340 ;
      LAYER via ;
        RECT 1070.520 110.200 1070.780 110.460 ;
        RECT 1071.440 110.200 1071.700 110.460 ;
        RECT 1071.440 96.260 1071.700 96.520 ;
        RECT 1071.440 48.320 1071.700 48.580 ;
        RECT 651.000 46.280 651.260 46.540 ;
        RECT 1071.440 46.280 1071.700 46.540 ;
      LAYER met2 ;
        RECT 1073.190 1100.650 1073.470 1104.000 ;
        RECT 1072.420 1100.510 1073.470 1100.650 ;
        RECT 1072.420 1088.410 1072.560 1100.510 ;
        RECT 1073.190 1100.000 1073.470 1100.510 ;
        RECT 1070.580 1088.270 1072.560 1088.410 ;
        RECT 1070.580 110.490 1070.720 1088.270 ;
        RECT 1070.520 110.170 1070.780 110.490 ;
        RECT 1071.440 110.170 1071.700 110.490 ;
        RECT 1071.500 96.550 1071.640 110.170 ;
        RECT 1071.440 96.230 1071.700 96.550 ;
        RECT 1071.440 48.290 1071.700 48.610 ;
        RECT 1071.500 46.570 1071.640 48.290 ;
        RECT 651.000 46.250 651.260 46.570 ;
        RECT 1071.440 46.250 1071.700 46.570 ;
        RECT 651.060 2.000 651.200 46.250 ;
        RECT 650.850 -4.000 651.410 2.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 989.990 25.740 990.310 25.800 ;
        RECT 1188.250 25.740 1188.570 25.800 ;
        RECT 989.990 25.600 1188.570 25.740 ;
        RECT 989.990 25.540 990.310 25.600 ;
        RECT 1188.250 25.540 1188.570 25.600 ;
      LAYER via ;
        RECT 990.020 25.540 990.280 25.800 ;
        RECT 1188.280 25.540 1188.540 25.800 ;
      LAYER met2 ;
        RECT 1189.570 1100.650 1189.850 1104.000 ;
        RECT 1188.340 1100.510 1189.850 1100.650 ;
        RECT 1188.340 25.830 1188.480 1100.510 ;
        RECT 1189.570 1100.000 1189.850 1100.510 ;
        RECT 990.020 25.510 990.280 25.830 ;
        RECT 1188.280 25.510 1188.540 25.830 ;
        RECT 990.080 2.000 990.220 25.510 ;
        RECT 989.870 -4.000 990.430 2.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1007.470 26.080 1007.790 26.140 ;
        RECT 1194.690 26.080 1195.010 26.140 ;
        RECT 1007.470 25.940 1195.010 26.080 ;
        RECT 1007.470 25.880 1007.790 25.940 ;
        RECT 1194.690 25.880 1195.010 25.940 ;
      LAYER via ;
        RECT 1007.500 25.880 1007.760 26.140 ;
        RECT 1194.720 25.880 1194.980 26.140 ;
      LAYER met2 ;
        RECT 1195.550 1100.650 1195.830 1104.000 ;
        RECT 1194.780 1100.510 1195.830 1100.650 ;
        RECT 1194.780 26.170 1194.920 1100.510 ;
        RECT 1195.550 1100.000 1195.830 1100.510 ;
        RECT 1007.500 25.850 1007.760 26.170 ;
        RECT 1194.720 25.850 1194.980 26.170 ;
        RECT 1007.560 2.000 1007.700 25.850 ;
        RECT 1007.350 -4.000 1007.910 2.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1025.410 26.420 1025.730 26.480 ;
        RECT 1201.590 26.420 1201.910 26.480 ;
        RECT 1025.410 26.280 1201.910 26.420 ;
        RECT 1025.410 26.220 1025.730 26.280 ;
        RECT 1201.590 26.220 1201.910 26.280 ;
      LAYER via ;
        RECT 1025.440 26.220 1025.700 26.480 ;
        RECT 1201.620 26.220 1201.880 26.480 ;
      LAYER met2 ;
        RECT 1201.990 1100.650 1202.270 1104.000 ;
        RECT 1201.680 1100.510 1202.270 1100.650 ;
        RECT 1201.680 26.510 1201.820 1100.510 ;
        RECT 1201.990 1100.000 1202.270 1100.510 ;
        RECT 1025.440 26.190 1025.700 26.510 ;
        RECT 1201.620 26.190 1201.880 26.510 ;
        RECT 1025.500 2.000 1025.640 26.190 ;
        RECT 1025.290 -4.000 1025.850 2.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1043.350 26.760 1043.670 26.820 ;
        RECT 1208.490 26.760 1208.810 26.820 ;
        RECT 1043.350 26.620 1208.810 26.760 ;
        RECT 1043.350 26.560 1043.670 26.620 ;
        RECT 1208.490 26.560 1208.810 26.620 ;
      LAYER via ;
        RECT 1043.380 26.560 1043.640 26.820 ;
        RECT 1208.520 26.560 1208.780 26.820 ;
      LAYER met2 ;
        RECT 1207.970 1100.650 1208.250 1104.000 ;
        RECT 1207.970 1100.510 1208.720 1100.650 ;
        RECT 1207.970 1100.000 1208.250 1100.510 ;
        RECT 1208.580 26.850 1208.720 1100.510 ;
        RECT 1043.380 26.530 1043.640 26.850 ;
        RECT 1208.520 26.530 1208.780 26.850 ;
        RECT 1043.440 2.000 1043.580 26.530 ;
        RECT 1043.230 -4.000 1043.790 2.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1061.825 1062.585 1061.995 1088.595 ;
        RECT 1062.285 772.905 1062.455 821.015 ;
        RECT 1061.365 655.605 1061.535 703.715 ;
        RECT 1061.365 565.505 1061.535 607.155 ;
        RECT 1062.285 186.405 1062.455 241.315 ;
        RECT 1061.365 96.305 1061.535 137.955 ;
        RECT 1061.365 48.365 1061.535 62.815 ;
      LAYER mcon ;
        RECT 1061.825 1088.425 1061.995 1088.595 ;
        RECT 1062.285 820.845 1062.455 821.015 ;
        RECT 1061.365 703.545 1061.535 703.715 ;
        RECT 1061.365 606.985 1061.535 607.155 ;
        RECT 1062.285 241.145 1062.455 241.315 ;
        RECT 1061.365 137.785 1061.535 137.955 ;
        RECT 1061.365 62.645 1061.535 62.815 ;
      LAYER met1 ;
        RECT 1061.765 1088.580 1062.055 1088.625 ;
        RECT 1214.010 1088.580 1214.330 1088.640 ;
        RECT 1061.765 1088.440 1214.330 1088.580 ;
        RECT 1061.765 1088.395 1062.055 1088.440 ;
        RECT 1214.010 1088.380 1214.330 1088.440 ;
        RECT 1061.750 1062.740 1062.070 1062.800 ;
        RECT 1061.555 1062.600 1062.070 1062.740 ;
        RECT 1061.750 1062.540 1062.070 1062.600 ;
        RECT 1060.830 1014.460 1061.150 1014.520 ;
        RECT 1062.210 1014.460 1062.530 1014.520 ;
        RECT 1060.830 1014.320 1062.530 1014.460 ;
        RECT 1060.830 1014.260 1061.150 1014.320 ;
        RECT 1062.210 1014.260 1062.530 1014.320 ;
        RECT 1062.210 821.000 1062.530 821.060 ;
        RECT 1062.015 820.860 1062.530 821.000 ;
        RECT 1062.210 820.800 1062.530 820.860 ;
        RECT 1062.210 773.060 1062.530 773.120 ;
        RECT 1062.015 772.920 1062.530 773.060 ;
        RECT 1062.210 772.860 1062.530 772.920 ;
        RECT 1061.305 703.700 1061.595 703.745 ;
        RECT 1061.750 703.700 1062.070 703.760 ;
        RECT 1061.305 703.560 1062.070 703.700 ;
        RECT 1061.305 703.515 1061.595 703.560 ;
        RECT 1061.750 703.500 1062.070 703.560 ;
        RECT 1061.305 655.760 1061.595 655.805 ;
        RECT 1061.750 655.760 1062.070 655.820 ;
        RECT 1061.305 655.620 1062.070 655.760 ;
        RECT 1061.305 655.575 1061.595 655.620 ;
        RECT 1061.750 655.560 1062.070 655.620 ;
        RECT 1061.305 607.140 1061.595 607.185 ;
        RECT 1061.750 607.140 1062.070 607.200 ;
        RECT 1061.305 607.000 1062.070 607.140 ;
        RECT 1061.305 606.955 1061.595 607.000 ;
        RECT 1061.750 606.940 1062.070 607.000 ;
        RECT 1061.305 565.660 1061.595 565.705 ;
        RECT 1061.750 565.660 1062.070 565.720 ;
        RECT 1061.305 565.520 1062.070 565.660 ;
        RECT 1061.305 565.475 1061.595 565.520 ;
        RECT 1061.750 565.460 1062.070 565.520 ;
        RECT 1061.290 427.620 1061.610 427.680 ;
        RECT 1062.210 427.620 1062.530 427.680 ;
        RECT 1061.290 427.480 1062.530 427.620 ;
        RECT 1061.290 427.420 1061.610 427.480 ;
        RECT 1062.210 427.420 1062.530 427.480 ;
        RECT 1061.290 331.060 1061.610 331.120 ;
        RECT 1061.750 331.060 1062.070 331.120 ;
        RECT 1061.290 330.920 1062.070 331.060 ;
        RECT 1061.290 330.860 1061.610 330.920 ;
        RECT 1061.750 330.860 1062.070 330.920 ;
        RECT 1062.210 241.300 1062.530 241.360 ;
        RECT 1062.015 241.160 1062.530 241.300 ;
        RECT 1062.210 241.100 1062.530 241.160 ;
        RECT 1061.750 186.560 1062.070 186.620 ;
        RECT 1062.225 186.560 1062.515 186.605 ;
        RECT 1061.750 186.420 1062.515 186.560 ;
        RECT 1061.750 186.360 1062.070 186.420 ;
        RECT 1062.225 186.375 1062.515 186.420 ;
        RECT 1061.290 137.940 1061.610 138.000 ;
        RECT 1061.290 137.800 1061.805 137.940 ;
        RECT 1061.290 137.740 1061.610 137.800 ;
        RECT 1061.290 96.460 1061.610 96.520 ;
        RECT 1061.095 96.320 1061.610 96.460 ;
        RECT 1061.290 96.260 1061.610 96.320 ;
        RECT 1061.290 62.800 1061.610 62.860 ;
        RECT 1061.095 62.660 1061.610 62.800 ;
        RECT 1061.290 62.600 1061.610 62.660 ;
        RECT 1061.290 48.520 1061.610 48.580 ;
        RECT 1061.095 48.380 1061.610 48.520 ;
        RECT 1061.290 48.320 1061.610 48.380 ;
      LAYER via ;
        RECT 1214.040 1088.380 1214.300 1088.640 ;
        RECT 1061.780 1062.540 1062.040 1062.800 ;
        RECT 1060.860 1014.260 1061.120 1014.520 ;
        RECT 1062.240 1014.260 1062.500 1014.520 ;
        RECT 1062.240 820.800 1062.500 821.060 ;
        RECT 1062.240 772.860 1062.500 773.120 ;
        RECT 1061.780 703.500 1062.040 703.760 ;
        RECT 1061.780 655.560 1062.040 655.820 ;
        RECT 1061.780 606.940 1062.040 607.200 ;
        RECT 1061.780 565.460 1062.040 565.720 ;
        RECT 1061.320 427.420 1061.580 427.680 ;
        RECT 1062.240 427.420 1062.500 427.680 ;
        RECT 1061.320 330.860 1061.580 331.120 ;
        RECT 1061.780 330.860 1062.040 331.120 ;
        RECT 1062.240 241.100 1062.500 241.360 ;
        RECT 1061.780 186.360 1062.040 186.620 ;
        RECT 1061.320 137.740 1061.580 138.000 ;
        RECT 1061.320 96.260 1061.580 96.520 ;
        RECT 1061.320 62.600 1061.580 62.860 ;
        RECT 1061.320 48.320 1061.580 48.580 ;
      LAYER met2 ;
        RECT 1213.950 1100.580 1214.230 1104.000 ;
        RECT 1213.950 1100.000 1214.240 1100.580 ;
        RECT 1214.100 1088.670 1214.240 1100.000 ;
        RECT 1214.040 1088.350 1214.300 1088.670 ;
        RECT 1061.780 1062.685 1062.040 1062.830 ;
        RECT 1060.850 1062.315 1061.130 1062.685 ;
        RECT 1061.770 1062.315 1062.050 1062.685 ;
        RECT 1060.920 1014.550 1061.060 1062.315 ;
        RECT 1060.860 1014.230 1061.120 1014.550 ;
        RECT 1062.240 1014.230 1062.500 1014.550 ;
        RECT 1062.300 821.090 1062.440 1014.230 ;
        RECT 1062.240 820.770 1062.500 821.090 ;
        RECT 1062.240 772.830 1062.500 773.150 ;
        RECT 1062.300 748.410 1062.440 772.830 ;
        RECT 1061.840 748.270 1062.440 748.410 ;
        RECT 1061.840 703.790 1061.980 748.270 ;
        RECT 1061.780 703.470 1062.040 703.790 ;
        RECT 1061.780 655.530 1062.040 655.850 ;
        RECT 1061.840 607.230 1061.980 655.530 ;
        RECT 1061.780 606.910 1062.040 607.230 ;
        RECT 1061.780 565.430 1062.040 565.750 ;
        RECT 1061.840 541.690 1061.980 565.430 ;
        RECT 1061.380 541.550 1061.980 541.690 ;
        RECT 1061.380 451.930 1061.520 541.550 ;
        RECT 1061.380 451.790 1062.440 451.930 ;
        RECT 1062.300 427.710 1062.440 451.790 ;
        RECT 1061.320 427.390 1061.580 427.710 ;
        RECT 1062.240 427.390 1062.500 427.710 ;
        RECT 1061.380 331.150 1061.520 427.390 ;
        RECT 1061.320 330.830 1061.580 331.150 ;
        RECT 1061.780 330.830 1062.040 331.150 ;
        RECT 1061.840 241.810 1061.980 330.830 ;
        RECT 1061.840 241.670 1062.440 241.810 ;
        RECT 1062.300 241.390 1062.440 241.670 ;
        RECT 1062.240 241.070 1062.500 241.390 ;
        RECT 1061.780 186.330 1062.040 186.650 ;
        RECT 1061.840 138.450 1061.980 186.330 ;
        RECT 1061.380 138.310 1061.980 138.450 ;
        RECT 1061.380 138.030 1061.520 138.310 ;
        RECT 1061.320 137.710 1061.580 138.030 ;
        RECT 1061.320 96.230 1061.580 96.550 ;
        RECT 1061.380 62.890 1061.520 96.230 ;
        RECT 1061.320 62.570 1061.580 62.890 ;
        RECT 1061.320 48.290 1061.580 48.610 ;
        RECT 1061.380 2.000 1061.520 48.290 ;
        RECT 1061.170 -4.000 1061.730 2.000 ;
      LAYER via2 ;
        RECT 1060.850 1062.360 1061.130 1062.640 ;
        RECT 1061.770 1062.360 1062.050 1062.640 ;
      LAYER met3 ;
        RECT 1060.825 1062.650 1061.155 1062.665 ;
        RECT 1061.745 1062.650 1062.075 1062.665 ;
        RECT 1060.825 1062.350 1062.075 1062.650 ;
        RECT 1060.825 1062.335 1061.155 1062.350 ;
        RECT 1061.745 1062.335 1062.075 1062.350 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1193.845 19.125 1194.015 20.315 ;
      LAYER mcon ;
        RECT 1193.845 20.145 1194.015 20.315 ;
      LAYER met1 ;
        RECT 1214.930 1052.200 1215.250 1052.260 ;
        RECT 1219.070 1052.200 1219.390 1052.260 ;
        RECT 1214.930 1052.060 1219.390 1052.200 ;
        RECT 1214.930 1052.000 1215.250 1052.060 ;
        RECT 1219.070 1052.000 1219.390 1052.060 ;
        RECT 1079.230 20.300 1079.550 20.360 ;
        RECT 1193.785 20.300 1194.075 20.345 ;
        RECT 1079.230 20.160 1194.075 20.300 ;
        RECT 1079.230 20.100 1079.550 20.160 ;
        RECT 1193.785 20.115 1194.075 20.160 ;
        RECT 1193.785 19.280 1194.075 19.325 ;
        RECT 1214.930 19.280 1215.250 19.340 ;
        RECT 1193.785 19.140 1215.250 19.280 ;
        RECT 1193.785 19.095 1194.075 19.140 ;
        RECT 1214.930 19.080 1215.250 19.140 ;
      LAYER via ;
        RECT 1214.960 1052.000 1215.220 1052.260 ;
        RECT 1219.100 1052.000 1219.360 1052.260 ;
        RECT 1079.260 20.100 1079.520 20.360 ;
        RECT 1214.960 19.080 1215.220 19.340 ;
      LAYER met2 ;
        RECT 1220.390 1100.650 1220.670 1104.000 ;
        RECT 1219.160 1100.510 1220.670 1100.650 ;
        RECT 1219.160 1052.290 1219.300 1100.510 ;
        RECT 1220.390 1100.000 1220.670 1100.510 ;
        RECT 1214.960 1051.970 1215.220 1052.290 ;
        RECT 1219.100 1051.970 1219.360 1052.290 ;
        RECT 1079.260 20.070 1079.520 20.390 ;
        RECT 1079.320 2.000 1079.460 20.070 ;
        RECT 1215.020 19.370 1215.160 1051.970 ;
        RECT 1214.960 19.050 1215.220 19.370 ;
        RECT 1079.110 -4.000 1079.670 2.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1096.710 1086.200 1097.030 1086.260 ;
        RECT 1226.430 1086.200 1226.750 1086.260 ;
        RECT 1096.710 1086.060 1226.750 1086.200 ;
        RECT 1096.710 1086.000 1097.030 1086.060 ;
        RECT 1226.430 1086.000 1226.750 1086.060 ;
      LAYER via ;
        RECT 1096.740 1086.000 1097.000 1086.260 ;
        RECT 1226.460 1086.000 1226.720 1086.260 ;
      LAYER met2 ;
        RECT 1226.370 1100.580 1226.650 1104.000 ;
        RECT 1226.370 1100.000 1226.660 1100.580 ;
        RECT 1226.520 1086.290 1226.660 1100.000 ;
        RECT 1096.740 1085.970 1097.000 1086.290 ;
        RECT 1226.460 1085.970 1226.720 1086.290 ;
        RECT 1096.800 2.000 1096.940 1085.970 ;
        RECT 1096.590 -4.000 1097.150 2.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1148.690 1084.840 1149.010 1084.900 ;
        RECT 1232.410 1084.840 1232.730 1084.900 ;
        RECT 1148.690 1084.700 1232.730 1084.840 ;
        RECT 1148.690 1084.640 1149.010 1084.700 ;
        RECT 1232.410 1084.640 1232.730 1084.700 ;
        RECT 1114.650 15.200 1114.970 15.260 ;
        RECT 1148.690 15.200 1149.010 15.260 ;
        RECT 1114.650 15.060 1149.010 15.200 ;
        RECT 1114.650 15.000 1114.970 15.060 ;
        RECT 1148.690 15.000 1149.010 15.060 ;
      LAYER via ;
        RECT 1148.720 1084.640 1148.980 1084.900 ;
        RECT 1232.440 1084.640 1232.700 1084.900 ;
        RECT 1114.680 15.000 1114.940 15.260 ;
        RECT 1148.720 15.000 1148.980 15.260 ;
      LAYER met2 ;
        RECT 1232.350 1100.580 1232.630 1104.000 ;
        RECT 1232.350 1100.000 1232.640 1100.580 ;
        RECT 1232.500 1084.930 1232.640 1100.000 ;
        RECT 1148.720 1084.610 1148.980 1084.930 ;
        RECT 1232.440 1084.610 1232.700 1084.930 ;
        RECT 1148.780 15.290 1148.920 1084.610 ;
        RECT 1114.680 14.970 1114.940 15.290 ;
        RECT 1148.720 14.970 1148.980 15.290 ;
        RECT 1114.740 2.000 1114.880 14.970 ;
        RECT 1114.530 -4.000 1115.090 2.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1138.110 1085.520 1138.430 1085.580 ;
        RECT 1238.390 1085.520 1238.710 1085.580 ;
        RECT 1138.110 1085.380 1238.710 1085.520 ;
        RECT 1138.110 1085.320 1138.430 1085.380 ;
        RECT 1238.390 1085.320 1238.710 1085.380 ;
        RECT 1132.590 17.240 1132.910 17.300 ;
        RECT 1138.110 17.240 1138.430 17.300 ;
        RECT 1132.590 17.100 1138.430 17.240 ;
        RECT 1132.590 17.040 1132.910 17.100 ;
        RECT 1138.110 17.040 1138.430 17.100 ;
      LAYER via ;
        RECT 1138.140 1085.320 1138.400 1085.580 ;
        RECT 1238.420 1085.320 1238.680 1085.580 ;
        RECT 1132.620 17.040 1132.880 17.300 ;
        RECT 1138.140 17.040 1138.400 17.300 ;
      LAYER met2 ;
        RECT 1238.330 1100.580 1238.610 1104.000 ;
        RECT 1238.330 1100.000 1238.620 1100.580 ;
        RECT 1238.480 1085.610 1238.620 1100.000 ;
        RECT 1138.140 1085.290 1138.400 1085.610 ;
        RECT 1238.420 1085.290 1238.680 1085.610 ;
        RECT 1138.200 17.330 1138.340 1085.290 ;
        RECT 1132.620 17.010 1132.880 17.330 ;
        RECT 1138.140 17.010 1138.400 17.330 ;
        RECT 1132.680 2.000 1132.820 17.010 ;
        RECT 1132.470 -4.000 1133.030 2.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1151.910 1085.180 1152.230 1085.240 ;
        RECT 1244.830 1085.180 1245.150 1085.240 ;
        RECT 1151.910 1085.040 1245.150 1085.180 ;
        RECT 1151.910 1084.980 1152.230 1085.040 ;
        RECT 1244.830 1084.980 1245.150 1085.040 ;
      LAYER via ;
        RECT 1151.940 1084.980 1152.200 1085.240 ;
        RECT 1244.860 1084.980 1245.120 1085.240 ;
      LAYER met2 ;
        RECT 1244.770 1100.580 1245.050 1104.000 ;
        RECT 1244.770 1100.000 1245.060 1100.580 ;
        RECT 1244.920 1085.270 1245.060 1100.000 ;
        RECT 1151.940 1084.950 1152.200 1085.270 ;
        RECT 1244.860 1084.950 1245.120 1085.270 ;
        RECT 1152.000 2.450 1152.140 1084.950 ;
        RECT 1150.620 2.310 1152.140 2.450 ;
        RECT 1150.620 2.000 1150.760 2.310 ;
        RECT 1150.410 -4.000 1150.970 2.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 668.910 46.820 669.230 46.880 ;
        RECT 1077.850 46.820 1078.170 46.880 ;
        RECT 668.910 46.680 1078.170 46.820 ;
        RECT 668.910 46.620 669.230 46.680 ;
        RECT 1077.850 46.620 1078.170 46.680 ;
      LAYER via ;
        RECT 668.940 46.620 669.200 46.880 ;
        RECT 1077.880 46.620 1078.140 46.880 ;
      LAYER met2 ;
        RECT 1079.170 1100.650 1079.450 1104.000 ;
        RECT 1077.940 1100.510 1079.450 1100.650 ;
        RECT 1077.940 46.910 1078.080 1100.510 ;
        RECT 1079.170 1100.000 1079.450 1100.510 ;
        RECT 668.940 46.590 669.200 46.910 ;
        RECT 1077.880 46.590 1078.140 46.910 ;
        RECT 669.000 2.000 669.140 46.590 ;
        RECT 668.790 -4.000 669.350 2.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1203.890 1086.880 1204.210 1086.940 ;
        RECT 1249.430 1086.880 1249.750 1086.940 ;
        RECT 1203.890 1086.740 1249.750 1086.880 ;
        RECT 1203.890 1086.680 1204.210 1086.740 ;
        RECT 1249.430 1086.680 1249.750 1086.740 ;
        RECT 1168.470 19.620 1168.790 19.680 ;
        RECT 1203.430 19.620 1203.750 19.680 ;
        RECT 1168.470 19.480 1203.750 19.620 ;
        RECT 1168.470 19.420 1168.790 19.480 ;
        RECT 1203.430 19.420 1203.750 19.480 ;
      LAYER via ;
        RECT 1203.920 1086.680 1204.180 1086.940 ;
        RECT 1249.460 1086.680 1249.720 1086.940 ;
        RECT 1168.500 19.420 1168.760 19.680 ;
        RECT 1203.460 19.420 1203.720 19.680 ;
      LAYER met2 ;
        RECT 1250.750 1100.650 1251.030 1104.000 ;
        RECT 1249.520 1100.510 1251.030 1100.650 ;
        RECT 1249.520 1086.970 1249.660 1100.510 ;
        RECT 1250.750 1100.000 1251.030 1100.510 ;
        RECT 1203.920 1086.650 1204.180 1086.970 ;
        RECT 1249.460 1086.650 1249.720 1086.970 ;
        RECT 1203.980 20.810 1204.120 1086.650 ;
        RECT 1203.520 20.670 1204.120 20.810 ;
        RECT 1203.520 19.710 1203.660 20.670 ;
        RECT 1168.500 19.390 1168.760 19.710 ;
        RECT 1203.460 19.390 1203.720 19.710 ;
        RECT 1168.560 2.000 1168.700 19.390 ;
        RECT 1168.350 -4.000 1168.910 2.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1186.410 1084.500 1186.730 1084.560 ;
        RECT 1256.790 1084.500 1257.110 1084.560 ;
        RECT 1186.410 1084.360 1257.110 1084.500 ;
        RECT 1186.410 1084.300 1186.730 1084.360 ;
        RECT 1256.790 1084.300 1257.110 1084.360 ;
      LAYER via ;
        RECT 1186.440 1084.300 1186.700 1084.560 ;
        RECT 1256.820 1084.300 1257.080 1084.560 ;
      LAYER met2 ;
        RECT 1256.730 1100.580 1257.010 1104.000 ;
        RECT 1256.730 1100.000 1257.020 1100.580 ;
        RECT 1256.880 1084.590 1257.020 1100.000 ;
        RECT 1186.440 1084.270 1186.700 1084.590 ;
        RECT 1256.820 1084.270 1257.080 1084.590 ;
        RECT 1186.500 2.450 1186.640 1084.270 ;
        RECT 1186.040 2.310 1186.640 2.450 ;
        RECT 1186.040 2.000 1186.180 2.310 ;
        RECT 1185.830 -4.000 1186.390 2.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1207.110 1086.540 1207.430 1086.600 ;
        RECT 1263.230 1086.540 1263.550 1086.600 ;
        RECT 1207.110 1086.400 1263.550 1086.540 ;
        RECT 1207.110 1086.340 1207.430 1086.400 ;
        RECT 1263.230 1086.340 1263.550 1086.400 ;
        RECT 1203.890 20.300 1204.210 20.360 ;
        RECT 1207.110 20.300 1207.430 20.360 ;
        RECT 1203.890 20.160 1207.430 20.300 ;
        RECT 1203.890 20.100 1204.210 20.160 ;
        RECT 1207.110 20.100 1207.430 20.160 ;
      LAYER via ;
        RECT 1207.140 1086.340 1207.400 1086.600 ;
        RECT 1263.260 1086.340 1263.520 1086.600 ;
        RECT 1203.920 20.100 1204.180 20.360 ;
        RECT 1207.140 20.100 1207.400 20.360 ;
      LAYER met2 ;
        RECT 1263.170 1100.580 1263.450 1104.000 ;
        RECT 1263.170 1100.000 1263.460 1100.580 ;
        RECT 1263.320 1086.630 1263.460 1100.000 ;
        RECT 1207.140 1086.310 1207.400 1086.630 ;
        RECT 1263.260 1086.310 1263.520 1086.630 ;
        RECT 1207.200 20.390 1207.340 1086.310 ;
        RECT 1203.920 20.070 1204.180 20.390 ;
        RECT 1207.140 20.070 1207.400 20.390 ;
        RECT 1203.980 2.000 1204.120 20.070 ;
        RECT 1203.770 -4.000 1204.330 2.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1227.810 1087.900 1228.130 1087.960 ;
        RECT 1269.210 1087.900 1269.530 1087.960 ;
        RECT 1227.810 1087.760 1269.530 1087.900 ;
        RECT 1227.810 1087.700 1228.130 1087.760 ;
        RECT 1269.210 1087.700 1269.530 1087.760 ;
        RECT 1221.830 17.920 1222.150 17.980 ;
        RECT 1227.810 17.920 1228.130 17.980 ;
        RECT 1221.830 17.780 1228.130 17.920 ;
        RECT 1221.830 17.720 1222.150 17.780 ;
        RECT 1227.810 17.720 1228.130 17.780 ;
      LAYER via ;
        RECT 1227.840 1087.700 1228.100 1087.960 ;
        RECT 1269.240 1087.700 1269.500 1087.960 ;
        RECT 1221.860 17.720 1222.120 17.980 ;
        RECT 1227.840 17.720 1228.100 17.980 ;
      LAYER met2 ;
        RECT 1269.150 1100.580 1269.430 1104.000 ;
        RECT 1269.150 1100.000 1269.440 1100.580 ;
        RECT 1269.300 1087.990 1269.440 1100.000 ;
        RECT 1227.840 1087.670 1228.100 1087.990 ;
        RECT 1269.240 1087.670 1269.500 1087.990 ;
        RECT 1227.900 18.010 1228.040 1087.670 ;
        RECT 1221.860 17.690 1222.120 18.010 ;
        RECT 1227.840 17.690 1228.100 18.010 ;
        RECT 1221.920 2.000 1222.060 17.690 ;
        RECT 1221.710 -4.000 1222.270 2.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1241.610 1087.560 1241.930 1087.620 ;
        RECT 1275.190 1087.560 1275.510 1087.620 ;
        RECT 1241.610 1087.420 1275.510 1087.560 ;
        RECT 1241.610 1087.360 1241.930 1087.420 ;
        RECT 1275.190 1087.360 1275.510 1087.420 ;
      LAYER via ;
        RECT 1241.640 1087.360 1241.900 1087.620 ;
        RECT 1275.220 1087.360 1275.480 1087.620 ;
      LAYER met2 ;
        RECT 1275.130 1100.580 1275.410 1104.000 ;
        RECT 1275.130 1100.000 1275.420 1100.580 ;
        RECT 1275.280 1087.650 1275.420 1100.000 ;
        RECT 1241.640 1087.330 1241.900 1087.650 ;
        RECT 1275.220 1087.330 1275.480 1087.650 ;
        RECT 1241.700 2.450 1241.840 1087.330 ;
        RECT 1239.860 2.310 1241.840 2.450 ;
        RECT 1239.860 2.000 1240.000 2.310 ;
        RECT 1239.650 -4.000 1240.210 2.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1262.310 1084.840 1262.630 1084.900 ;
        RECT 1281.630 1084.840 1281.950 1084.900 ;
        RECT 1262.310 1084.700 1281.950 1084.840 ;
        RECT 1262.310 1084.640 1262.630 1084.700 ;
        RECT 1281.630 1084.640 1281.950 1084.700 ;
        RECT 1257.250 17.580 1257.570 17.640 ;
        RECT 1262.310 17.580 1262.630 17.640 ;
        RECT 1257.250 17.440 1262.630 17.580 ;
        RECT 1257.250 17.380 1257.570 17.440 ;
        RECT 1262.310 17.380 1262.630 17.440 ;
      LAYER via ;
        RECT 1262.340 1084.640 1262.600 1084.900 ;
        RECT 1281.660 1084.640 1281.920 1084.900 ;
        RECT 1257.280 17.380 1257.540 17.640 ;
        RECT 1262.340 17.380 1262.600 17.640 ;
      LAYER met2 ;
        RECT 1281.570 1100.580 1281.850 1104.000 ;
        RECT 1281.570 1100.000 1281.860 1100.580 ;
        RECT 1281.720 1084.930 1281.860 1100.000 ;
        RECT 1262.340 1084.610 1262.600 1084.930 ;
        RECT 1281.660 1084.610 1281.920 1084.930 ;
        RECT 1262.400 17.670 1262.540 1084.610 ;
        RECT 1257.280 17.350 1257.540 17.670 ;
        RECT 1262.340 17.350 1262.600 17.670 ;
        RECT 1257.340 2.000 1257.480 17.350 ;
        RECT 1257.130 -4.000 1257.690 2.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1276.110 1088.240 1276.430 1088.300 ;
        RECT 1287.610 1088.240 1287.930 1088.300 ;
        RECT 1276.110 1088.100 1287.930 1088.240 ;
        RECT 1276.110 1088.040 1276.430 1088.100 ;
        RECT 1287.610 1088.040 1287.930 1088.100 ;
      LAYER via ;
        RECT 1276.140 1088.040 1276.400 1088.300 ;
        RECT 1287.640 1088.040 1287.900 1088.300 ;
      LAYER met2 ;
        RECT 1287.550 1100.580 1287.830 1104.000 ;
        RECT 1287.550 1100.000 1287.840 1100.580 ;
        RECT 1287.700 1088.330 1287.840 1100.000 ;
        RECT 1276.140 1088.010 1276.400 1088.330 ;
        RECT 1287.640 1088.010 1287.900 1088.330 ;
        RECT 1276.200 2.450 1276.340 1088.010 ;
        RECT 1275.280 2.310 1276.340 2.450 ;
        RECT 1275.280 2.000 1275.420 2.310 ;
        RECT 1275.070 -4.000 1275.630 2.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1291.365 1014.305 1291.535 1038.615 ;
        RECT 1291.365 786.505 1291.535 821.015 ;
        RECT 1291.365 689.605 1291.535 724.455 ;
        RECT 1291.365 593.045 1291.535 627.895 ;
        RECT 1291.365 496.485 1291.535 531.335 ;
        RECT 1291.365 386.325 1291.535 434.775 ;
        RECT 1291.365 158.525 1291.535 193.035 ;
      LAYER mcon ;
        RECT 1291.365 1038.445 1291.535 1038.615 ;
        RECT 1291.365 820.845 1291.535 821.015 ;
        RECT 1291.365 724.285 1291.535 724.455 ;
        RECT 1291.365 627.725 1291.535 627.895 ;
        RECT 1291.365 531.165 1291.535 531.335 ;
        RECT 1291.365 434.605 1291.535 434.775 ;
        RECT 1291.365 192.865 1291.535 193.035 ;
      LAYER met1 ;
        RECT 1291.290 1038.600 1291.610 1038.660 ;
        RECT 1291.095 1038.460 1291.610 1038.600 ;
        RECT 1291.290 1038.400 1291.610 1038.460 ;
        RECT 1291.305 1014.460 1291.595 1014.505 ;
        RECT 1291.750 1014.460 1292.070 1014.520 ;
        RECT 1291.305 1014.320 1292.070 1014.460 ;
        RECT 1291.305 1014.275 1291.595 1014.320 ;
        RECT 1291.750 1014.260 1292.070 1014.320 ;
        RECT 1290.830 835.280 1291.150 835.340 ;
        RECT 1291.750 835.280 1292.070 835.340 ;
        RECT 1290.830 835.140 1292.070 835.280 ;
        RECT 1290.830 835.080 1291.150 835.140 ;
        RECT 1291.750 835.080 1292.070 835.140 ;
        RECT 1291.290 821.000 1291.610 821.060 ;
        RECT 1291.095 820.860 1291.610 821.000 ;
        RECT 1291.290 820.800 1291.610 820.860 ;
        RECT 1291.290 786.660 1291.610 786.720 ;
        RECT 1291.095 786.520 1291.610 786.660 ;
        RECT 1291.290 786.460 1291.610 786.520 ;
        RECT 1290.830 738.380 1291.150 738.440 ;
        RECT 1291.750 738.380 1292.070 738.440 ;
        RECT 1290.830 738.240 1292.070 738.380 ;
        RECT 1290.830 738.180 1291.150 738.240 ;
        RECT 1291.750 738.180 1292.070 738.240 ;
        RECT 1291.290 724.440 1291.610 724.500 ;
        RECT 1291.095 724.300 1291.610 724.440 ;
        RECT 1291.290 724.240 1291.610 724.300 ;
        RECT 1291.290 689.760 1291.610 689.820 ;
        RECT 1291.095 689.620 1291.610 689.760 ;
        RECT 1291.290 689.560 1291.610 689.620 ;
        RECT 1290.830 641.820 1291.150 641.880 ;
        RECT 1291.750 641.820 1292.070 641.880 ;
        RECT 1290.830 641.680 1292.070 641.820 ;
        RECT 1290.830 641.620 1291.150 641.680 ;
        RECT 1291.750 641.620 1292.070 641.680 ;
        RECT 1291.290 627.880 1291.610 627.940 ;
        RECT 1291.095 627.740 1291.610 627.880 ;
        RECT 1291.290 627.680 1291.610 627.740 ;
        RECT 1291.290 593.200 1291.610 593.260 ;
        RECT 1291.095 593.060 1291.610 593.200 ;
        RECT 1291.290 593.000 1291.610 593.060 ;
        RECT 1290.830 545.260 1291.150 545.320 ;
        RECT 1291.750 545.260 1292.070 545.320 ;
        RECT 1290.830 545.120 1292.070 545.260 ;
        RECT 1290.830 545.060 1291.150 545.120 ;
        RECT 1291.750 545.060 1292.070 545.120 ;
        RECT 1291.290 531.320 1291.610 531.380 ;
        RECT 1291.095 531.180 1291.610 531.320 ;
        RECT 1291.290 531.120 1291.610 531.180 ;
        RECT 1291.290 496.640 1291.610 496.700 ;
        RECT 1291.095 496.500 1291.610 496.640 ;
        RECT 1291.290 496.440 1291.610 496.500 ;
        RECT 1290.830 448.700 1291.150 448.760 ;
        RECT 1291.750 448.700 1292.070 448.760 ;
        RECT 1290.830 448.560 1292.070 448.700 ;
        RECT 1290.830 448.500 1291.150 448.560 ;
        RECT 1291.750 448.500 1292.070 448.560 ;
        RECT 1291.290 434.760 1291.610 434.820 ;
        RECT 1291.095 434.620 1291.610 434.760 ;
        RECT 1291.290 434.560 1291.610 434.620 ;
        RECT 1291.305 386.480 1291.595 386.525 ;
        RECT 1291.750 386.480 1292.070 386.540 ;
        RECT 1291.305 386.340 1292.070 386.480 ;
        RECT 1291.305 386.295 1291.595 386.340 ;
        RECT 1291.750 386.280 1292.070 386.340 ;
        RECT 1290.830 352.140 1291.150 352.200 ;
        RECT 1290.830 352.000 1291.520 352.140 ;
        RECT 1290.830 351.940 1291.150 352.000 ;
        RECT 1291.380 351.860 1291.520 352.000 ;
        RECT 1291.290 351.600 1291.610 351.860 ;
        RECT 1291.290 241.640 1291.610 241.700 ;
        RECT 1291.750 241.640 1292.070 241.700 ;
        RECT 1291.290 241.500 1292.070 241.640 ;
        RECT 1291.290 241.440 1291.610 241.500 ;
        RECT 1291.750 241.440 1292.070 241.500 ;
        RECT 1291.305 193.020 1291.595 193.065 ;
        RECT 1291.750 193.020 1292.070 193.080 ;
        RECT 1291.305 192.880 1292.070 193.020 ;
        RECT 1291.305 192.835 1291.595 192.880 ;
        RECT 1291.750 192.820 1292.070 192.880 ;
        RECT 1291.290 158.680 1291.610 158.740 ;
        RECT 1291.095 158.540 1291.610 158.680 ;
        RECT 1291.290 158.480 1291.610 158.540 ;
        RECT 1290.830 20.640 1291.150 20.700 ;
        RECT 1293.130 20.640 1293.450 20.700 ;
        RECT 1290.830 20.500 1293.450 20.640 ;
        RECT 1290.830 20.440 1291.150 20.500 ;
        RECT 1293.130 20.440 1293.450 20.500 ;
      LAYER via ;
        RECT 1291.320 1038.400 1291.580 1038.660 ;
        RECT 1291.780 1014.260 1292.040 1014.520 ;
        RECT 1290.860 835.080 1291.120 835.340 ;
        RECT 1291.780 835.080 1292.040 835.340 ;
        RECT 1291.320 820.800 1291.580 821.060 ;
        RECT 1291.320 786.460 1291.580 786.720 ;
        RECT 1290.860 738.180 1291.120 738.440 ;
        RECT 1291.780 738.180 1292.040 738.440 ;
        RECT 1291.320 724.240 1291.580 724.500 ;
        RECT 1291.320 689.560 1291.580 689.820 ;
        RECT 1290.860 641.620 1291.120 641.880 ;
        RECT 1291.780 641.620 1292.040 641.880 ;
        RECT 1291.320 627.680 1291.580 627.940 ;
        RECT 1291.320 593.000 1291.580 593.260 ;
        RECT 1290.860 545.060 1291.120 545.320 ;
        RECT 1291.780 545.060 1292.040 545.320 ;
        RECT 1291.320 531.120 1291.580 531.380 ;
        RECT 1291.320 496.440 1291.580 496.700 ;
        RECT 1290.860 448.500 1291.120 448.760 ;
        RECT 1291.780 448.500 1292.040 448.760 ;
        RECT 1291.320 434.560 1291.580 434.820 ;
        RECT 1291.780 386.280 1292.040 386.540 ;
        RECT 1290.860 351.940 1291.120 352.200 ;
        RECT 1291.320 351.600 1291.580 351.860 ;
        RECT 1291.320 241.440 1291.580 241.700 ;
        RECT 1291.780 241.440 1292.040 241.700 ;
        RECT 1291.780 192.820 1292.040 193.080 ;
        RECT 1291.320 158.480 1291.580 158.740 ;
        RECT 1290.860 20.440 1291.120 20.700 ;
        RECT 1293.160 20.440 1293.420 20.700 ;
      LAYER met2 ;
        RECT 1293.530 1100.650 1293.810 1104.000 ;
        RECT 1293.220 1100.510 1293.810 1100.650 ;
        RECT 1293.220 1088.410 1293.360 1100.510 ;
        RECT 1293.530 1100.000 1293.810 1100.510 ;
        RECT 1291.380 1088.270 1293.360 1088.410 ;
        RECT 1291.380 1038.690 1291.520 1088.270 ;
        RECT 1291.320 1038.370 1291.580 1038.690 ;
        RECT 1291.780 1014.230 1292.040 1014.550 ;
        RECT 1291.840 835.370 1291.980 1014.230 ;
        RECT 1290.860 835.050 1291.120 835.370 ;
        RECT 1291.780 835.050 1292.040 835.370 ;
        RECT 1290.920 834.770 1291.060 835.050 ;
        RECT 1290.920 834.630 1291.520 834.770 ;
        RECT 1291.380 821.090 1291.520 834.630 ;
        RECT 1291.320 820.770 1291.580 821.090 ;
        RECT 1291.320 786.430 1291.580 786.750 ;
        RECT 1291.380 772.890 1291.520 786.430 ;
        RECT 1291.380 772.750 1291.980 772.890 ;
        RECT 1291.840 738.470 1291.980 772.750 ;
        RECT 1290.860 738.210 1291.120 738.470 ;
        RECT 1290.860 738.150 1291.520 738.210 ;
        RECT 1291.780 738.150 1292.040 738.470 ;
        RECT 1290.920 738.070 1291.520 738.150 ;
        RECT 1291.380 724.530 1291.520 738.070 ;
        RECT 1291.320 724.210 1291.580 724.530 ;
        RECT 1291.320 689.530 1291.580 689.850 ;
        RECT 1291.380 676.330 1291.520 689.530 ;
        RECT 1291.380 676.190 1291.980 676.330 ;
        RECT 1291.840 641.910 1291.980 676.190 ;
        RECT 1290.860 641.650 1291.120 641.910 ;
        RECT 1290.860 641.590 1291.520 641.650 ;
        RECT 1291.780 641.590 1292.040 641.910 ;
        RECT 1290.920 641.510 1291.520 641.590 ;
        RECT 1291.380 627.970 1291.520 641.510 ;
        RECT 1291.320 627.650 1291.580 627.970 ;
        RECT 1291.320 592.970 1291.580 593.290 ;
        RECT 1291.380 579.770 1291.520 592.970 ;
        RECT 1291.380 579.630 1291.980 579.770 ;
        RECT 1291.840 545.350 1291.980 579.630 ;
        RECT 1290.860 545.090 1291.120 545.350 ;
        RECT 1290.860 545.030 1291.520 545.090 ;
        RECT 1291.780 545.030 1292.040 545.350 ;
        RECT 1290.920 544.950 1291.520 545.030 ;
        RECT 1291.380 531.410 1291.520 544.950 ;
        RECT 1291.320 531.090 1291.580 531.410 ;
        RECT 1291.320 496.410 1291.580 496.730 ;
        RECT 1291.380 483.210 1291.520 496.410 ;
        RECT 1291.380 483.070 1291.980 483.210 ;
        RECT 1291.840 448.790 1291.980 483.070 ;
        RECT 1290.860 448.530 1291.120 448.790 ;
        RECT 1290.860 448.470 1291.520 448.530 ;
        RECT 1291.780 448.470 1292.040 448.790 ;
        RECT 1290.920 448.390 1291.520 448.470 ;
        RECT 1291.380 434.850 1291.520 448.390 ;
        RECT 1291.320 434.530 1291.580 434.850 ;
        RECT 1291.780 386.250 1292.040 386.570 ;
        RECT 1291.840 386.085 1291.980 386.250 ;
        RECT 1290.850 385.715 1291.130 386.085 ;
        RECT 1291.770 385.715 1292.050 386.085 ;
        RECT 1290.920 352.230 1291.060 385.715 ;
        RECT 1290.860 351.910 1291.120 352.230 ;
        RECT 1291.320 351.570 1291.580 351.890 ;
        RECT 1291.380 303.690 1291.520 351.570 ;
        RECT 1291.380 303.550 1291.980 303.690 ;
        RECT 1291.840 241.730 1291.980 303.550 ;
        RECT 1291.320 241.410 1291.580 241.730 ;
        RECT 1291.780 241.410 1292.040 241.730 ;
        RECT 1291.380 207.130 1291.520 241.410 ;
        RECT 1291.380 206.990 1291.980 207.130 ;
        RECT 1291.840 193.110 1291.980 206.990 ;
        RECT 1291.780 192.790 1292.040 193.110 ;
        RECT 1291.320 158.450 1291.580 158.770 ;
        RECT 1291.380 110.570 1291.520 158.450 ;
        RECT 1291.380 110.430 1291.980 110.570 ;
        RECT 1291.840 62.290 1291.980 110.430 ;
        RECT 1290.920 62.150 1291.980 62.290 ;
        RECT 1290.920 20.730 1291.060 62.150 ;
        RECT 1290.860 20.410 1291.120 20.730 ;
        RECT 1293.160 20.410 1293.420 20.730 ;
        RECT 1293.220 2.000 1293.360 20.410 ;
        RECT 1293.010 -4.000 1293.570 2.000 ;
      LAYER via2 ;
        RECT 1290.850 385.760 1291.130 386.040 ;
        RECT 1291.770 385.760 1292.050 386.040 ;
      LAYER met3 ;
        RECT 1290.825 386.050 1291.155 386.065 ;
        RECT 1291.745 386.050 1292.075 386.065 ;
        RECT 1290.825 385.750 1292.075 386.050 ;
        RECT 1290.825 385.735 1291.155 385.750 ;
        RECT 1291.745 385.735 1292.075 385.750 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1300.030 1087.220 1300.350 1087.280 ;
        RECT 1307.390 1087.220 1307.710 1087.280 ;
        RECT 1300.030 1087.080 1307.710 1087.220 ;
        RECT 1300.030 1087.020 1300.350 1087.080 ;
        RECT 1307.390 1087.020 1307.710 1087.080 ;
        RECT 1307.390 20.640 1307.710 20.700 ;
        RECT 1311.070 20.640 1311.390 20.700 ;
        RECT 1307.390 20.500 1311.390 20.640 ;
        RECT 1307.390 20.440 1307.710 20.500 ;
        RECT 1311.070 20.440 1311.390 20.500 ;
      LAYER via ;
        RECT 1300.060 1087.020 1300.320 1087.280 ;
        RECT 1307.420 1087.020 1307.680 1087.280 ;
        RECT 1307.420 20.440 1307.680 20.700 ;
        RECT 1311.100 20.440 1311.360 20.700 ;
      LAYER met2 ;
        RECT 1299.970 1100.580 1300.250 1104.000 ;
        RECT 1299.970 1100.000 1300.260 1100.580 ;
        RECT 1300.120 1087.310 1300.260 1100.000 ;
        RECT 1300.060 1086.990 1300.320 1087.310 ;
        RECT 1307.420 1086.990 1307.680 1087.310 ;
        RECT 1307.480 20.730 1307.620 1086.990 ;
        RECT 1307.420 20.410 1307.680 20.730 ;
        RECT 1311.100 20.410 1311.360 20.730 ;
        RECT 1311.160 2.000 1311.300 20.410 ;
        RECT 1310.950 -4.000 1311.510 2.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1306.010 1085.520 1306.330 1085.580 ;
        RECT 1306.010 1085.380 1317.740 1085.520 ;
        RECT 1306.010 1085.320 1306.330 1085.380 ;
        RECT 1317.600 1085.180 1317.740 1085.380 ;
        RECT 1326.250 1085.180 1326.570 1085.240 ;
        RECT 1317.600 1085.040 1326.570 1085.180 ;
        RECT 1326.250 1084.980 1326.570 1085.040 ;
        RECT 1326.250 62.120 1326.570 62.180 ;
        RECT 1329.010 62.120 1329.330 62.180 ;
        RECT 1326.250 61.980 1329.330 62.120 ;
        RECT 1326.250 61.920 1326.570 61.980 ;
        RECT 1329.010 61.920 1329.330 61.980 ;
      LAYER via ;
        RECT 1306.040 1085.320 1306.300 1085.580 ;
        RECT 1326.280 1084.980 1326.540 1085.240 ;
        RECT 1326.280 61.920 1326.540 62.180 ;
        RECT 1329.040 61.920 1329.300 62.180 ;
      LAYER met2 ;
        RECT 1305.950 1100.580 1306.230 1104.000 ;
        RECT 1305.950 1100.000 1306.240 1100.580 ;
        RECT 1306.100 1085.610 1306.240 1100.000 ;
        RECT 1306.040 1085.290 1306.300 1085.610 ;
        RECT 1326.280 1084.950 1326.540 1085.270 ;
        RECT 1326.340 62.210 1326.480 1084.950 ;
        RECT 1326.280 61.890 1326.540 62.210 ;
        RECT 1329.040 61.890 1329.300 62.210 ;
        RECT 1329.100 2.000 1329.240 61.890 ;
        RECT 1328.890 -4.000 1329.450 2.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1084.825 1062.585 1084.995 1076.695 ;
      LAYER mcon ;
        RECT 1084.825 1076.525 1084.995 1076.695 ;
      LAYER met1 ;
        RECT 1084.765 1076.680 1085.055 1076.725 ;
        RECT 1085.670 1076.680 1085.990 1076.740 ;
        RECT 1084.765 1076.540 1085.990 1076.680 ;
        RECT 1084.765 1076.495 1085.055 1076.540 ;
        RECT 1085.670 1076.480 1085.990 1076.540 ;
        RECT 1084.750 1062.740 1085.070 1062.800 ;
        RECT 1084.555 1062.600 1085.070 1062.740 ;
        RECT 1084.750 1062.540 1085.070 1062.600 ;
        RECT 1083.370 966.180 1083.690 966.240 ;
        RECT 1084.750 966.180 1085.070 966.240 ;
        RECT 1083.370 966.040 1085.070 966.180 ;
        RECT 1083.370 965.980 1083.690 966.040 ;
        RECT 1084.750 965.980 1085.070 966.040 ;
        RECT 1083.370 869.620 1083.690 869.680 ;
        RECT 1084.750 869.620 1085.070 869.680 ;
        RECT 1083.370 869.480 1085.070 869.620 ;
        RECT 1083.370 869.420 1083.690 869.480 ;
        RECT 1084.750 869.420 1085.070 869.480 ;
        RECT 1084.750 47.980 1085.070 48.240 ;
        RECT 686.390 47.840 686.710 47.900 ;
        RECT 686.390 47.700 1077.620 47.840 ;
        RECT 686.390 47.640 686.710 47.700 ;
        RECT 1077.480 47.500 1077.620 47.700 ;
        RECT 1084.840 47.500 1084.980 47.980 ;
        RECT 1077.480 47.360 1084.980 47.500 ;
      LAYER via ;
        RECT 1085.700 1076.480 1085.960 1076.740 ;
        RECT 1084.780 1062.540 1085.040 1062.800 ;
        RECT 1083.400 965.980 1083.660 966.240 ;
        RECT 1084.780 965.980 1085.040 966.240 ;
        RECT 1083.400 869.420 1083.660 869.680 ;
        RECT 1084.780 869.420 1085.040 869.680 ;
        RECT 1084.780 47.980 1085.040 48.240 ;
        RECT 686.420 47.640 686.680 47.900 ;
      LAYER met2 ;
        RECT 1085.610 1100.580 1085.890 1104.000 ;
        RECT 1085.610 1100.000 1085.900 1100.580 ;
        RECT 1085.760 1076.770 1085.900 1100.000 ;
        RECT 1085.700 1076.450 1085.960 1076.770 ;
        RECT 1084.780 1062.510 1085.040 1062.830 ;
        RECT 1084.840 1014.405 1084.980 1062.510 ;
        RECT 1083.390 1014.035 1083.670 1014.405 ;
        RECT 1084.770 1014.035 1085.050 1014.405 ;
        RECT 1083.460 966.270 1083.600 1014.035 ;
        RECT 1083.400 965.950 1083.660 966.270 ;
        RECT 1084.780 965.950 1085.040 966.270 ;
        RECT 1084.840 917.845 1084.980 965.950 ;
        RECT 1083.390 917.475 1083.670 917.845 ;
        RECT 1084.770 917.475 1085.050 917.845 ;
        RECT 1083.460 869.710 1083.600 917.475 ;
        RECT 1083.400 869.390 1083.660 869.710 ;
        RECT 1084.780 869.390 1085.040 869.710 ;
        RECT 1084.840 48.270 1084.980 869.390 ;
        RECT 1084.780 47.950 1085.040 48.270 ;
        RECT 686.420 47.610 686.680 47.930 ;
        RECT 686.480 2.000 686.620 47.610 ;
        RECT 686.270 -4.000 686.830 2.000 ;
      LAYER via2 ;
        RECT 1083.390 1014.080 1083.670 1014.360 ;
        RECT 1084.770 1014.080 1085.050 1014.360 ;
        RECT 1083.390 917.520 1083.670 917.800 ;
        RECT 1084.770 917.520 1085.050 917.800 ;
      LAYER met3 ;
        RECT 1083.365 1014.370 1083.695 1014.385 ;
        RECT 1084.745 1014.370 1085.075 1014.385 ;
        RECT 1083.365 1014.070 1085.075 1014.370 ;
        RECT 1083.365 1014.055 1083.695 1014.070 ;
        RECT 1084.745 1014.055 1085.075 1014.070 ;
        RECT 1083.365 917.810 1083.695 917.825 ;
        RECT 1084.745 917.810 1085.075 917.825 ;
        RECT 1083.365 917.510 1085.075 917.810 ;
        RECT 1083.365 917.495 1083.695 917.510 ;
        RECT 1084.745 917.495 1085.075 917.510 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1311.990 1085.180 1312.310 1085.240 ;
        RECT 1317.050 1085.180 1317.370 1085.240 ;
        RECT 1311.990 1085.040 1317.370 1085.180 ;
        RECT 1311.990 1084.980 1312.310 1085.040 ;
        RECT 1317.050 1084.980 1317.370 1085.040 ;
        RECT 1317.050 17.920 1317.370 17.980 ;
        RECT 1346.490 17.920 1346.810 17.980 ;
        RECT 1317.050 17.780 1346.810 17.920 ;
        RECT 1317.050 17.720 1317.370 17.780 ;
        RECT 1346.490 17.720 1346.810 17.780 ;
      LAYER via ;
        RECT 1312.020 1084.980 1312.280 1085.240 ;
        RECT 1317.080 1084.980 1317.340 1085.240 ;
        RECT 1317.080 17.720 1317.340 17.980 ;
        RECT 1346.520 17.720 1346.780 17.980 ;
      LAYER met2 ;
        RECT 1311.930 1100.580 1312.210 1104.000 ;
        RECT 1311.930 1100.000 1312.220 1100.580 ;
        RECT 1312.080 1085.270 1312.220 1100.000 ;
        RECT 1312.020 1084.950 1312.280 1085.270 ;
        RECT 1317.080 1084.950 1317.340 1085.270 ;
        RECT 1317.140 18.010 1317.280 1084.950 ;
        RECT 1317.080 17.690 1317.340 18.010 ;
        RECT 1346.520 17.690 1346.780 18.010 ;
        RECT 1346.580 2.000 1346.720 17.690 ;
        RECT 1346.370 -4.000 1346.930 2.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1318.430 1084.500 1318.750 1084.560 ;
        RECT 1348.790 1084.500 1349.110 1084.560 ;
        RECT 1318.430 1084.360 1349.110 1084.500 ;
        RECT 1318.430 1084.300 1318.750 1084.360 ;
        RECT 1348.790 1084.300 1349.110 1084.360 ;
        RECT 1348.790 20.640 1349.110 20.700 ;
        RECT 1364.430 20.640 1364.750 20.700 ;
        RECT 1348.790 20.500 1364.750 20.640 ;
        RECT 1348.790 20.440 1349.110 20.500 ;
        RECT 1364.430 20.440 1364.750 20.500 ;
      LAYER via ;
        RECT 1318.460 1084.300 1318.720 1084.560 ;
        RECT 1348.820 1084.300 1349.080 1084.560 ;
        RECT 1348.820 20.440 1349.080 20.700 ;
        RECT 1364.460 20.440 1364.720 20.700 ;
      LAYER met2 ;
        RECT 1318.370 1100.580 1318.650 1104.000 ;
        RECT 1318.370 1100.000 1318.660 1100.580 ;
        RECT 1318.520 1084.590 1318.660 1100.000 ;
        RECT 1318.460 1084.270 1318.720 1084.590 ;
        RECT 1348.820 1084.270 1349.080 1084.590 ;
        RECT 1348.880 20.730 1349.020 1084.270 ;
        RECT 1348.820 20.410 1349.080 20.730 ;
        RECT 1364.460 20.410 1364.720 20.730 ;
        RECT 1364.520 2.000 1364.660 20.410 ;
        RECT 1364.310 -4.000 1364.870 2.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1365.425 19.125 1365.595 20.315 ;
      LAYER mcon ;
        RECT 1365.425 20.145 1365.595 20.315 ;
      LAYER met1 ;
        RECT 1324.410 1088.580 1324.730 1088.640 ;
        RECT 1328.090 1088.580 1328.410 1088.640 ;
        RECT 1324.410 1088.440 1328.410 1088.580 ;
        RECT 1324.410 1088.380 1324.730 1088.440 ;
        RECT 1328.090 1088.380 1328.410 1088.440 ;
        RECT 1365.365 20.300 1365.655 20.345 ;
        RECT 1382.370 20.300 1382.690 20.360 ;
        RECT 1365.365 20.160 1382.690 20.300 ;
        RECT 1365.365 20.115 1365.655 20.160 ;
        RECT 1382.370 20.100 1382.690 20.160 ;
        RECT 1328.090 19.280 1328.410 19.340 ;
        RECT 1365.365 19.280 1365.655 19.325 ;
        RECT 1328.090 19.140 1365.655 19.280 ;
        RECT 1328.090 19.080 1328.410 19.140 ;
        RECT 1365.365 19.095 1365.655 19.140 ;
      LAYER via ;
        RECT 1324.440 1088.380 1324.700 1088.640 ;
        RECT 1328.120 1088.380 1328.380 1088.640 ;
        RECT 1382.400 20.100 1382.660 20.360 ;
        RECT 1328.120 19.080 1328.380 19.340 ;
      LAYER met2 ;
        RECT 1324.350 1100.580 1324.630 1104.000 ;
        RECT 1324.350 1100.000 1324.640 1100.580 ;
        RECT 1324.500 1088.670 1324.640 1100.000 ;
        RECT 1324.440 1088.350 1324.700 1088.670 ;
        RECT 1328.120 1088.350 1328.380 1088.670 ;
        RECT 1328.180 19.370 1328.320 1088.350 ;
        RECT 1382.400 20.070 1382.660 20.390 ;
        RECT 1328.120 19.050 1328.380 19.370 ;
        RECT 1382.460 2.000 1382.600 20.070 ;
        RECT 1382.250 -4.000 1382.810 2.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1331.310 17.580 1331.630 17.640 ;
        RECT 1331.310 17.440 1359.140 17.580 ;
        RECT 1331.310 17.380 1331.630 17.440 ;
        RECT 1359.000 17.240 1359.140 17.440 ;
        RECT 1359.000 17.100 1383.520 17.240 ;
        RECT 1383.380 16.900 1383.520 17.100 ;
        RECT 1400.310 16.900 1400.630 16.960 ;
        RECT 1383.380 16.760 1400.630 16.900 ;
        RECT 1400.310 16.700 1400.630 16.760 ;
      LAYER via ;
        RECT 1331.340 17.380 1331.600 17.640 ;
        RECT 1400.340 16.700 1400.600 16.960 ;
      LAYER met2 ;
        RECT 1330.330 1100.650 1330.610 1104.000 ;
        RECT 1330.330 1100.510 1331.540 1100.650 ;
        RECT 1330.330 1100.000 1330.610 1100.510 ;
        RECT 1331.400 17.670 1331.540 1100.510 ;
        RECT 1331.340 17.350 1331.600 17.670 ;
        RECT 1400.340 16.670 1400.600 16.990 ;
        RECT 1400.400 2.000 1400.540 16.670 ;
        RECT 1400.190 -4.000 1400.750 2.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1390.725 19.465 1390.895 20.315 ;
      LAYER mcon ;
        RECT 1390.725 20.145 1390.895 20.315 ;
      LAYER met1 ;
        RECT 1364.980 20.500 1383.060 20.640 ;
        RECT 1364.980 20.300 1365.120 20.500 ;
        RECT 1353.020 20.160 1365.120 20.300 ;
        RECT 1382.920 20.300 1383.060 20.500 ;
        RECT 1390.665 20.300 1390.955 20.345 ;
        RECT 1382.920 20.160 1390.955 20.300 ;
        RECT 1337.750 19.960 1338.070 20.020 ;
        RECT 1353.020 19.960 1353.160 20.160 ;
        RECT 1390.665 20.115 1390.955 20.160 ;
        RECT 1337.750 19.820 1353.160 19.960 ;
        RECT 1337.750 19.760 1338.070 19.820 ;
        RECT 1390.665 19.620 1390.955 19.665 ;
        RECT 1418.250 19.620 1418.570 19.680 ;
        RECT 1390.665 19.480 1418.570 19.620 ;
        RECT 1390.665 19.435 1390.955 19.480 ;
        RECT 1418.250 19.420 1418.570 19.480 ;
      LAYER via ;
        RECT 1337.780 19.760 1338.040 20.020 ;
        RECT 1418.280 19.420 1418.540 19.680 ;
      LAYER met2 ;
        RECT 1336.310 1100.650 1336.590 1104.000 ;
        RECT 1336.310 1100.510 1337.980 1100.650 ;
        RECT 1336.310 1100.000 1336.590 1100.510 ;
        RECT 1337.840 20.050 1337.980 1100.510 ;
        RECT 1337.780 19.730 1338.040 20.050 ;
        RECT 1418.280 19.390 1418.540 19.710 ;
        RECT 1418.340 2.000 1418.480 19.390 ;
        RECT 1418.130 -4.000 1418.690 2.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1371.865 16.405 1372.035 19.295 ;
      LAYER mcon ;
        RECT 1371.865 19.125 1372.035 19.295 ;
      LAYER met1 ;
        RECT 1371.805 19.280 1372.095 19.325 ;
        RECT 1435.730 19.280 1436.050 19.340 ;
        RECT 1371.805 19.140 1436.050 19.280 ;
        RECT 1371.805 19.095 1372.095 19.140 ;
        RECT 1435.730 19.080 1436.050 19.140 ;
        RECT 1344.190 16.560 1344.510 16.620 ;
        RECT 1371.805 16.560 1372.095 16.605 ;
        RECT 1344.190 16.420 1372.095 16.560 ;
        RECT 1344.190 16.360 1344.510 16.420 ;
        RECT 1371.805 16.375 1372.095 16.420 ;
      LAYER via ;
        RECT 1435.760 19.080 1436.020 19.340 ;
        RECT 1344.220 16.360 1344.480 16.620 ;
      LAYER met2 ;
        RECT 1342.750 1100.650 1343.030 1104.000 ;
        RECT 1342.750 1100.510 1344.420 1100.650 ;
        RECT 1342.750 1100.000 1343.030 1100.510 ;
        RECT 1344.280 16.650 1344.420 1100.510 ;
        RECT 1435.760 19.050 1436.020 19.370 ;
        RECT 1344.220 16.330 1344.480 16.650 ;
        RECT 1435.820 2.000 1435.960 19.050 ;
        RECT 1435.610 -4.000 1436.170 2.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1350.630 1052.200 1350.950 1052.260 ;
        RECT 1351.550 1052.200 1351.870 1052.260 ;
        RECT 1350.630 1052.060 1351.870 1052.200 ;
        RECT 1350.630 1052.000 1350.950 1052.060 ;
        RECT 1351.550 1052.000 1351.870 1052.060 ;
        RECT 1350.630 949.520 1350.950 949.580 ;
        RECT 1351.550 949.520 1351.870 949.580 ;
        RECT 1350.630 949.380 1351.870 949.520 ;
        RECT 1350.630 949.320 1350.950 949.380 ;
        RECT 1351.550 949.320 1351.870 949.380 ;
        RECT 1350.630 907.360 1350.950 907.420 ;
        RECT 1351.550 907.360 1351.870 907.420 ;
        RECT 1350.630 907.220 1351.870 907.360 ;
        RECT 1350.630 907.160 1350.950 907.220 ;
        RECT 1351.550 907.160 1351.870 907.220 ;
        RECT 1350.630 852.960 1350.950 853.020 ;
        RECT 1351.550 852.960 1351.870 853.020 ;
        RECT 1350.630 852.820 1351.870 852.960 ;
        RECT 1350.630 852.760 1350.950 852.820 ;
        RECT 1351.550 852.760 1351.870 852.820 ;
        RECT 1350.630 810.800 1350.950 810.860 ;
        RECT 1351.550 810.800 1351.870 810.860 ;
        RECT 1350.630 810.660 1351.870 810.800 ;
        RECT 1350.630 810.600 1350.950 810.660 ;
        RECT 1351.550 810.600 1351.870 810.660 ;
        RECT 1350.630 762.520 1350.950 762.580 ;
        RECT 1351.550 762.520 1351.870 762.580 ;
        RECT 1350.630 762.380 1351.870 762.520 ;
        RECT 1350.630 762.320 1350.950 762.380 ;
        RECT 1351.550 762.320 1351.870 762.380 ;
        RECT 1350.630 714.240 1350.950 714.300 ;
        RECT 1351.550 714.240 1351.870 714.300 ;
        RECT 1350.630 714.100 1351.870 714.240 ;
        RECT 1350.630 714.040 1350.950 714.100 ;
        RECT 1351.550 714.040 1351.870 714.100 ;
        RECT 1350.630 659.840 1350.950 659.900 ;
        RECT 1351.550 659.840 1351.870 659.900 ;
        RECT 1350.630 659.700 1351.870 659.840 ;
        RECT 1350.630 659.640 1350.950 659.700 ;
        RECT 1351.550 659.640 1351.870 659.700 ;
        RECT 1350.630 617.680 1350.950 617.740 ;
        RECT 1351.550 617.680 1351.870 617.740 ;
        RECT 1350.630 617.540 1351.870 617.680 ;
        RECT 1350.630 617.480 1350.950 617.540 ;
        RECT 1351.550 617.480 1351.870 617.540 ;
        RECT 1350.630 569.400 1350.950 569.460 ;
        RECT 1351.550 569.400 1351.870 569.460 ;
        RECT 1350.630 569.260 1351.870 569.400 ;
        RECT 1350.630 569.200 1350.950 569.260 ;
        RECT 1351.550 569.200 1351.870 569.260 ;
        RECT 1350.630 527.240 1350.950 527.300 ;
        RECT 1351.550 527.240 1351.870 527.300 ;
        RECT 1350.630 527.100 1351.870 527.240 ;
        RECT 1350.630 527.040 1350.950 527.100 ;
        RECT 1351.550 527.040 1351.870 527.100 ;
        RECT 1350.630 472.840 1350.950 472.900 ;
        RECT 1351.550 472.840 1351.870 472.900 ;
        RECT 1350.630 472.700 1351.870 472.840 ;
        RECT 1350.630 472.640 1350.950 472.700 ;
        RECT 1351.550 472.640 1351.870 472.700 ;
        RECT 1350.630 430.680 1350.950 430.740 ;
        RECT 1351.550 430.680 1351.870 430.740 ;
        RECT 1350.630 430.540 1351.870 430.680 ;
        RECT 1350.630 430.480 1350.950 430.540 ;
        RECT 1351.550 430.480 1351.870 430.540 ;
        RECT 1350.630 376.280 1350.950 376.340 ;
        RECT 1351.550 376.280 1351.870 376.340 ;
        RECT 1350.630 376.140 1351.870 376.280 ;
        RECT 1350.630 376.080 1350.950 376.140 ;
        RECT 1351.550 376.080 1351.870 376.140 ;
        RECT 1350.630 327.660 1350.950 327.720 ;
        RECT 1351.550 327.660 1351.870 327.720 ;
        RECT 1350.630 327.520 1351.870 327.660 ;
        RECT 1350.630 327.460 1350.950 327.520 ;
        RECT 1351.550 327.460 1351.870 327.520 ;
        RECT 1350.630 273.260 1350.950 273.320 ;
        RECT 1351.550 273.260 1351.870 273.320 ;
        RECT 1350.630 273.120 1351.870 273.260 ;
        RECT 1350.630 273.060 1350.950 273.120 ;
        RECT 1351.550 273.060 1351.870 273.120 ;
        RECT 1350.630 237.220 1350.950 237.280 ;
        RECT 1351.550 237.220 1351.870 237.280 ;
        RECT 1350.630 237.080 1351.870 237.220 ;
        RECT 1350.630 237.020 1350.950 237.080 ;
        RECT 1351.550 237.020 1351.870 237.080 ;
        RECT 1350.630 176.700 1350.950 176.760 ;
        RECT 1351.550 176.700 1351.870 176.760 ;
        RECT 1350.630 176.560 1351.870 176.700 ;
        RECT 1350.630 176.500 1350.950 176.560 ;
        RECT 1351.550 176.500 1351.870 176.560 ;
        RECT 1350.630 134.540 1350.950 134.600 ;
        RECT 1351.550 134.540 1351.870 134.600 ;
        RECT 1350.630 134.400 1351.870 134.540 ;
        RECT 1350.630 134.340 1350.950 134.400 ;
        RECT 1351.550 134.340 1351.870 134.400 ;
        RECT 1350.630 86.260 1350.950 86.320 ;
        RECT 1351.550 86.260 1351.870 86.320 ;
        RECT 1350.630 86.120 1351.870 86.260 ;
        RECT 1350.630 86.060 1350.950 86.120 ;
        RECT 1351.550 86.060 1351.870 86.120 ;
        RECT 1350.630 17.920 1350.950 17.980 ;
        RECT 1453.670 17.920 1453.990 17.980 ;
        RECT 1350.630 17.780 1453.990 17.920 ;
        RECT 1350.630 17.720 1350.950 17.780 ;
        RECT 1453.670 17.720 1453.990 17.780 ;
      LAYER via ;
        RECT 1350.660 1052.000 1350.920 1052.260 ;
        RECT 1351.580 1052.000 1351.840 1052.260 ;
        RECT 1350.660 949.320 1350.920 949.580 ;
        RECT 1351.580 949.320 1351.840 949.580 ;
        RECT 1350.660 907.160 1350.920 907.420 ;
        RECT 1351.580 907.160 1351.840 907.420 ;
        RECT 1350.660 852.760 1350.920 853.020 ;
        RECT 1351.580 852.760 1351.840 853.020 ;
        RECT 1350.660 810.600 1350.920 810.860 ;
        RECT 1351.580 810.600 1351.840 810.860 ;
        RECT 1350.660 762.320 1350.920 762.580 ;
        RECT 1351.580 762.320 1351.840 762.580 ;
        RECT 1350.660 714.040 1350.920 714.300 ;
        RECT 1351.580 714.040 1351.840 714.300 ;
        RECT 1350.660 659.640 1350.920 659.900 ;
        RECT 1351.580 659.640 1351.840 659.900 ;
        RECT 1350.660 617.480 1350.920 617.740 ;
        RECT 1351.580 617.480 1351.840 617.740 ;
        RECT 1350.660 569.200 1350.920 569.460 ;
        RECT 1351.580 569.200 1351.840 569.460 ;
        RECT 1350.660 527.040 1350.920 527.300 ;
        RECT 1351.580 527.040 1351.840 527.300 ;
        RECT 1350.660 472.640 1350.920 472.900 ;
        RECT 1351.580 472.640 1351.840 472.900 ;
        RECT 1350.660 430.480 1350.920 430.740 ;
        RECT 1351.580 430.480 1351.840 430.740 ;
        RECT 1350.660 376.080 1350.920 376.340 ;
        RECT 1351.580 376.080 1351.840 376.340 ;
        RECT 1350.660 327.460 1350.920 327.720 ;
        RECT 1351.580 327.460 1351.840 327.720 ;
        RECT 1350.660 273.060 1350.920 273.320 ;
        RECT 1351.580 273.060 1351.840 273.320 ;
        RECT 1350.660 237.020 1350.920 237.280 ;
        RECT 1351.580 237.020 1351.840 237.280 ;
        RECT 1350.660 176.500 1350.920 176.760 ;
        RECT 1351.580 176.500 1351.840 176.760 ;
        RECT 1350.660 134.340 1350.920 134.600 ;
        RECT 1351.580 134.340 1351.840 134.600 ;
        RECT 1350.660 86.060 1350.920 86.320 ;
        RECT 1351.580 86.060 1351.840 86.320 ;
        RECT 1350.660 17.720 1350.920 17.980 ;
        RECT 1453.700 17.720 1453.960 17.980 ;
      LAYER met2 ;
        RECT 1348.730 1100.650 1349.010 1104.000 ;
        RECT 1348.730 1100.510 1350.860 1100.650 ;
        RECT 1348.730 1100.000 1349.010 1100.510 ;
        RECT 1350.720 1052.290 1350.860 1100.510 ;
        RECT 1350.660 1051.970 1350.920 1052.290 ;
        RECT 1351.580 1051.970 1351.840 1052.290 ;
        RECT 1351.640 949.610 1351.780 1051.970 ;
        RECT 1350.660 949.290 1350.920 949.610 ;
        RECT 1351.580 949.290 1351.840 949.610 ;
        RECT 1350.720 907.450 1350.860 949.290 ;
        RECT 1350.660 907.130 1350.920 907.450 ;
        RECT 1351.580 907.130 1351.840 907.450 ;
        RECT 1351.640 853.050 1351.780 907.130 ;
        RECT 1350.660 852.730 1350.920 853.050 ;
        RECT 1351.580 852.730 1351.840 853.050 ;
        RECT 1350.720 810.890 1350.860 852.730 ;
        RECT 1350.660 810.570 1350.920 810.890 ;
        RECT 1351.580 810.570 1351.840 810.890 ;
        RECT 1351.640 762.610 1351.780 810.570 ;
        RECT 1350.660 762.290 1350.920 762.610 ;
        RECT 1351.580 762.290 1351.840 762.610 ;
        RECT 1350.720 714.330 1350.860 762.290 ;
        RECT 1350.660 714.010 1350.920 714.330 ;
        RECT 1351.580 714.010 1351.840 714.330 ;
        RECT 1351.640 659.930 1351.780 714.010 ;
        RECT 1350.660 659.610 1350.920 659.930 ;
        RECT 1351.580 659.610 1351.840 659.930 ;
        RECT 1350.720 617.770 1350.860 659.610 ;
        RECT 1350.660 617.450 1350.920 617.770 ;
        RECT 1351.580 617.450 1351.840 617.770 ;
        RECT 1351.640 569.490 1351.780 617.450 ;
        RECT 1350.660 569.170 1350.920 569.490 ;
        RECT 1351.580 569.170 1351.840 569.490 ;
        RECT 1350.720 527.330 1350.860 569.170 ;
        RECT 1350.660 527.010 1350.920 527.330 ;
        RECT 1351.580 527.010 1351.840 527.330 ;
        RECT 1351.640 472.930 1351.780 527.010 ;
        RECT 1350.660 472.610 1350.920 472.930 ;
        RECT 1351.580 472.610 1351.840 472.930 ;
        RECT 1350.720 430.770 1350.860 472.610 ;
        RECT 1350.660 430.450 1350.920 430.770 ;
        RECT 1351.580 430.450 1351.840 430.770 ;
        RECT 1351.640 376.370 1351.780 430.450 ;
        RECT 1350.660 376.050 1350.920 376.370 ;
        RECT 1351.580 376.050 1351.840 376.370 ;
        RECT 1350.720 327.750 1350.860 376.050 ;
        RECT 1350.660 327.430 1350.920 327.750 ;
        RECT 1351.580 327.430 1351.840 327.750 ;
        RECT 1351.640 273.350 1351.780 327.430 ;
        RECT 1350.660 273.030 1350.920 273.350 ;
        RECT 1351.580 273.030 1351.840 273.350 ;
        RECT 1350.720 237.310 1350.860 273.030 ;
        RECT 1350.660 236.990 1350.920 237.310 ;
        RECT 1351.580 236.990 1351.840 237.310 ;
        RECT 1351.640 176.790 1351.780 236.990 ;
        RECT 1350.660 176.470 1350.920 176.790 ;
        RECT 1351.580 176.470 1351.840 176.790 ;
        RECT 1350.720 134.630 1350.860 176.470 ;
        RECT 1350.660 134.310 1350.920 134.630 ;
        RECT 1351.580 134.310 1351.840 134.630 ;
        RECT 1351.640 86.350 1351.780 134.310 ;
        RECT 1350.660 86.030 1350.920 86.350 ;
        RECT 1351.580 86.030 1351.840 86.350 ;
        RECT 1350.720 18.010 1350.860 86.030 ;
        RECT 1350.660 17.690 1350.920 18.010 ;
        RECT 1453.700 17.690 1453.960 18.010 ;
        RECT 1453.760 2.000 1453.900 17.690 ;
        RECT 1453.550 -4.000 1454.110 2.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1354.770 1084.840 1355.090 1084.900 ;
        RECT 1417.790 1084.840 1418.110 1084.900 ;
        RECT 1354.770 1084.700 1418.110 1084.840 ;
        RECT 1354.770 1084.640 1355.090 1084.700 ;
        RECT 1417.790 1084.640 1418.110 1084.700 ;
        RECT 1471.610 14.180 1471.930 14.240 ;
        RECT 1424.320 14.040 1471.930 14.180 ;
        RECT 1417.790 13.840 1418.110 13.900 ;
        RECT 1424.320 13.840 1424.460 14.040 ;
        RECT 1471.610 13.980 1471.930 14.040 ;
        RECT 1417.790 13.700 1424.460 13.840 ;
        RECT 1417.790 13.640 1418.110 13.700 ;
      LAYER via ;
        RECT 1354.800 1084.640 1355.060 1084.900 ;
        RECT 1417.820 1084.640 1418.080 1084.900 ;
        RECT 1417.820 13.640 1418.080 13.900 ;
        RECT 1471.640 13.980 1471.900 14.240 ;
      LAYER met2 ;
        RECT 1354.710 1100.580 1354.990 1104.000 ;
        RECT 1354.710 1100.000 1355.000 1100.580 ;
        RECT 1354.860 1084.930 1355.000 1100.000 ;
        RECT 1354.800 1084.610 1355.060 1084.930 ;
        RECT 1417.820 1084.610 1418.080 1084.930 ;
        RECT 1417.880 13.930 1418.020 1084.610 ;
        RECT 1471.640 13.950 1471.900 14.270 ;
        RECT 1417.820 13.610 1418.080 13.930 ;
        RECT 1471.700 2.000 1471.840 13.950 ;
        RECT 1471.490 -4.000 1472.050 2.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1361.210 1085.180 1361.530 1085.240 ;
        RECT 1361.210 1085.040 1432.740 1085.180 ;
        RECT 1361.210 1084.980 1361.530 1085.040 ;
        RECT 1432.600 1084.840 1432.740 1085.040 ;
        RECT 1452.290 1084.840 1452.610 1084.900 ;
        RECT 1432.600 1084.700 1452.610 1084.840 ;
        RECT 1452.290 1084.640 1452.610 1084.700 ;
        RECT 1452.290 14.520 1452.610 14.580 ;
        RECT 1489.550 14.520 1489.870 14.580 ;
        RECT 1452.290 14.380 1489.870 14.520 ;
        RECT 1452.290 14.320 1452.610 14.380 ;
        RECT 1489.550 14.320 1489.870 14.380 ;
      LAYER via ;
        RECT 1361.240 1084.980 1361.500 1085.240 ;
        RECT 1452.320 1084.640 1452.580 1084.900 ;
        RECT 1452.320 14.320 1452.580 14.580 ;
        RECT 1489.580 14.320 1489.840 14.580 ;
      LAYER met2 ;
        RECT 1361.150 1100.580 1361.430 1104.000 ;
        RECT 1361.150 1100.000 1361.440 1100.580 ;
        RECT 1361.300 1085.270 1361.440 1100.000 ;
        RECT 1361.240 1084.950 1361.500 1085.270 ;
        RECT 1452.320 1084.610 1452.580 1084.930 ;
        RECT 1452.380 14.610 1452.520 1084.610 ;
        RECT 1452.320 14.290 1452.580 14.610 ;
        RECT 1489.580 14.290 1489.840 14.610 ;
        RECT 1489.640 2.000 1489.780 14.290 ;
        RECT 1489.430 -4.000 1489.990 2.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1410.045 1084.345 1410.215 1085.535 ;
      LAYER mcon ;
        RECT 1410.045 1085.365 1410.215 1085.535 ;
      LAYER met1 ;
        RECT 1409.985 1085.520 1410.275 1085.565 ;
        RECT 1409.985 1085.380 1464.940 1085.520 ;
        RECT 1409.985 1085.335 1410.275 1085.380 ;
        RECT 1464.800 1084.840 1464.940 1085.380 ;
        RECT 1486.790 1084.840 1487.110 1084.900 ;
        RECT 1464.800 1084.700 1487.110 1084.840 ;
        RECT 1486.790 1084.640 1487.110 1084.700 ;
        RECT 1367.190 1084.500 1367.510 1084.560 ;
        RECT 1409.985 1084.500 1410.275 1084.545 ;
        RECT 1367.190 1084.360 1410.275 1084.500 ;
        RECT 1367.190 1084.300 1367.510 1084.360 ;
        RECT 1409.985 1084.315 1410.275 1084.360 ;
        RECT 1486.790 17.240 1487.110 17.300 ;
        RECT 1507.030 17.240 1507.350 17.300 ;
        RECT 1486.790 17.100 1507.350 17.240 ;
        RECT 1486.790 17.040 1487.110 17.100 ;
        RECT 1507.030 17.040 1507.350 17.100 ;
      LAYER via ;
        RECT 1486.820 1084.640 1487.080 1084.900 ;
        RECT 1367.220 1084.300 1367.480 1084.560 ;
        RECT 1486.820 17.040 1487.080 17.300 ;
        RECT 1507.060 17.040 1507.320 17.300 ;
      LAYER met2 ;
        RECT 1367.130 1100.580 1367.410 1104.000 ;
        RECT 1367.130 1100.000 1367.420 1100.580 ;
        RECT 1367.280 1084.590 1367.420 1100.000 ;
        RECT 1486.820 1084.610 1487.080 1084.930 ;
        RECT 1367.220 1084.270 1367.480 1084.590 ;
        RECT 1486.880 17.330 1487.020 1084.610 ;
        RECT 1486.820 17.010 1487.080 17.330 ;
        RECT 1507.060 17.010 1507.320 17.330 ;
        RECT 1507.120 2.000 1507.260 17.010 ;
        RECT 1506.910 -4.000 1507.470 2.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 704.330 44.440 704.650 44.500 ;
        RECT 1090.730 44.440 1091.050 44.500 ;
        RECT 704.330 44.300 1091.050 44.440 ;
        RECT 704.330 44.240 704.650 44.300 ;
        RECT 1090.730 44.240 1091.050 44.300 ;
      LAYER via ;
        RECT 704.360 44.240 704.620 44.500 ;
        RECT 1090.760 44.240 1091.020 44.500 ;
      LAYER met2 ;
        RECT 1091.590 1100.650 1091.870 1104.000 ;
        RECT 1090.820 1100.510 1091.870 1100.650 ;
        RECT 1090.820 44.530 1090.960 1100.510 ;
        RECT 1091.590 1100.000 1091.870 1100.510 ;
        RECT 704.360 44.210 704.620 44.530 ;
        RECT 1090.760 44.210 1091.020 44.530 ;
        RECT 704.420 2.000 704.560 44.210 ;
        RECT 704.210 -4.000 704.770 2.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1500.590 1085.860 1500.910 1085.920 ;
        RECT 1409.600 1085.720 1481.960 1085.860 ;
        RECT 1373.170 1085.520 1373.490 1085.580 ;
        RECT 1409.600 1085.520 1409.740 1085.720 ;
        RECT 1373.170 1085.380 1409.740 1085.520 ;
        RECT 1481.820 1085.520 1481.960 1085.720 ;
        RECT 1489.640 1085.720 1500.910 1085.860 ;
        RECT 1489.640 1085.520 1489.780 1085.720 ;
        RECT 1500.590 1085.660 1500.910 1085.720 ;
        RECT 1481.820 1085.380 1489.780 1085.520 ;
        RECT 1373.170 1085.320 1373.490 1085.380 ;
        RECT 1500.590 15.540 1500.910 15.600 ;
        RECT 1524.970 15.540 1525.290 15.600 ;
        RECT 1500.590 15.400 1525.290 15.540 ;
        RECT 1500.590 15.340 1500.910 15.400 ;
        RECT 1524.970 15.340 1525.290 15.400 ;
      LAYER via ;
        RECT 1373.200 1085.320 1373.460 1085.580 ;
        RECT 1500.620 1085.660 1500.880 1085.920 ;
        RECT 1500.620 15.340 1500.880 15.600 ;
        RECT 1525.000 15.340 1525.260 15.600 ;
      LAYER met2 ;
        RECT 1373.110 1100.580 1373.390 1104.000 ;
        RECT 1373.110 1100.000 1373.400 1100.580 ;
        RECT 1373.260 1085.610 1373.400 1100.000 ;
        RECT 1500.620 1085.630 1500.880 1085.950 ;
        RECT 1373.200 1085.290 1373.460 1085.610 ;
        RECT 1500.680 15.630 1500.820 1085.630 ;
        RECT 1500.620 15.310 1500.880 15.630 ;
        RECT 1525.000 15.310 1525.260 15.630 ;
        RECT 1525.060 2.000 1525.200 15.310 ;
        RECT 1524.850 -4.000 1525.410 2.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1407.745 1088.425 1407.915 1089.275 ;
        RECT 1462.945 1088.425 1463.575 1088.595 ;
        RECT 1463.405 1087.065 1463.575 1088.425 ;
      LAYER mcon ;
        RECT 1407.745 1089.105 1407.915 1089.275 ;
      LAYER met1 ;
        RECT 1407.685 1089.260 1407.975 1089.305 ;
        RECT 1379.700 1089.120 1407.975 1089.260 ;
        RECT 1379.700 1088.980 1379.840 1089.120 ;
        RECT 1407.685 1089.075 1407.975 1089.120 ;
        RECT 1379.610 1088.720 1379.930 1088.980 ;
        RECT 1407.685 1088.580 1407.975 1088.625 ;
        RECT 1462.885 1088.580 1463.175 1088.625 ;
        RECT 1407.685 1088.440 1463.175 1088.580 ;
        RECT 1407.685 1088.395 1407.975 1088.440 ;
        RECT 1462.885 1088.395 1463.175 1088.440 ;
        RECT 1463.345 1087.220 1463.635 1087.265 ;
        RECT 1507.490 1087.220 1507.810 1087.280 ;
        RECT 1463.345 1087.080 1507.810 1087.220 ;
        RECT 1463.345 1087.035 1463.635 1087.080 ;
        RECT 1507.490 1087.020 1507.810 1087.080 ;
        RECT 1507.490 15.880 1507.810 15.940 ;
        RECT 1507.490 15.740 1525.660 15.880 ;
        RECT 1507.490 15.680 1507.810 15.740 ;
        RECT 1525.520 15.200 1525.660 15.740 ;
        RECT 1542.910 15.200 1543.230 15.260 ;
        RECT 1525.520 15.060 1543.230 15.200 ;
        RECT 1542.910 15.000 1543.230 15.060 ;
      LAYER via ;
        RECT 1379.640 1088.720 1379.900 1088.980 ;
        RECT 1507.520 1087.020 1507.780 1087.280 ;
        RECT 1507.520 15.680 1507.780 15.940 ;
        RECT 1542.940 15.000 1543.200 15.260 ;
      LAYER met2 ;
        RECT 1379.550 1100.580 1379.830 1104.000 ;
        RECT 1379.550 1100.000 1379.840 1100.580 ;
        RECT 1379.700 1089.885 1379.840 1100.000 ;
        RECT 1379.630 1089.515 1379.910 1089.885 ;
        RECT 1379.640 1088.690 1379.900 1089.010 ;
        RECT 1379.700 1088.525 1379.840 1088.690 ;
        RECT 1379.630 1088.155 1379.910 1088.525 ;
        RECT 1507.520 1086.990 1507.780 1087.310 ;
        RECT 1507.580 15.970 1507.720 1086.990 ;
        RECT 1507.520 15.650 1507.780 15.970 ;
        RECT 1542.940 14.970 1543.200 15.290 ;
        RECT 1543.000 2.000 1543.140 14.970 ;
        RECT 1542.790 -4.000 1543.350 2.000 ;
      LAYER via2 ;
        RECT 1379.630 1089.560 1379.910 1089.840 ;
        RECT 1379.630 1088.200 1379.910 1088.480 ;
      LAYER met3 ;
        RECT 1379.605 1089.860 1379.935 1089.865 ;
        RECT 1379.350 1089.850 1379.935 1089.860 ;
        RECT 1379.150 1089.550 1379.935 1089.850 ;
        RECT 1379.350 1089.540 1379.935 1089.550 ;
        RECT 1379.605 1089.535 1379.935 1089.540 ;
        RECT 1379.605 1088.500 1379.935 1088.505 ;
        RECT 1379.350 1088.490 1379.935 1088.500 ;
        RECT 1379.150 1088.190 1379.935 1088.490 ;
        RECT 1379.350 1088.180 1379.935 1088.190 ;
        RECT 1379.605 1088.175 1379.935 1088.180 ;
      LAYER via3 ;
        RECT 1379.380 1089.540 1379.700 1089.860 ;
        RECT 1379.380 1088.180 1379.700 1088.500 ;
      LAYER met4 ;
        RECT 1379.375 1089.535 1379.705 1089.865 ;
        RECT 1379.390 1088.505 1379.690 1089.535 ;
        RECT 1379.375 1088.175 1379.705 1088.505 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1514.390 1088.240 1514.710 1088.300 ;
        RECT 1503.440 1088.100 1514.710 1088.240 ;
        RECT 1385.590 1087.900 1385.910 1087.960 ;
        RECT 1503.440 1087.900 1503.580 1088.100 ;
        RECT 1514.390 1088.040 1514.710 1088.100 ;
        RECT 1385.590 1087.760 1503.580 1087.900 ;
        RECT 1385.590 1087.700 1385.910 1087.760 ;
        RECT 1514.390 14.180 1514.710 14.240 ;
        RECT 1560.850 14.180 1561.170 14.240 ;
        RECT 1514.390 14.040 1561.170 14.180 ;
        RECT 1514.390 13.980 1514.710 14.040 ;
        RECT 1560.850 13.980 1561.170 14.040 ;
      LAYER via ;
        RECT 1385.620 1087.700 1385.880 1087.960 ;
        RECT 1514.420 1088.040 1514.680 1088.300 ;
        RECT 1514.420 13.980 1514.680 14.240 ;
        RECT 1560.880 13.980 1561.140 14.240 ;
      LAYER met2 ;
        RECT 1385.530 1100.580 1385.810 1104.000 ;
        RECT 1385.530 1100.000 1385.820 1100.580 ;
        RECT 1385.680 1087.990 1385.820 1100.000 ;
        RECT 1514.420 1088.010 1514.680 1088.330 ;
        RECT 1385.620 1087.670 1385.880 1087.990 ;
        RECT 1514.480 14.270 1514.620 1088.010 ;
        RECT 1514.420 13.950 1514.680 14.270 ;
        RECT 1560.880 13.950 1561.140 14.270 ;
        RECT 1560.940 2.000 1561.080 13.950 ;
        RECT 1560.730 -4.000 1561.290 2.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1391.570 1088.920 1391.890 1088.980 ;
        RECT 1521.290 1088.920 1521.610 1088.980 ;
        RECT 1391.570 1088.780 1521.610 1088.920 ;
        RECT 1391.570 1088.720 1391.890 1088.780 ;
        RECT 1521.290 1088.720 1521.610 1088.780 ;
        RECT 1521.290 14.520 1521.610 14.580 ;
        RECT 1578.790 14.520 1579.110 14.580 ;
        RECT 1521.290 14.380 1579.110 14.520 ;
        RECT 1521.290 14.320 1521.610 14.380 ;
        RECT 1578.790 14.320 1579.110 14.380 ;
      LAYER via ;
        RECT 1391.600 1088.720 1391.860 1088.980 ;
        RECT 1521.320 1088.720 1521.580 1088.980 ;
        RECT 1521.320 14.320 1521.580 14.580 ;
        RECT 1578.820 14.320 1579.080 14.580 ;
      LAYER met2 ;
        RECT 1391.510 1100.580 1391.790 1104.000 ;
        RECT 1391.510 1100.000 1391.800 1100.580 ;
        RECT 1391.660 1089.010 1391.800 1100.000 ;
        RECT 1391.600 1088.690 1391.860 1089.010 ;
        RECT 1521.320 1088.690 1521.580 1089.010 ;
        RECT 1521.380 14.610 1521.520 1088.690 ;
        RECT 1521.320 14.290 1521.580 14.610 ;
        RECT 1578.820 14.290 1579.080 14.610 ;
        RECT 1578.880 2.000 1579.020 14.290 ;
        RECT 1578.670 -4.000 1579.230 2.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1476.745 1085.025 1476.915 1088.255 ;
        RECT 1541.605 14.705 1541.775 15.555 ;
      LAYER mcon ;
        RECT 1476.745 1088.085 1476.915 1088.255 ;
        RECT 1541.605 15.385 1541.775 15.555 ;
      LAYER met1 ;
        RECT 1398.010 1088.240 1398.330 1088.300 ;
        RECT 1476.685 1088.240 1476.975 1088.285 ;
        RECT 1398.010 1088.100 1476.975 1088.240 ;
        RECT 1398.010 1088.040 1398.330 1088.100 ;
        RECT 1476.685 1088.055 1476.975 1088.100 ;
        RECT 1476.685 1085.180 1476.975 1085.225 ;
        RECT 1476.685 1085.040 1487.480 1085.180 ;
        RECT 1476.685 1084.995 1476.975 1085.040 ;
        RECT 1487.340 1084.840 1487.480 1085.040 ;
        RECT 1528.190 1084.840 1528.510 1084.900 ;
        RECT 1487.340 1084.700 1528.510 1084.840 ;
        RECT 1528.190 1084.640 1528.510 1084.700 ;
        RECT 1528.190 15.540 1528.510 15.600 ;
        RECT 1541.545 15.540 1541.835 15.585 ;
        RECT 1528.190 15.400 1541.835 15.540 ;
        RECT 1528.190 15.340 1528.510 15.400 ;
        RECT 1541.545 15.355 1541.835 15.400 ;
        RECT 1541.545 14.860 1541.835 14.905 ;
        RECT 1596.270 14.860 1596.590 14.920 ;
        RECT 1541.545 14.720 1596.590 14.860 ;
        RECT 1541.545 14.675 1541.835 14.720 ;
        RECT 1596.270 14.660 1596.590 14.720 ;
      LAYER via ;
        RECT 1398.040 1088.040 1398.300 1088.300 ;
        RECT 1528.220 1084.640 1528.480 1084.900 ;
        RECT 1528.220 15.340 1528.480 15.600 ;
        RECT 1596.300 14.660 1596.560 14.920 ;
      LAYER met2 ;
        RECT 1397.950 1100.580 1398.230 1104.000 ;
        RECT 1397.950 1100.000 1398.240 1100.580 ;
        RECT 1398.100 1088.330 1398.240 1100.000 ;
        RECT 1398.040 1088.010 1398.300 1088.330 ;
        RECT 1528.220 1084.610 1528.480 1084.930 ;
        RECT 1528.280 15.630 1528.420 1084.610 ;
        RECT 1528.220 15.310 1528.480 15.630 ;
        RECT 1596.300 14.630 1596.560 14.950 ;
        RECT 1596.360 2.000 1596.500 14.630 ;
        RECT 1596.150 -4.000 1596.710 2.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1531.485 14.705 1531.655 16.235 ;
      LAYER mcon ;
        RECT 1531.485 16.065 1531.655 16.235 ;
      LAYER met1 ;
        RECT 1403.990 1086.540 1404.310 1086.600 ;
        RECT 1403.990 1086.400 1438.720 1086.540 ;
        RECT 1403.990 1086.340 1404.310 1086.400 ;
        RECT 1438.580 1086.200 1438.720 1086.400 ;
        RECT 1528.650 1086.200 1528.970 1086.260 ;
        RECT 1438.580 1086.060 1528.970 1086.200 ;
        RECT 1528.650 1086.000 1528.970 1086.060 ;
        RECT 1531.425 16.220 1531.715 16.265 ;
        RECT 1614.210 16.220 1614.530 16.280 ;
        RECT 1531.425 16.080 1614.530 16.220 ;
        RECT 1531.425 16.035 1531.715 16.080 ;
        RECT 1614.210 16.020 1614.530 16.080 ;
        RECT 1528.650 14.860 1528.970 14.920 ;
        RECT 1531.425 14.860 1531.715 14.905 ;
        RECT 1528.650 14.720 1531.715 14.860 ;
        RECT 1528.650 14.660 1528.970 14.720 ;
        RECT 1531.425 14.675 1531.715 14.720 ;
      LAYER via ;
        RECT 1404.020 1086.340 1404.280 1086.600 ;
        RECT 1528.680 1086.000 1528.940 1086.260 ;
        RECT 1614.240 16.020 1614.500 16.280 ;
        RECT 1528.680 14.660 1528.940 14.920 ;
      LAYER met2 ;
        RECT 1403.930 1100.580 1404.210 1104.000 ;
        RECT 1403.930 1100.000 1404.220 1100.580 ;
        RECT 1404.080 1086.630 1404.220 1100.000 ;
        RECT 1404.020 1086.310 1404.280 1086.630 ;
        RECT 1528.680 1085.970 1528.940 1086.290 ;
        RECT 1528.740 14.950 1528.880 1085.970 ;
        RECT 1614.240 15.990 1614.500 16.310 ;
        RECT 1528.680 14.630 1528.940 14.950 ;
        RECT 1614.300 2.000 1614.440 15.990 ;
        RECT 1614.090 -4.000 1614.650 2.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1567.825 15.385 1567.995 16.575 ;
      LAYER mcon ;
        RECT 1567.825 16.405 1567.995 16.575 ;
      LAYER met1 ;
        RECT 1409.970 1089.940 1410.290 1090.000 ;
        RECT 1541.990 1089.940 1542.310 1090.000 ;
        RECT 1409.970 1089.800 1542.310 1089.940 ;
        RECT 1409.970 1089.740 1410.290 1089.800 ;
        RECT 1541.990 1089.740 1542.310 1089.800 ;
        RECT 1567.765 16.560 1568.055 16.605 ;
        RECT 1632.150 16.560 1632.470 16.620 ;
        RECT 1567.765 16.420 1632.470 16.560 ;
        RECT 1567.765 16.375 1568.055 16.420 ;
        RECT 1632.150 16.360 1632.470 16.420 ;
        RECT 1541.990 15.540 1542.310 15.600 ;
        RECT 1567.765 15.540 1568.055 15.585 ;
        RECT 1541.990 15.400 1568.055 15.540 ;
        RECT 1541.990 15.340 1542.310 15.400 ;
        RECT 1567.765 15.355 1568.055 15.400 ;
      LAYER via ;
        RECT 1410.000 1089.740 1410.260 1090.000 ;
        RECT 1542.020 1089.740 1542.280 1090.000 ;
        RECT 1632.180 16.360 1632.440 16.620 ;
        RECT 1542.020 15.340 1542.280 15.600 ;
      LAYER met2 ;
        RECT 1409.910 1100.580 1410.190 1104.000 ;
        RECT 1409.910 1100.000 1410.200 1100.580 ;
        RECT 1410.060 1090.030 1410.200 1100.000 ;
        RECT 1410.000 1089.710 1410.260 1090.030 ;
        RECT 1542.020 1089.710 1542.280 1090.030 ;
        RECT 1542.080 15.630 1542.220 1089.710 ;
        RECT 1632.180 16.330 1632.440 16.650 ;
        RECT 1542.020 15.310 1542.280 15.630 ;
        RECT 1632.240 2.000 1632.380 16.330 ;
        RECT 1632.030 -4.000 1632.590 2.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1415.950 1089.600 1416.270 1089.660 ;
        RECT 1420.550 1089.600 1420.870 1089.660 ;
        RECT 1415.950 1089.460 1420.870 1089.600 ;
        RECT 1415.950 1089.400 1416.270 1089.460 ;
        RECT 1420.550 1089.400 1420.870 1089.460 ;
        RECT 1420.550 193.500 1420.870 193.760 ;
        RECT 1420.640 193.080 1420.780 193.500 ;
        RECT 1420.550 192.820 1420.870 193.080 ;
        RECT 1420.550 169.020 1420.870 169.280 ;
        RECT 1420.640 168.600 1420.780 169.020 ;
        RECT 1420.550 168.340 1420.870 168.600 ;
        RECT 1420.550 22.000 1420.870 22.060 ;
        RECT 1650.090 22.000 1650.410 22.060 ;
        RECT 1420.550 21.860 1650.410 22.000 ;
        RECT 1420.550 21.800 1420.870 21.860 ;
        RECT 1650.090 21.800 1650.410 21.860 ;
      LAYER via ;
        RECT 1415.980 1089.400 1416.240 1089.660 ;
        RECT 1420.580 1089.400 1420.840 1089.660 ;
        RECT 1420.580 193.500 1420.840 193.760 ;
        RECT 1420.580 192.820 1420.840 193.080 ;
        RECT 1420.580 169.020 1420.840 169.280 ;
        RECT 1420.580 168.340 1420.840 168.600 ;
        RECT 1420.580 21.800 1420.840 22.060 ;
        RECT 1650.120 21.800 1650.380 22.060 ;
      LAYER met2 ;
        RECT 1415.890 1100.580 1416.170 1104.000 ;
        RECT 1415.890 1100.000 1416.180 1100.580 ;
        RECT 1416.040 1089.690 1416.180 1100.000 ;
        RECT 1415.980 1089.370 1416.240 1089.690 ;
        RECT 1420.580 1089.370 1420.840 1089.690 ;
        RECT 1420.640 193.790 1420.780 1089.370 ;
        RECT 1420.580 193.470 1420.840 193.790 ;
        RECT 1420.580 192.790 1420.840 193.110 ;
        RECT 1420.640 169.310 1420.780 192.790 ;
        RECT 1420.580 168.990 1420.840 169.310 ;
        RECT 1420.580 168.310 1420.840 168.630 ;
        RECT 1420.640 22.090 1420.780 168.310 ;
        RECT 1420.580 21.770 1420.840 22.090 ;
        RECT 1650.120 21.770 1650.380 22.090 ;
        RECT 1650.180 2.000 1650.320 21.770 ;
        RECT 1649.970 -4.000 1650.530 2.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1422.390 1089.600 1422.710 1089.660 ;
        RECT 1427.450 1089.600 1427.770 1089.660 ;
        RECT 1422.390 1089.460 1427.770 1089.600 ;
        RECT 1422.390 1089.400 1422.710 1089.460 ;
        RECT 1427.450 1089.400 1427.770 1089.460 ;
        RECT 1427.450 22.340 1427.770 22.400 ;
        RECT 1668.030 22.340 1668.350 22.400 ;
        RECT 1427.450 22.200 1668.350 22.340 ;
        RECT 1427.450 22.140 1427.770 22.200 ;
        RECT 1668.030 22.140 1668.350 22.200 ;
      LAYER via ;
        RECT 1422.420 1089.400 1422.680 1089.660 ;
        RECT 1427.480 1089.400 1427.740 1089.660 ;
        RECT 1427.480 22.140 1427.740 22.400 ;
        RECT 1668.060 22.140 1668.320 22.400 ;
      LAYER met2 ;
        RECT 1422.330 1100.580 1422.610 1104.000 ;
        RECT 1422.330 1100.000 1422.620 1100.580 ;
        RECT 1422.480 1089.690 1422.620 1100.000 ;
        RECT 1422.420 1089.370 1422.680 1089.690 ;
        RECT 1427.480 1089.370 1427.740 1089.690 ;
        RECT 1427.540 22.430 1427.680 1089.370 ;
        RECT 1427.480 22.110 1427.740 22.430 ;
        RECT 1668.060 22.110 1668.320 22.430 ;
        RECT 1668.120 2.000 1668.260 22.110 ;
        RECT 1667.910 -4.000 1668.470 2.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1428.370 1086.200 1428.690 1086.260 ;
        RECT 1434.350 1086.200 1434.670 1086.260 ;
        RECT 1428.370 1086.060 1434.670 1086.200 ;
        RECT 1428.370 1086.000 1428.690 1086.060 ;
        RECT 1434.350 1086.000 1434.670 1086.060 ;
        RECT 1434.350 23.360 1434.670 23.420 ;
        RECT 1685.510 23.360 1685.830 23.420 ;
        RECT 1434.350 23.220 1685.830 23.360 ;
        RECT 1434.350 23.160 1434.670 23.220 ;
        RECT 1685.510 23.160 1685.830 23.220 ;
      LAYER via ;
        RECT 1428.400 1086.000 1428.660 1086.260 ;
        RECT 1434.380 1086.000 1434.640 1086.260 ;
        RECT 1434.380 23.160 1434.640 23.420 ;
        RECT 1685.540 23.160 1685.800 23.420 ;
      LAYER met2 ;
        RECT 1428.310 1100.580 1428.590 1104.000 ;
        RECT 1428.310 1100.000 1428.600 1100.580 ;
        RECT 1428.460 1086.290 1428.600 1100.000 ;
        RECT 1428.400 1085.970 1428.660 1086.290 ;
        RECT 1434.380 1085.970 1434.640 1086.290 ;
        RECT 1434.440 23.450 1434.580 1085.970 ;
        RECT 1434.380 23.130 1434.640 23.450 ;
        RECT 1685.540 23.130 1685.800 23.450 ;
        RECT 1685.600 2.000 1685.740 23.130 ;
        RECT 1685.390 -4.000 1685.950 2.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 722.270 23.020 722.590 23.080 ;
        RECT 1097.170 23.020 1097.490 23.080 ;
        RECT 722.270 22.880 1097.490 23.020 ;
        RECT 722.270 22.820 722.590 22.880 ;
        RECT 1097.170 22.820 1097.490 22.880 ;
      LAYER via ;
        RECT 722.300 22.820 722.560 23.080 ;
        RECT 1097.200 22.820 1097.460 23.080 ;
      LAYER met2 ;
        RECT 1097.570 1100.650 1097.850 1104.000 ;
        RECT 1097.260 1100.510 1097.850 1100.650 ;
        RECT 1097.260 23.110 1097.400 1100.510 ;
        RECT 1097.570 1100.000 1097.850 1100.510 ;
        RECT 722.300 22.790 722.560 23.110 ;
        RECT 1097.200 22.790 1097.460 23.110 ;
        RECT 722.360 2.000 722.500 22.790 ;
        RECT 722.150 -4.000 722.710 2.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1433.890 27.100 1434.210 27.160 ;
        RECT 1703.450 27.100 1703.770 27.160 ;
        RECT 1433.890 26.960 1703.770 27.100 ;
        RECT 1433.890 26.900 1434.210 26.960 ;
        RECT 1703.450 26.900 1703.770 26.960 ;
      LAYER via ;
        RECT 1433.920 26.900 1434.180 27.160 ;
        RECT 1703.480 26.900 1703.740 27.160 ;
      LAYER met2 ;
        RECT 1434.290 1100.650 1434.570 1104.000 ;
        RECT 1433.980 1100.510 1434.570 1100.650 ;
        RECT 1433.980 27.190 1434.120 1100.510 ;
        RECT 1434.290 1100.000 1434.570 1100.510 ;
        RECT 1433.920 26.870 1434.180 27.190 ;
        RECT 1703.480 26.870 1703.740 27.190 ;
        RECT 1703.540 2.000 1703.680 26.870 ;
        RECT 1703.330 -4.000 1703.890 2.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1440.790 26.420 1441.110 26.480 ;
        RECT 1721.390 26.420 1721.710 26.480 ;
        RECT 1440.790 26.280 1721.710 26.420 ;
        RECT 1440.790 26.220 1441.110 26.280 ;
        RECT 1721.390 26.220 1721.710 26.280 ;
      LAYER via ;
        RECT 1440.820 26.220 1441.080 26.480 ;
        RECT 1721.420 26.220 1721.680 26.480 ;
      LAYER met2 ;
        RECT 1440.730 1100.580 1441.010 1104.000 ;
        RECT 1440.730 1100.000 1441.020 1100.580 ;
        RECT 1440.880 26.510 1441.020 1100.000 ;
        RECT 1440.820 26.190 1441.080 26.510 ;
        RECT 1721.420 26.190 1721.680 26.510 ;
        RECT 1721.480 2.000 1721.620 26.190 ;
        RECT 1721.270 -4.000 1721.830 2.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1446.770 1089.600 1447.090 1089.660 ;
        RECT 1448.610 1089.600 1448.930 1089.660 ;
        RECT 1446.770 1089.460 1448.930 1089.600 ;
        RECT 1446.770 1089.400 1447.090 1089.460 ;
        RECT 1448.610 1089.400 1448.930 1089.460 ;
        RECT 1448.610 26.080 1448.930 26.140 ;
        RECT 1739.330 26.080 1739.650 26.140 ;
        RECT 1448.610 25.940 1739.650 26.080 ;
        RECT 1448.610 25.880 1448.930 25.940 ;
        RECT 1739.330 25.880 1739.650 25.940 ;
      LAYER via ;
        RECT 1446.800 1089.400 1447.060 1089.660 ;
        RECT 1448.640 1089.400 1448.900 1089.660 ;
        RECT 1448.640 25.880 1448.900 26.140 ;
        RECT 1739.360 25.880 1739.620 26.140 ;
      LAYER met2 ;
        RECT 1446.710 1100.580 1446.990 1104.000 ;
        RECT 1446.710 1100.000 1447.000 1100.580 ;
        RECT 1446.860 1089.690 1447.000 1100.000 ;
        RECT 1446.800 1089.370 1447.060 1089.690 ;
        RECT 1448.640 1089.370 1448.900 1089.690 ;
        RECT 1448.700 26.170 1448.840 1089.370 ;
        RECT 1448.640 25.850 1448.900 26.170 ;
        RECT 1739.360 25.850 1739.620 26.170 ;
        RECT 1739.420 2.000 1739.560 25.850 ;
        RECT 1739.210 -4.000 1739.770 2.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1452.750 1089.600 1453.070 1089.660 ;
        RECT 1455.050 1089.600 1455.370 1089.660 ;
        RECT 1452.750 1089.460 1455.370 1089.600 ;
        RECT 1452.750 1089.400 1453.070 1089.460 ;
        RECT 1455.050 1089.400 1455.370 1089.460 ;
        RECT 1455.050 25.740 1455.370 25.800 ;
        RECT 1756.810 25.740 1757.130 25.800 ;
        RECT 1455.050 25.600 1757.130 25.740 ;
        RECT 1455.050 25.540 1455.370 25.600 ;
        RECT 1756.810 25.540 1757.130 25.600 ;
      LAYER via ;
        RECT 1452.780 1089.400 1453.040 1089.660 ;
        RECT 1455.080 1089.400 1455.340 1089.660 ;
        RECT 1455.080 25.540 1455.340 25.800 ;
        RECT 1756.840 25.540 1757.100 25.800 ;
      LAYER met2 ;
        RECT 1452.690 1100.580 1452.970 1104.000 ;
        RECT 1452.690 1100.000 1452.980 1100.580 ;
        RECT 1452.840 1089.690 1452.980 1100.000 ;
        RECT 1452.780 1089.370 1453.040 1089.690 ;
        RECT 1455.080 1089.370 1455.340 1089.690 ;
        RECT 1455.140 25.830 1455.280 1089.370 ;
        RECT 1455.080 25.510 1455.340 25.830 ;
        RECT 1756.840 25.510 1757.100 25.830 ;
        RECT 1756.900 2.000 1757.040 25.510 ;
        RECT 1756.690 -4.000 1757.250 2.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1459.190 1083.820 1459.510 1083.880 ;
        RECT 1461.950 1083.820 1462.270 1083.880 ;
        RECT 1459.190 1083.680 1462.270 1083.820 ;
        RECT 1459.190 1083.620 1459.510 1083.680 ;
        RECT 1461.950 1083.620 1462.270 1083.680 ;
        RECT 1461.950 25.400 1462.270 25.460 ;
        RECT 1774.750 25.400 1775.070 25.460 ;
        RECT 1461.950 25.260 1775.070 25.400 ;
        RECT 1461.950 25.200 1462.270 25.260 ;
        RECT 1774.750 25.200 1775.070 25.260 ;
      LAYER via ;
        RECT 1459.220 1083.620 1459.480 1083.880 ;
        RECT 1461.980 1083.620 1462.240 1083.880 ;
        RECT 1461.980 25.200 1462.240 25.460 ;
        RECT 1774.780 25.200 1775.040 25.460 ;
      LAYER met2 ;
        RECT 1459.130 1100.580 1459.410 1104.000 ;
        RECT 1459.130 1100.000 1459.420 1100.580 ;
        RECT 1459.280 1083.910 1459.420 1100.000 ;
        RECT 1459.220 1083.590 1459.480 1083.910 ;
        RECT 1461.980 1083.590 1462.240 1083.910 ;
        RECT 1462.040 25.490 1462.180 1083.590 ;
        RECT 1461.980 25.170 1462.240 25.490 ;
        RECT 1774.780 25.170 1775.040 25.490 ;
        RECT 1774.840 2.000 1774.980 25.170 ;
        RECT 1774.630 -4.000 1775.190 2.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1465.170 1085.520 1465.490 1085.580 ;
        RECT 1468.850 1085.520 1469.170 1085.580 ;
        RECT 1465.170 1085.380 1469.170 1085.520 ;
        RECT 1465.170 1085.320 1465.490 1085.380 ;
        RECT 1468.850 1085.320 1469.170 1085.380 ;
        RECT 1468.850 25.060 1469.170 25.120 ;
        RECT 1792.690 25.060 1793.010 25.120 ;
        RECT 1468.850 24.920 1793.010 25.060 ;
        RECT 1468.850 24.860 1469.170 24.920 ;
        RECT 1792.690 24.860 1793.010 24.920 ;
      LAYER via ;
        RECT 1465.200 1085.320 1465.460 1085.580 ;
        RECT 1468.880 1085.320 1469.140 1085.580 ;
        RECT 1468.880 24.860 1469.140 25.120 ;
        RECT 1792.720 24.860 1792.980 25.120 ;
      LAYER met2 ;
        RECT 1465.110 1100.580 1465.390 1104.000 ;
        RECT 1465.110 1100.000 1465.400 1100.580 ;
        RECT 1465.260 1085.610 1465.400 1100.000 ;
        RECT 1465.200 1085.290 1465.460 1085.610 ;
        RECT 1468.880 1085.290 1469.140 1085.610 ;
        RECT 1468.940 25.150 1469.080 1085.290 ;
        RECT 1468.880 24.830 1469.140 25.150 ;
        RECT 1792.720 24.830 1792.980 25.150 ;
        RECT 1792.780 2.000 1792.920 24.830 ;
        RECT 1792.570 -4.000 1793.130 2.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1471.150 1085.180 1471.470 1085.240 ;
        RECT 1476.210 1085.180 1476.530 1085.240 ;
        RECT 1471.150 1085.040 1476.530 1085.180 ;
        RECT 1471.150 1084.980 1471.470 1085.040 ;
        RECT 1476.210 1084.980 1476.530 1085.040 ;
        RECT 1476.210 24.720 1476.530 24.780 ;
        RECT 1810.630 24.720 1810.950 24.780 ;
        RECT 1476.210 24.580 1810.950 24.720 ;
        RECT 1476.210 24.520 1476.530 24.580 ;
        RECT 1810.630 24.520 1810.950 24.580 ;
      LAYER via ;
        RECT 1471.180 1084.980 1471.440 1085.240 ;
        RECT 1476.240 1084.980 1476.500 1085.240 ;
        RECT 1476.240 24.520 1476.500 24.780 ;
        RECT 1810.660 24.520 1810.920 24.780 ;
      LAYER met2 ;
        RECT 1471.090 1100.580 1471.370 1104.000 ;
        RECT 1471.090 1100.000 1471.380 1100.580 ;
        RECT 1471.240 1085.270 1471.380 1100.000 ;
        RECT 1471.180 1084.950 1471.440 1085.270 ;
        RECT 1476.240 1084.950 1476.500 1085.270 ;
        RECT 1476.300 24.810 1476.440 1084.950 ;
        RECT 1476.240 24.490 1476.500 24.810 ;
        RECT 1810.660 24.490 1810.920 24.810 ;
        RECT 1810.720 2.000 1810.860 24.490 ;
        RECT 1810.510 -4.000 1811.070 2.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1477.590 1088.240 1477.910 1088.300 ;
        RECT 1483.110 1088.240 1483.430 1088.300 ;
        RECT 1477.590 1088.100 1483.430 1088.240 ;
        RECT 1477.590 1088.040 1477.910 1088.100 ;
        RECT 1483.110 1088.040 1483.430 1088.100 ;
        RECT 1483.110 24.380 1483.430 24.440 ;
        RECT 1828.570 24.380 1828.890 24.440 ;
        RECT 1483.110 24.240 1828.890 24.380 ;
        RECT 1483.110 24.180 1483.430 24.240 ;
        RECT 1828.570 24.180 1828.890 24.240 ;
      LAYER via ;
        RECT 1477.620 1088.040 1477.880 1088.300 ;
        RECT 1483.140 1088.040 1483.400 1088.300 ;
        RECT 1483.140 24.180 1483.400 24.440 ;
        RECT 1828.600 24.180 1828.860 24.440 ;
      LAYER met2 ;
        RECT 1477.530 1100.580 1477.810 1104.000 ;
        RECT 1477.530 1100.000 1477.820 1100.580 ;
        RECT 1477.680 1088.330 1477.820 1100.000 ;
        RECT 1477.620 1088.010 1477.880 1088.330 ;
        RECT 1483.140 1088.010 1483.400 1088.330 ;
        RECT 1483.200 24.470 1483.340 1088.010 ;
        RECT 1483.140 24.150 1483.400 24.470 ;
        RECT 1828.600 24.150 1828.860 24.470 ;
        RECT 1828.660 2.000 1828.800 24.150 ;
        RECT 1828.450 -4.000 1829.010 2.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1483.570 1088.580 1483.890 1088.640 ;
        RECT 1490.010 1088.580 1490.330 1088.640 ;
        RECT 1483.570 1088.440 1490.330 1088.580 ;
        RECT 1483.570 1088.380 1483.890 1088.440 ;
        RECT 1490.010 1088.380 1490.330 1088.440 ;
        RECT 1490.010 24.040 1490.330 24.100 ;
        RECT 1846.050 24.040 1846.370 24.100 ;
        RECT 1490.010 23.900 1846.370 24.040 ;
        RECT 1490.010 23.840 1490.330 23.900 ;
        RECT 1846.050 23.840 1846.370 23.900 ;
      LAYER via ;
        RECT 1483.600 1088.380 1483.860 1088.640 ;
        RECT 1490.040 1088.380 1490.300 1088.640 ;
        RECT 1490.040 23.840 1490.300 24.100 ;
        RECT 1846.080 23.840 1846.340 24.100 ;
      LAYER met2 ;
        RECT 1483.510 1100.580 1483.790 1104.000 ;
        RECT 1483.510 1100.000 1483.800 1100.580 ;
        RECT 1483.660 1088.670 1483.800 1100.000 ;
        RECT 1483.600 1088.350 1483.860 1088.670 ;
        RECT 1490.040 1088.350 1490.300 1088.670 ;
        RECT 1490.100 24.130 1490.240 1088.350 ;
        RECT 1490.040 23.810 1490.300 24.130 ;
        RECT 1846.080 23.810 1846.340 24.130 ;
        RECT 1846.140 2.000 1846.280 23.810 ;
        RECT 1845.930 -4.000 1846.490 2.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1489.490 1100.580 1489.770 1104.000 ;
        RECT 1489.490 1100.000 1489.780 1100.580 ;
        RECT 1489.640 24.325 1489.780 1100.000 ;
        RECT 1489.570 23.955 1489.850 24.325 ;
        RECT 1864.010 23.955 1864.290 24.325 ;
        RECT 1864.080 2.000 1864.220 23.955 ;
        RECT 1863.870 -4.000 1864.430 2.000 ;
      LAYER via2 ;
        RECT 1489.570 24.000 1489.850 24.280 ;
        RECT 1864.010 24.000 1864.290 24.280 ;
      LAYER met3 ;
        RECT 1489.545 24.290 1489.875 24.305 ;
        RECT 1863.985 24.290 1864.315 24.305 ;
        RECT 1489.545 23.990 1864.315 24.290 ;
        RECT 1489.545 23.975 1489.875 23.990 ;
        RECT 1863.985 23.975 1864.315 23.990 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 740.210 22.680 740.530 22.740 ;
        RECT 1104.070 22.680 1104.390 22.740 ;
        RECT 740.210 22.540 1104.390 22.680 ;
        RECT 740.210 22.480 740.530 22.540 ;
        RECT 1104.070 22.480 1104.390 22.540 ;
      LAYER via ;
        RECT 740.240 22.480 740.500 22.740 ;
        RECT 1104.100 22.480 1104.360 22.740 ;
      LAYER met2 ;
        RECT 1104.010 1100.580 1104.290 1104.000 ;
        RECT 1104.010 1100.000 1104.300 1100.580 ;
        RECT 1104.160 22.770 1104.300 1100.000 ;
        RECT 740.240 22.450 740.500 22.770 ;
        RECT 1104.100 22.450 1104.360 22.770 ;
        RECT 740.300 2.000 740.440 22.450 ;
        RECT 740.090 -4.000 740.650 2.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1496.910 49.540 1497.230 49.600 ;
        RECT 1876.870 49.540 1877.190 49.600 ;
        RECT 1496.910 49.400 1877.190 49.540 ;
        RECT 1496.910 49.340 1497.230 49.400 ;
        RECT 1876.870 49.340 1877.190 49.400 ;
        RECT 1876.870 2.620 1877.190 2.680 ;
        RECT 1881.930 2.620 1882.250 2.680 ;
        RECT 1876.870 2.480 1882.250 2.620 ;
        RECT 1876.870 2.420 1877.190 2.480 ;
        RECT 1881.930 2.420 1882.250 2.480 ;
      LAYER via ;
        RECT 1496.940 49.340 1497.200 49.600 ;
        RECT 1876.900 49.340 1877.160 49.600 ;
        RECT 1876.900 2.420 1877.160 2.680 ;
        RECT 1881.960 2.420 1882.220 2.680 ;
      LAYER met2 ;
        RECT 1495.930 1100.650 1496.210 1104.000 ;
        RECT 1495.930 1100.510 1497.140 1100.650 ;
        RECT 1495.930 1100.000 1496.210 1100.510 ;
        RECT 1497.000 49.630 1497.140 1100.510 ;
        RECT 1496.940 49.310 1497.200 49.630 ;
        RECT 1876.900 49.310 1877.160 49.630 ;
        RECT 1876.960 2.710 1877.100 49.310 ;
        RECT 1876.900 2.390 1877.160 2.710 ;
        RECT 1881.960 2.390 1882.220 2.710 ;
        RECT 1882.020 2.000 1882.160 2.390 ;
        RECT 1881.810 -4.000 1882.370 2.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1501.970 1088.580 1502.290 1088.640 ;
        RECT 1503.810 1088.580 1504.130 1088.640 ;
        RECT 1501.970 1088.440 1504.130 1088.580 ;
        RECT 1501.970 1088.380 1502.290 1088.440 ;
        RECT 1503.810 1088.380 1504.130 1088.440 ;
        RECT 1503.810 49.880 1504.130 49.940 ;
        RECT 1897.570 49.880 1897.890 49.940 ;
        RECT 1503.810 49.740 1897.890 49.880 ;
        RECT 1503.810 49.680 1504.130 49.740 ;
        RECT 1897.570 49.680 1897.890 49.740 ;
      LAYER via ;
        RECT 1502.000 1088.380 1502.260 1088.640 ;
        RECT 1503.840 1088.380 1504.100 1088.640 ;
        RECT 1503.840 49.680 1504.100 49.940 ;
        RECT 1897.600 49.680 1897.860 49.940 ;
      LAYER met2 ;
        RECT 1501.910 1100.580 1502.190 1104.000 ;
        RECT 1501.910 1100.000 1502.200 1100.580 ;
        RECT 1502.060 1088.670 1502.200 1100.000 ;
        RECT 1502.000 1088.350 1502.260 1088.670 ;
        RECT 1503.840 1088.350 1504.100 1088.670 ;
        RECT 1503.900 49.970 1504.040 1088.350 ;
        RECT 1503.840 49.650 1504.100 49.970 ;
        RECT 1897.600 49.650 1897.860 49.970 ;
        RECT 1897.660 2.450 1897.800 49.650 ;
        RECT 1897.660 2.310 1900.100 2.450 ;
        RECT 1899.960 2.000 1900.100 2.310 ;
        RECT 1899.750 -4.000 1900.310 2.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1507.950 1088.580 1508.270 1088.640 ;
        RECT 1510.710 1088.580 1511.030 1088.640 ;
        RECT 1507.950 1088.440 1511.030 1088.580 ;
        RECT 1507.950 1088.380 1508.270 1088.440 ;
        RECT 1510.710 1088.380 1511.030 1088.440 ;
        RECT 1510.710 50.220 1511.030 50.280 ;
        RECT 1911.830 50.220 1912.150 50.280 ;
        RECT 1510.710 50.080 1912.150 50.220 ;
        RECT 1510.710 50.020 1511.030 50.080 ;
        RECT 1911.830 50.020 1912.150 50.080 ;
        RECT 1911.830 14.520 1912.150 14.580 ;
        RECT 1917.810 14.520 1918.130 14.580 ;
        RECT 1911.830 14.380 1918.130 14.520 ;
        RECT 1911.830 14.320 1912.150 14.380 ;
        RECT 1917.810 14.320 1918.130 14.380 ;
      LAYER via ;
        RECT 1507.980 1088.380 1508.240 1088.640 ;
        RECT 1510.740 1088.380 1511.000 1088.640 ;
        RECT 1510.740 50.020 1511.000 50.280 ;
        RECT 1911.860 50.020 1912.120 50.280 ;
        RECT 1911.860 14.320 1912.120 14.580 ;
        RECT 1917.840 14.320 1918.100 14.580 ;
      LAYER met2 ;
        RECT 1507.890 1100.580 1508.170 1104.000 ;
        RECT 1507.890 1100.000 1508.180 1100.580 ;
        RECT 1508.040 1088.670 1508.180 1100.000 ;
        RECT 1507.980 1088.350 1508.240 1088.670 ;
        RECT 1510.740 1088.350 1511.000 1088.670 ;
        RECT 1510.800 50.310 1510.940 1088.350 ;
        RECT 1510.740 49.990 1511.000 50.310 ;
        RECT 1911.860 49.990 1912.120 50.310 ;
        RECT 1911.920 14.610 1912.060 49.990 ;
        RECT 1911.860 14.290 1912.120 14.610 ;
        RECT 1917.840 14.290 1918.100 14.610 ;
        RECT 1917.900 2.000 1918.040 14.290 ;
        RECT 1917.690 -4.000 1918.250 2.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1513.930 1083.820 1514.250 1083.880 ;
        RECT 1517.610 1083.820 1517.930 1083.880 ;
        RECT 1513.930 1083.680 1517.930 1083.820 ;
        RECT 1513.930 1083.620 1514.250 1083.680 ;
        RECT 1517.610 1083.620 1517.930 1083.680 ;
        RECT 1517.610 50.560 1517.930 50.620 ;
        RECT 1932.070 50.560 1932.390 50.620 ;
        RECT 1517.610 50.420 1932.390 50.560 ;
        RECT 1517.610 50.360 1517.930 50.420 ;
        RECT 1932.070 50.360 1932.390 50.420 ;
      LAYER via ;
        RECT 1513.960 1083.620 1514.220 1083.880 ;
        RECT 1517.640 1083.620 1517.900 1083.880 ;
        RECT 1517.640 50.360 1517.900 50.620 ;
        RECT 1932.100 50.360 1932.360 50.620 ;
      LAYER met2 ;
        RECT 1513.870 1100.580 1514.150 1104.000 ;
        RECT 1513.870 1100.000 1514.160 1100.580 ;
        RECT 1514.020 1083.910 1514.160 1100.000 ;
        RECT 1513.960 1083.590 1514.220 1083.910 ;
        RECT 1517.640 1083.590 1517.900 1083.910 ;
        RECT 1517.700 50.650 1517.840 1083.590 ;
        RECT 1517.640 50.330 1517.900 50.650 ;
        RECT 1932.100 50.330 1932.360 50.650 ;
        RECT 1932.160 2.450 1932.300 50.330 ;
        RECT 1932.160 2.310 1935.520 2.450 ;
        RECT 1935.380 2.000 1935.520 2.310 ;
        RECT 1935.170 -4.000 1935.730 2.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1520.370 1083.820 1520.690 1083.880 ;
        RECT 1524.510 1083.820 1524.830 1083.880 ;
        RECT 1520.370 1083.680 1524.830 1083.820 ;
        RECT 1520.370 1083.620 1520.690 1083.680 ;
        RECT 1524.510 1083.620 1524.830 1083.680 ;
        RECT 1524.510 50.900 1524.830 50.960 ;
        RECT 1953.230 50.900 1953.550 50.960 ;
        RECT 1524.510 50.760 1953.550 50.900 ;
        RECT 1524.510 50.700 1524.830 50.760 ;
        RECT 1953.230 50.700 1953.550 50.760 ;
      LAYER via ;
        RECT 1520.400 1083.620 1520.660 1083.880 ;
        RECT 1524.540 1083.620 1524.800 1083.880 ;
        RECT 1524.540 50.700 1524.800 50.960 ;
        RECT 1953.260 50.700 1953.520 50.960 ;
      LAYER met2 ;
        RECT 1520.310 1100.580 1520.590 1104.000 ;
        RECT 1520.310 1100.000 1520.600 1100.580 ;
        RECT 1520.460 1083.910 1520.600 1100.000 ;
        RECT 1520.400 1083.590 1520.660 1083.910 ;
        RECT 1524.540 1083.590 1524.800 1083.910 ;
        RECT 1524.600 50.990 1524.740 1083.590 ;
        RECT 1524.540 50.670 1524.800 50.990 ;
        RECT 1953.260 50.670 1953.520 50.990 ;
        RECT 1953.320 2.000 1953.460 50.670 ;
        RECT 1953.110 -4.000 1953.670 2.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1526.350 1083.820 1526.670 1083.880 ;
        RECT 1530.950 1083.820 1531.270 1083.880 ;
        RECT 1526.350 1083.680 1531.270 1083.820 ;
        RECT 1526.350 1083.620 1526.670 1083.680 ;
        RECT 1530.950 1083.620 1531.270 1083.680 ;
        RECT 1530.950 51.240 1531.270 51.300 ;
        RECT 1966.570 51.240 1966.890 51.300 ;
        RECT 1530.950 51.100 1966.890 51.240 ;
        RECT 1530.950 51.040 1531.270 51.100 ;
        RECT 1966.570 51.040 1966.890 51.100 ;
      LAYER via ;
        RECT 1526.380 1083.620 1526.640 1083.880 ;
        RECT 1530.980 1083.620 1531.240 1083.880 ;
        RECT 1530.980 51.040 1531.240 51.300 ;
        RECT 1966.600 51.040 1966.860 51.300 ;
      LAYER met2 ;
        RECT 1526.290 1100.580 1526.570 1104.000 ;
        RECT 1526.290 1100.000 1526.580 1100.580 ;
        RECT 1526.440 1083.910 1526.580 1100.000 ;
        RECT 1526.380 1083.590 1526.640 1083.910 ;
        RECT 1530.980 1083.590 1531.240 1083.910 ;
        RECT 1531.040 51.330 1531.180 1083.590 ;
        RECT 1530.980 51.010 1531.240 51.330 ;
        RECT 1966.600 51.010 1966.860 51.330 ;
        RECT 1966.660 16.730 1966.800 51.010 ;
        RECT 1966.660 16.590 1971.400 16.730 ;
        RECT 1971.260 2.000 1971.400 16.590 ;
        RECT 1971.050 -4.000 1971.610 2.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1532.330 1083.820 1532.650 1083.880 ;
        RECT 1537.850 1083.820 1538.170 1083.880 ;
        RECT 1532.330 1083.680 1538.170 1083.820 ;
        RECT 1532.330 1083.620 1532.650 1083.680 ;
        RECT 1537.850 1083.620 1538.170 1083.680 ;
        RECT 1537.850 54.980 1538.170 55.040 ;
        RECT 1987.270 54.980 1987.590 55.040 ;
        RECT 1537.850 54.840 1987.590 54.980 ;
        RECT 1537.850 54.780 1538.170 54.840 ;
        RECT 1987.270 54.780 1987.590 54.840 ;
      LAYER via ;
        RECT 1532.360 1083.620 1532.620 1083.880 ;
        RECT 1537.880 1083.620 1538.140 1083.880 ;
        RECT 1537.880 54.780 1538.140 55.040 ;
        RECT 1987.300 54.780 1987.560 55.040 ;
      LAYER met2 ;
        RECT 1532.270 1100.580 1532.550 1104.000 ;
        RECT 1532.270 1100.000 1532.560 1100.580 ;
        RECT 1532.420 1083.910 1532.560 1100.000 ;
        RECT 1532.360 1083.590 1532.620 1083.910 ;
        RECT 1537.880 1083.590 1538.140 1083.910 ;
        RECT 1537.940 55.070 1538.080 1083.590 ;
        RECT 1537.880 54.750 1538.140 55.070 ;
        RECT 1987.300 54.750 1987.560 55.070 ;
        RECT 1987.360 16.730 1987.500 54.750 ;
        RECT 1987.360 16.590 1989.340 16.730 ;
        RECT 1989.200 2.000 1989.340 16.590 ;
        RECT 1988.990 -4.000 1989.550 2.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1538.770 1083.820 1539.090 1083.880 ;
        RECT 1544.290 1083.820 1544.610 1083.880 ;
        RECT 1538.770 1083.680 1544.610 1083.820 ;
        RECT 1538.770 1083.620 1539.090 1083.680 ;
        RECT 1544.290 1083.620 1544.610 1083.680 ;
        RECT 1544.290 54.640 1544.610 54.700 ;
        RECT 2001.530 54.640 2001.850 54.700 ;
        RECT 1544.290 54.500 2001.850 54.640 ;
        RECT 1544.290 54.440 1544.610 54.500 ;
        RECT 2001.530 54.440 2001.850 54.500 ;
      LAYER via ;
        RECT 1538.800 1083.620 1539.060 1083.880 ;
        RECT 1544.320 1083.620 1544.580 1083.880 ;
        RECT 1544.320 54.440 1544.580 54.700 ;
        RECT 2001.560 54.440 2001.820 54.700 ;
      LAYER met2 ;
        RECT 1538.710 1100.580 1538.990 1104.000 ;
        RECT 1538.710 1100.000 1539.000 1100.580 ;
        RECT 1538.860 1083.910 1539.000 1100.000 ;
        RECT 1538.800 1083.590 1539.060 1083.910 ;
        RECT 1544.320 1083.590 1544.580 1083.910 ;
        RECT 1544.380 54.730 1544.520 1083.590 ;
        RECT 1544.320 54.410 1544.580 54.730 ;
        RECT 2001.560 54.410 2001.820 54.730 ;
        RECT 2001.620 16.730 2001.760 54.410 ;
        RECT 2001.620 16.590 2006.820 16.730 ;
        RECT 2006.680 2.000 2006.820 16.590 ;
        RECT 2006.470 -4.000 2007.030 2.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1545.210 27.780 1545.530 27.840 ;
        RECT 2024.530 27.780 2024.850 27.840 ;
        RECT 1545.210 27.640 2024.850 27.780 ;
        RECT 1545.210 27.580 1545.530 27.640 ;
        RECT 2024.530 27.580 2024.850 27.640 ;
      LAYER via ;
        RECT 1545.240 27.580 1545.500 27.840 ;
        RECT 2024.560 27.580 2024.820 27.840 ;
      LAYER met2 ;
        RECT 1544.690 1100.650 1544.970 1104.000 ;
        RECT 1544.690 1100.510 1545.440 1100.650 ;
        RECT 1544.690 1100.000 1544.970 1100.510 ;
        RECT 1545.300 27.870 1545.440 1100.510 ;
        RECT 1545.240 27.550 1545.500 27.870 ;
        RECT 2024.560 27.550 2024.820 27.870 ;
        RECT 2024.620 2.000 2024.760 27.550 ;
        RECT 2024.410 -4.000 2024.970 2.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1552.110 28.120 1552.430 28.180 ;
        RECT 2042.470 28.120 2042.790 28.180 ;
        RECT 1552.110 27.980 2042.790 28.120 ;
        RECT 1552.110 27.920 1552.430 27.980 ;
        RECT 2042.470 27.920 2042.790 27.980 ;
      LAYER via ;
        RECT 1552.140 27.920 1552.400 28.180 ;
        RECT 2042.500 27.920 2042.760 28.180 ;
      LAYER met2 ;
        RECT 1550.670 1100.650 1550.950 1104.000 ;
        RECT 1550.670 1100.510 1552.340 1100.650 ;
        RECT 1550.670 1100.000 1550.950 1100.510 ;
        RECT 1552.200 28.210 1552.340 1100.510 ;
        RECT 1552.140 27.890 1552.400 28.210 ;
        RECT 2042.500 27.890 2042.760 28.210 ;
        RECT 2042.560 2.000 2042.700 27.890 ;
        RECT 2042.350 -4.000 2042.910 2.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1104.530 1052.540 1104.850 1052.600 ;
        RECT 1108.670 1052.540 1108.990 1052.600 ;
        RECT 1104.530 1052.400 1108.990 1052.540 ;
        RECT 1104.530 1052.340 1104.850 1052.400 ;
        RECT 1108.670 1052.340 1108.990 1052.400 ;
        RECT 757.690 22.340 758.010 22.400 ;
        RECT 1104.530 22.340 1104.850 22.400 ;
        RECT 757.690 22.200 1104.850 22.340 ;
        RECT 757.690 22.140 758.010 22.200 ;
        RECT 1104.530 22.140 1104.850 22.200 ;
      LAYER via ;
        RECT 1104.560 1052.340 1104.820 1052.600 ;
        RECT 1108.700 1052.340 1108.960 1052.600 ;
        RECT 757.720 22.140 757.980 22.400 ;
        RECT 1104.560 22.140 1104.820 22.400 ;
      LAYER met2 ;
        RECT 1109.990 1100.650 1110.270 1104.000 ;
        RECT 1108.760 1100.510 1110.270 1100.650 ;
        RECT 1108.760 1052.630 1108.900 1100.510 ;
        RECT 1109.990 1100.000 1110.270 1100.510 ;
        RECT 1104.560 1052.310 1104.820 1052.630 ;
        RECT 1108.700 1052.310 1108.960 1052.630 ;
        RECT 1104.620 22.430 1104.760 1052.310 ;
        RECT 757.720 22.110 757.980 22.430 ;
        RECT 1104.560 22.110 1104.820 22.430 ;
        RECT 757.780 2.000 757.920 22.110 ;
        RECT 757.570 -4.000 758.130 2.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1557.170 1083.820 1557.490 1083.880 ;
        RECT 1559.010 1083.820 1559.330 1083.880 ;
        RECT 1557.170 1083.680 1559.330 1083.820 ;
        RECT 1557.170 1083.620 1557.490 1083.680 ;
        RECT 1559.010 1083.620 1559.330 1083.680 ;
        RECT 1559.010 28.460 1559.330 28.520 ;
        RECT 2060.410 28.460 2060.730 28.520 ;
        RECT 1559.010 28.320 2060.730 28.460 ;
        RECT 1559.010 28.260 1559.330 28.320 ;
        RECT 2060.410 28.260 2060.730 28.320 ;
      LAYER via ;
        RECT 1557.200 1083.620 1557.460 1083.880 ;
        RECT 1559.040 1083.620 1559.300 1083.880 ;
        RECT 1559.040 28.260 1559.300 28.520 ;
        RECT 2060.440 28.260 2060.700 28.520 ;
      LAYER met2 ;
        RECT 1557.110 1100.580 1557.390 1104.000 ;
        RECT 1557.110 1100.000 1557.400 1100.580 ;
        RECT 1557.260 1083.910 1557.400 1100.000 ;
        RECT 1557.200 1083.590 1557.460 1083.910 ;
        RECT 1559.040 1083.590 1559.300 1083.910 ;
        RECT 1559.100 28.550 1559.240 1083.590 ;
        RECT 1559.040 28.230 1559.300 28.550 ;
        RECT 2060.440 28.230 2060.700 28.550 ;
        RECT 2060.500 2.000 2060.640 28.230 ;
        RECT 2060.290 -4.000 2060.850 2.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1563.150 1083.480 1563.470 1083.540 ;
        RECT 1565.910 1083.480 1566.230 1083.540 ;
        RECT 1563.150 1083.340 1566.230 1083.480 ;
        RECT 1563.150 1083.280 1563.470 1083.340 ;
        RECT 1565.910 1083.280 1566.230 1083.340 ;
        RECT 1565.910 28.800 1566.230 28.860 ;
        RECT 2078.350 28.800 2078.670 28.860 ;
        RECT 1565.910 28.660 2078.670 28.800 ;
        RECT 1565.910 28.600 1566.230 28.660 ;
        RECT 2078.350 28.600 2078.670 28.660 ;
      LAYER via ;
        RECT 1563.180 1083.280 1563.440 1083.540 ;
        RECT 1565.940 1083.280 1566.200 1083.540 ;
        RECT 1565.940 28.600 1566.200 28.860 ;
        RECT 2078.380 28.600 2078.640 28.860 ;
      LAYER met2 ;
        RECT 1563.090 1100.580 1563.370 1104.000 ;
        RECT 1563.090 1100.000 1563.380 1100.580 ;
        RECT 1563.240 1083.570 1563.380 1100.000 ;
        RECT 1563.180 1083.250 1563.440 1083.570 ;
        RECT 1565.940 1083.250 1566.200 1083.570 ;
        RECT 1566.000 28.890 1566.140 1083.250 ;
        RECT 1565.940 28.570 1566.200 28.890 ;
        RECT 2078.380 28.570 2078.640 28.890 ;
        RECT 2078.440 2.000 2078.580 28.570 ;
        RECT 2078.230 -4.000 2078.790 2.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1569.130 1086.200 1569.450 1086.260 ;
        RECT 1572.810 1086.200 1573.130 1086.260 ;
        RECT 1569.130 1086.060 1573.130 1086.200 ;
        RECT 1569.130 1086.000 1569.450 1086.060 ;
        RECT 1572.810 1086.000 1573.130 1086.060 ;
        RECT 1572.810 29.140 1573.130 29.200 ;
        RECT 2095.830 29.140 2096.150 29.200 ;
        RECT 1572.810 29.000 2096.150 29.140 ;
        RECT 1572.810 28.940 1573.130 29.000 ;
        RECT 2095.830 28.940 2096.150 29.000 ;
      LAYER via ;
        RECT 1569.160 1086.000 1569.420 1086.260 ;
        RECT 1572.840 1086.000 1573.100 1086.260 ;
        RECT 1572.840 28.940 1573.100 29.200 ;
        RECT 2095.860 28.940 2096.120 29.200 ;
      LAYER met2 ;
        RECT 1569.070 1100.580 1569.350 1104.000 ;
        RECT 1569.070 1100.000 1569.360 1100.580 ;
        RECT 1569.220 1086.290 1569.360 1100.000 ;
        RECT 1569.160 1085.970 1569.420 1086.290 ;
        RECT 1572.840 1085.970 1573.100 1086.290 ;
        RECT 1572.900 29.230 1573.040 1085.970 ;
        RECT 1572.840 28.910 1573.100 29.230 ;
        RECT 2095.860 28.910 2096.120 29.230 ;
        RECT 2095.920 2.000 2096.060 28.910 ;
        RECT 2095.710 -4.000 2096.270 2.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1575.570 1083.480 1575.890 1083.540 ;
        RECT 1579.710 1083.480 1580.030 1083.540 ;
        RECT 1575.570 1083.340 1580.030 1083.480 ;
        RECT 1575.570 1083.280 1575.890 1083.340 ;
        RECT 1579.710 1083.280 1580.030 1083.340 ;
        RECT 1579.710 29.480 1580.030 29.540 ;
        RECT 2113.770 29.480 2114.090 29.540 ;
        RECT 1579.710 29.340 2114.090 29.480 ;
        RECT 1579.710 29.280 1580.030 29.340 ;
        RECT 2113.770 29.280 2114.090 29.340 ;
      LAYER via ;
        RECT 1575.600 1083.280 1575.860 1083.540 ;
        RECT 1579.740 1083.280 1580.000 1083.540 ;
        RECT 1579.740 29.280 1580.000 29.540 ;
        RECT 2113.800 29.280 2114.060 29.540 ;
      LAYER met2 ;
        RECT 1575.510 1100.580 1575.790 1104.000 ;
        RECT 1575.510 1100.000 1575.800 1100.580 ;
        RECT 1575.660 1083.570 1575.800 1100.000 ;
        RECT 1575.600 1083.250 1575.860 1083.570 ;
        RECT 1579.740 1083.250 1580.000 1083.570 ;
        RECT 1579.800 29.570 1579.940 1083.250 ;
        RECT 1579.740 29.250 1580.000 29.570 ;
        RECT 2113.800 29.250 2114.060 29.570 ;
        RECT 2113.860 2.000 2114.000 29.250 ;
        RECT 2113.650 -4.000 2114.210 2.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1581.550 1083.480 1581.870 1083.540 ;
        RECT 1586.610 1083.480 1586.930 1083.540 ;
        RECT 1581.550 1083.340 1586.930 1083.480 ;
        RECT 1581.550 1083.280 1581.870 1083.340 ;
        RECT 1586.610 1083.280 1586.930 1083.340 ;
        RECT 1586.610 29.820 1586.930 29.880 ;
        RECT 2131.710 29.820 2132.030 29.880 ;
        RECT 1586.610 29.680 2132.030 29.820 ;
        RECT 1586.610 29.620 1586.930 29.680 ;
        RECT 2131.710 29.620 2132.030 29.680 ;
      LAYER via ;
        RECT 1581.580 1083.280 1581.840 1083.540 ;
        RECT 1586.640 1083.280 1586.900 1083.540 ;
        RECT 1586.640 29.620 1586.900 29.880 ;
        RECT 2131.740 29.620 2132.000 29.880 ;
      LAYER met2 ;
        RECT 1581.490 1100.580 1581.770 1104.000 ;
        RECT 1581.490 1100.000 1581.780 1100.580 ;
        RECT 1581.640 1083.570 1581.780 1100.000 ;
        RECT 1581.580 1083.250 1581.840 1083.570 ;
        RECT 1586.640 1083.250 1586.900 1083.570 ;
        RECT 1586.700 29.910 1586.840 1083.250 ;
        RECT 1586.640 29.590 1586.900 29.910 ;
        RECT 2131.740 29.590 2132.000 29.910 ;
        RECT 2131.800 2.000 2131.940 29.590 ;
        RECT 2131.590 -4.000 2132.150 2.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1587.530 1083.480 1587.850 1083.540 ;
        RECT 1593.050 1083.480 1593.370 1083.540 ;
        RECT 1587.530 1083.340 1593.370 1083.480 ;
        RECT 1587.530 1083.280 1587.850 1083.340 ;
        RECT 1593.050 1083.280 1593.370 1083.340 ;
        RECT 1593.050 30.160 1593.370 30.220 ;
        RECT 2149.650 30.160 2149.970 30.220 ;
        RECT 1593.050 30.020 2149.970 30.160 ;
        RECT 1593.050 29.960 1593.370 30.020 ;
        RECT 2149.650 29.960 2149.970 30.020 ;
      LAYER via ;
        RECT 1587.560 1083.280 1587.820 1083.540 ;
        RECT 1593.080 1083.280 1593.340 1083.540 ;
        RECT 1593.080 29.960 1593.340 30.220 ;
        RECT 2149.680 29.960 2149.940 30.220 ;
      LAYER met2 ;
        RECT 1587.470 1100.580 1587.750 1104.000 ;
        RECT 1587.470 1100.000 1587.760 1100.580 ;
        RECT 1587.620 1083.570 1587.760 1100.000 ;
        RECT 1587.560 1083.250 1587.820 1083.570 ;
        RECT 1593.080 1083.250 1593.340 1083.570 ;
        RECT 1593.140 30.250 1593.280 1083.250 ;
        RECT 1593.080 29.930 1593.340 30.250 ;
        RECT 2149.680 29.930 2149.940 30.250 ;
        RECT 2149.740 2.000 2149.880 29.930 ;
        RECT 2149.530 -4.000 2150.090 2.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1593.510 30.500 1593.830 30.560 ;
        RECT 2167.590 30.500 2167.910 30.560 ;
        RECT 1593.510 30.360 2167.910 30.500 ;
        RECT 1593.510 30.300 1593.830 30.360 ;
        RECT 2167.590 30.300 2167.910 30.360 ;
      LAYER via ;
        RECT 1593.540 30.300 1593.800 30.560 ;
        RECT 2167.620 30.300 2167.880 30.560 ;
      LAYER met2 ;
        RECT 1593.450 1100.580 1593.730 1104.000 ;
        RECT 1593.450 1100.000 1593.740 1100.580 ;
        RECT 1593.600 30.590 1593.740 1100.000 ;
        RECT 1593.540 30.270 1593.800 30.590 ;
        RECT 2167.620 30.270 2167.880 30.590 ;
        RECT 2167.680 2.000 2167.820 30.270 ;
        RECT 2167.470 -4.000 2168.030 2.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1600.410 34.240 1600.730 34.300 ;
        RECT 2185.070 34.240 2185.390 34.300 ;
        RECT 1600.410 34.100 2185.390 34.240 ;
        RECT 1600.410 34.040 1600.730 34.100 ;
        RECT 2185.070 34.040 2185.390 34.100 ;
      LAYER via ;
        RECT 1600.440 34.040 1600.700 34.300 ;
        RECT 2185.100 34.040 2185.360 34.300 ;
      LAYER met2 ;
        RECT 1599.890 1100.650 1600.170 1104.000 ;
        RECT 1599.890 1100.510 1600.640 1100.650 ;
        RECT 1599.890 1100.000 1600.170 1100.510 ;
        RECT 1600.500 34.330 1600.640 1100.510 ;
        RECT 1600.440 34.010 1600.700 34.330 ;
        RECT 2185.100 34.010 2185.360 34.330 ;
        RECT 2185.160 2.000 2185.300 34.010 ;
        RECT 2184.950 -4.000 2185.510 2.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1607.310 33.900 1607.630 33.960 ;
        RECT 2203.010 33.900 2203.330 33.960 ;
        RECT 1607.310 33.760 2203.330 33.900 ;
        RECT 1607.310 33.700 1607.630 33.760 ;
        RECT 2203.010 33.700 2203.330 33.760 ;
      LAYER via ;
        RECT 1607.340 33.700 1607.600 33.960 ;
        RECT 2203.040 33.700 2203.300 33.960 ;
      LAYER met2 ;
        RECT 1605.870 1100.650 1606.150 1104.000 ;
        RECT 1605.870 1100.510 1607.540 1100.650 ;
        RECT 1605.870 1100.000 1606.150 1100.510 ;
        RECT 1607.400 33.990 1607.540 1100.510 ;
        RECT 1607.340 33.670 1607.600 33.990 ;
        RECT 2203.040 33.670 2203.300 33.990 ;
        RECT 2203.100 2.000 2203.240 33.670 ;
        RECT 2202.890 -4.000 2203.450 2.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1611.910 1087.900 1612.230 1087.960 ;
        RECT 1614.210 1087.900 1614.530 1087.960 ;
        RECT 1611.910 1087.760 1614.530 1087.900 ;
        RECT 1611.910 1087.700 1612.230 1087.760 ;
        RECT 1614.210 1087.700 1614.530 1087.760 ;
        RECT 1614.210 33.560 1614.530 33.620 ;
        RECT 2220.950 33.560 2221.270 33.620 ;
        RECT 1614.210 33.420 2221.270 33.560 ;
        RECT 1614.210 33.360 1614.530 33.420 ;
        RECT 2220.950 33.360 2221.270 33.420 ;
      LAYER via ;
        RECT 1611.940 1087.700 1612.200 1087.960 ;
        RECT 1614.240 1087.700 1614.500 1087.960 ;
        RECT 1614.240 33.360 1614.500 33.620 ;
        RECT 2220.980 33.360 2221.240 33.620 ;
      LAYER met2 ;
        RECT 1611.850 1100.580 1612.130 1104.000 ;
        RECT 1611.850 1100.000 1612.140 1100.580 ;
        RECT 1612.000 1087.990 1612.140 1100.000 ;
        RECT 1611.940 1087.670 1612.200 1087.990 ;
        RECT 1614.240 1087.670 1614.500 1087.990 ;
        RECT 1614.300 33.650 1614.440 1087.670 ;
        RECT 1614.240 33.330 1614.500 33.650 ;
        RECT 2220.980 33.330 2221.240 33.650 ;
        RECT 2221.040 2.000 2221.180 33.330 ;
        RECT 2220.830 -4.000 2221.390 2.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1110.970 1032.480 1111.290 1032.540 ;
        RECT 1114.650 1032.480 1114.970 1032.540 ;
        RECT 1110.970 1032.340 1114.970 1032.480 ;
        RECT 1110.970 1032.280 1111.290 1032.340 ;
        RECT 1114.650 1032.280 1114.970 1032.340 ;
        RECT 775.630 22.000 775.950 22.060 ;
        RECT 1110.970 22.000 1111.290 22.060 ;
        RECT 775.630 21.860 1111.290 22.000 ;
        RECT 775.630 21.800 775.950 21.860 ;
        RECT 1110.970 21.800 1111.290 21.860 ;
      LAYER via ;
        RECT 1111.000 1032.280 1111.260 1032.540 ;
        RECT 1114.680 1032.280 1114.940 1032.540 ;
        RECT 775.660 21.800 775.920 22.060 ;
        RECT 1111.000 21.800 1111.260 22.060 ;
      LAYER met2 ;
        RECT 1115.970 1100.650 1116.250 1104.000 ;
        RECT 1114.740 1100.510 1116.250 1100.650 ;
        RECT 1114.740 1032.570 1114.880 1100.510 ;
        RECT 1115.970 1100.000 1116.250 1100.510 ;
        RECT 1111.000 1032.250 1111.260 1032.570 ;
        RECT 1114.680 1032.250 1114.940 1032.570 ;
        RECT 1111.060 22.090 1111.200 1032.250 ;
        RECT 775.660 21.770 775.920 22.090 ;
        RECT 1111.000 21.770 1111.260 22.090 ;
        RECT 775.720 2.000 775.860 21.770 ;
        RECT 775.510 -4.000 776.070 2.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1618.350 1087.560 1618.670 1087.620 ;
        RECT 1621.110 1087.560 1621.430 1087.620 ;
        RECT 1618.350 1087.420 1621.430 1087.560 ;
        RECT 1618.350 1087.360 1618.670 1087.420 ;
        RECT 1621.110 1087.360 1621.430 1087.420 ;
        RECT 1621.110 33.220 1621.430 33.280 ;
        RECT 2238.890 33.220 2239.210 33.280 ;
        RECT 1621.110 33.080 2239.210 33.220 ;
        RECT 1621.110 33.020 1621.430 33.080 ;
        RECT 2238.890 33.020 2239.210 33.080 ;
      LAYER via ;
        RECT 1618.380 1087.360 1618.640 1087.620 ;
        RECT 1621.140 1087.360 1621.400 1087.620 ;
        RECT 1621.140 33.020 1621.400 33.280 ;
        RECT 2238.920 33.020 2239.180 33.280 ;
      LAYER met2 ;
        RECT 1618.290 1100.580 1618.570 1104.000 ;
        RECT 1618.290 1100.000 1618.580 1100.580 ;
        RECT 1618.440 1087.650 1618.580 1100.000 ;
        RECT 1618.380 1087.330 1618.640 1087.650 ;
        RECT 1621.140 1087.330 1621.400 1087.650 ;
        RECT 1621.200 33.310 1621.340 1087.330 ;
        RECT 1621.140 32.990 1621.400 33.310 ;
        RECT 2238.920 32.990 2239.180 33.310 ;
        RECT 2238.980 2.000 2239.120 32.990 ;
        RECT 2238.770 -4.000 2239.330 2.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1624.330 1087.900 1624.650 1087.960 ;
        RECT 1628.010 1087.900 1628.330 1087.960 ;
        RECT 1624.330 1087.760 1628.330 1087.900 ;
        RECT 1624.330 1087.700 1624.650 1087.760 ;
        RECT 1628.010 1087.700 1628.330 1087.760 ;
        RECT 1628.010 32.880 1628.330 32.940 ;
        RECT 2256.370 32.880 2256.690 32.940 ;
        RECT 1628.010 32.740 2256.690 32.880 ;
        RECT 1628.010 32.680 1628.330 32.740 ;
        RECT 2256.370 32.680 2256.690 32.740 ;
      LAYER via ;
        RECT 1624.360 1087.700 1624.620 1087.960 ;
        RECT 1628.040 1087.700 1628.300 1087.960 ;
        RECT 1628.040 32.680 1628.300 32.940 ;
        RECT 2256.400 32.680 2256.660 32.940 ;
      LAYER met2 ;
        RECT 1624.270 1100.580 1624.550 1104.000 ;
        RECT 1624.270 1100.000 1624.560 1100.580 ;
        RECT 1624.420 1087.990 1624.560 1100.000 ;
        RECT 1624.360 1087.670 1624.620 1087.990 ;
        RECT 1628.040 1087.670 1628.300 1087.990 ;
        RECT 1628.100 32.970 1628.240 1087.670 ;
        RECT 1628.040 32.650 1628.300 32.970 ;
        RECT 2256.400 32.650 2256.660 32.970 ;
        RECT 2256.460 2.000 2256.600 32.650 ;
        RECT 2256.250 -4.000 2256.810 2.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1630.310 1087.900 1630.630 1087.960 ;
        RECT 1634.910 1087.900 1635.230 1087.960 ;
        RECT 1630.310 1087.760 1635.230 1087.900 ;
        RECT 1630.310 1087.700 1630.630 1087.760 ;
        RECT 1634.910 1087.700 1635.230 1087.760 ;
        RECT 1634.910 32.540 1635.230 32.600 ;
        RECT 2274.310 32.540 2274.630 32.600 ;
        RECT 1634.910 32.400 2274.630 32.540 ;
        RECT 1634.910 32.340 1635.230 32.400 ;
        RECT 2274.310 32.340 2274.630 32.400 ;
      LAYER via ;
        RECT 1630.340 1087.700 1630.600 1087.960 ;
        RECT 1634.940 1087.700 1635.200 1087.960 ;
        RECT 1634.940 32.340 1635.200 32.600 ;
        RECT 2274.340 32.340 2274.600 32.600 ;
      LAYER met2 ;
        RECT 1630.250 1100.580 1630.530 1104.000 ;
        RECT 1630.250 1100.000 1630.540 1100.580 ;
        RECT 1630.400 1087.990 1630.540 1100.000 ;
        RECT 1630.340 1087.670 1630.600 1087.990 ;
        RECT 1634.940 1087.670 1635.200 1087.990 ;
        RECT 1635.000 32.630 1635.140 1087.670 ;
        RECT 1634.940 32.310 1635.200 32.630 ;
        RECT 2274.340 32.310 2274.600 32.630 ;
        RECT 2274.400 2.000 2274.540 32.310 ;
        RECT 2274.190 -4.000 2274.750 2.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1636.750 1087.900 1637.070 1087.960 ;
        RECT 1641.810 1087.900 1642.130 1087.960 ;
        RECT 1636.750 1087.760 1642.130 1087.900 ;
        RECT 1636.750 1087.700 1637.070 1087.760 ;
        RECT 1641.810 1087.700 1642.130 1087.760 ;
        RECT 1641.810 32.200 1642.130 32.260 ;
        RECT 2292.250 32.200 2292.570 32.260 ;
        RECT 1641.810 32.060 2292.570 32.200 ;
        RECT 1641.810 32.000 1642.130 32.060 ;
        RECT 2292.250 32.000 2292.570 32.060 ;
      LAYER via ;
        RECT 1636.780 1087.700 1637.040 1087.960 ;
        RECT 1641.840 1087.700 1642.100 1087.960 ;
        RECT 1641.840 32.000 1642.100 32.260 ;
        RECT 2292.280 32.000 2292.540 32.260 ;
      LAYER met2 ;
        RECT 1636.690 1100.580 1636.970 1104.000 ;
        RECT 1636.690 1100.000 1636.980 1100.580 ;
        RECT 1636.840 1087.990 1636.980 1100.000 ;
        RECT 1636.780 1087.670 1637.040 1087.990 ;
        RECT 1641.840 1087.670 1642.100 1087.990 ;
        RECT 1641.900 32.290 1642.040 1087.670 ;
        RECT 1641.840 31.970 1642.100 32.290 ;
        RECT 2292.280 31.970 2292.540 32.290 ;
        RECT 2292.340 2.000 2292.480 31.970 ;
        RECT 2292.130 -4.000 2292.690 2.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1642.730 1087.900 1643.050 1087.960 ;
        RECT 1648.250 1087.900 1648.570 1087.960 ;
        RECT 1642.730 1087.760 1648.570 1087.900 ;
        RECT 1642.730 1087.700 1643.050 1087.760 ;
        RECT 1648.250 1087.700 1648.570 1087.760 ;
        RECT 1648.250 31.860 1648.570 31.920 ;
        RECT 2310.190 31.860 2310.510 31.920 ;
        RECT 1648.250 31.720 2310.510 31.860 ;
        RECT 1648.250 31.660 1648.570 31.720 ;
        RECT 2310.190 31.660 2310.510 31.720 ;
      LAYER via ;
        RECT 1642.760 1087.700 1643.020 1087.960 ;
        RECT 1648.280 1087.700 1648.540 1087.960 ;
        RECT 1648.280 31.660 1648.540 31.920 ;
        RECT 2310.220 31.660 2310.480 31.920 ;
      LAYER met2 ;
        RECT 1642.670 1100.580 1642.950 1104.000 ;
        RECT 1642.670 1100.000 1642.960 1100.580 ;
        RECT 1642.820 1087.990 1642.960 1100.000 ;
        RECT 1642.760 1087.670 1643.020 1087.990 ;
        RECT 1648.280 1087.670 1648.540 1087.990 ;
        RECT 1648.340 31.950 1648.480 1087.670 ;
        RECT 1648.280 31.630 1648.540 31.950 ;
        RECT 2310.220 31.630 2310.480 31.950 ;
        RECT 2310.280 2.000 2310.420 31.630 ;
        RECT 2310.070 -4.000 2310.630 2.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1648.710 31.520 1649.030 31.580 ;
        RECT 2328.130 31.520 2328.450 31.580 ;
        RECT 1648.710 31.380 2328.450 31.520 ;
        RECT 1648.710 31.320 1649.030 31.380 ;
        RECT 2328.130 31.320 2328.450 31.380 ;
      LAYER via ;
        RECT 1648.740 31.320 1649.000 31.580 ;
        RECT 2328.160 31.320 2328.420 31.580 ;
      LAYER met2 ;
        RECT 1648.650 1100.580 1648.930 1104.000 ;
        RECT 1648.650 1100.000 1648.940 1100.580 ;
        RECT 1648.800 31.610 1648.940 1100.000 ;
        RECT 1648.740 31.290 1649.000 31.610 ;
        RECT 2328.160 31.290 2328.420 31.610 ;
        RECT 2328.220 2.000 2328.360 31.290 ;
        RECT 2328.010 -4.000 2328.570 2.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1655.610 31.180 1655.930 31.240 ;
        RECT 2345.610 31.180 2345.930 31.240 ;
        RECT 1655.610 31.040 2345.930 31.180 ;
        RECT 1655.610 30.980 1655.930 31.040 ;
        RECT 2345.610 30.980 2345.930 31.040 ;
      LAYER via ;
        RECT 1655.640 30.980 1655.900 31.240 ;
        RECT 2345.640 30.980 2345.900 31.240 ;
      LAYER met2 ;
        RECT 1655.090 1100.650 1655.370 1104.000 ;
        RECT 1655.090 1100.510 1655.840 1100.650 ;
        RECT 1655.090 1100.000 1655.370 1100.510 ;
        RECT 1655.700 31.270 1655.840 1100.510 ;
        RECT 1655.640 30.950 1655.900 31.270 ;
        RECT 2345.640 30.950 2345.900 31.270 ;
        RECT 2345.700 2.000 2345.840 30.950 ;
        RECT 2345.490 -4.000 2346.050 2.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1662.510 30.840 1662.830 30.900 ;
        RECT 2363.550 30.840 2363.870 30.900 ;
        RECT 1662.510 30.700 2363.870 30.840 ;
        RECT 1662.510 30.640 1662.830 30.700 ;
        RECT 2363.550 30.640 2363.870 30.700 ;
      LAYER via ;
        RECT 1662.540 30.640 1662.800 30.900 ;
        RECT 2363.580 30.640 2363.840 30.900 ;
      LAYER met2 ;
        RECT 1661.070 1100.650 1661.350 1104.000 ;
        RECT 1661.070 1100.510 1662.740 1100.650 ;
        RECT 1661.070 1100.000 1661.350 1100.510 ;
        RECT 1662.600 30.930 1662.740 1100.510 ;
        RECT 1662.540 30.610 1662.800 30.930 ;
        RECT 2363.580 30.610 2363.840 30.930 ;
        RECT 2363.640 2.000 2363.780 30.610 ;
        RECT 2363.430 -4.000 2363.990 2.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1667.110 1088.580 1667.430 1088.640 ;
        RECT 1668.950 1088.580 1669.270 1088.640 ;
        RECT 1667.110 1088.440 1669.270 1088.580 ;
        RECT 1667.110 1088.380 1667.430 1088.440 ;
        RECT 1668.950 1088.380 1669.270 1088.440 ;
      LAYER via ;
        RECT 1667.140 1088.380 1667.400 1088.640 ;
        RECT 1668.980 1088.380 1669.240 1088.640 ;
      LAYER met2 ;
        RECT 1667.050 1100.580 1667.330 1104.000 ;
        RECT 1667.050 1100.000 1667.340 1100.580 ;
        RECT 1667.200 1088.670 1667.340 1100.000 ;
        RECT 1667.140 1088.350 1667.400 1088.670 ;
        RECT 1668.980 1088.350 1669.240 1088.670 ;
        RECT 1669.040 31.125 1669.180 1088.350 ;
        RECT 1668.970 30.755 1669.250 31.125 ;
        RECT 2381.510 30.755 2381.790 31.125 ;
        RECT 2381.580 2.000 2381.720 30.755 ;
        RECT 2381.370 -4.000 2381.930 2.000 ;
      LAYER via2 ;
        RECT 1668.970 30.800 1669.250 31.080 ;
        RECT 2381.510 30.800 2381.790 31.080 ;
      LAYER met3 ;
        RECT 1668.945 31.090 1669.275 31.105 ;
        RECT 2381.485 31.090 2381.815 31.105 ;
        RECT 1668.945 30.790 2381.815 31.090 ;
        RECT 1668.945 30.775 1669.275 30.790 ;
        RECT 2381.485 30.775 2381.815 30.790 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1673.550 1088.580 1673.870 1088.640 ;
        RECT 1676.310 1088.580 1676.630 1088.640 ;
        RECT 1673.550 1088.440 1676.630 1088.580 ;
        RECT 1673.550 1088.380 1673.870 1088.440 ;
        RECT 1676.310 1088.380 1676.630 1088.440 ;
        RECT 1676.310 61.440 1676.630 61.500 ;
        RECT 2394.370 61.440 2394.690 61.500 ;
        RECT 1676.310 61.300 2394.690 61.440 ;
        RECT 1676.310 61.240 1676.630 61.300 ;
        RECT 2394.370 61.240 2394.690 61.300 ;
        RECT 2394.370 2.620 2394.690 2.680 ;
        RECT 2399.430 2.620 2399.750 2.680 ;
        RECT 2394.370 2.480 2399.750 2.620 ;
        RECT 2394.370 2.420 2394.690 2.480 ;
        RECT 2399.430 2.420 2399.750 2.480 ;
      LAYER via ;
        RECT 1673.580 1088.380 1673.840 1088.640 ;
        RECT 1676.340 1088.380 1676.600 1088.640 ;
        RECT 1676.340 61.240 1676.600 61.500 ;
        RECT 2394.400 61.240 2394.660 61.500 ;
        RECT 2394.400 2.420 2394.660 2.680 ;
        RECT 2399.460 2.420 2399.720 2.680 ;
      LAYER met2 ;
        RECT 1673.490 1100.580 1673.770 1104.000 ;
        RECT 1673.490 1100.000 1673.780 1100.580 ;
        RECT 1673.640 1088.670 1673.780 1100.000 ;
        RECT 1673.580 1088.350 1673.840 1088.670 ;
        RECT 1676.340 1088.350 1676.600 1088.670 ;
        RECT 1676.400 61.530 1676.540 1088.350 ;
        RECT 1676.340 61.210 1676.600 61.530 ;
        RECT 2394.400 61.210 2394.660 61.530 ;
        RECT 2394.460 2.710 2394.600 61.210 ;
        RECT 2394.400 2.390 2394.660 2.710 ;
        RECT 2399.460 2.390 2399.720 2.710 ;
        RECT 2399.520 2.000 2399.660 2.390 ;
        RECT 2399.310 -4.000 2399.870 2.000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1117.870 1042.680 1118.190 1042.740 ;
        RECT 1120.630 1042.680 1120.950 1042.740 ;
        RECT 1117.870 1042.540 1120.950 1042.680 ;
        RECT 1117.870 1042.480 1118.190 1042.540 ;
        RECT 1120.630 1042.480 1120.950 1042.540 ;
        RECT 793.570 21.660 793.890 21.720 ;
        RECT 1117.870 21.660 1118.190 21.720 ;
        RECT 793.570 21.520 1118.190 21.660 ;
        RECT 793.570 21.460 793.890 21.520 ;
        RECT 1117.870 21.460 1118.190 21.520 ;
      LAYER via ;
        RECT 1117.900 1042.480 1118.160 1042.740 ;
        RECT 1120.660 1042.480 1120.920 1042.740 ;
        RECT 793.600 21.460 793.860 21.720 ;
        RECT 1117.900 21.460 1118.160 21.720 ;
      LAYER met2 ;
        RECT 1122.410 1100.650 1122.690 1104.000 ;
        RECT 1120.720 1100.510 1122.690 1100.650 ;
        RECT 1120.720 1042.770 1120.860 1100.510 ;
        RECT 1122.410 1100.000 1122.690 1100.510 ;
        RECT 1117.900 1042.450 1118.160 1042.770 ;
        RECT 1120.660 1042.450 1120.920 1042.770 ;
        RECT 1117.960 21.750 1118.100 1042.450 ;
        RECT 793.600 21.430 793.860 21.750 ;
        RECT 1117.900 21.430 1118.160 21.750 ;
        RECT 793.660 2.000 793.800 21.430 ;
        RECT 793.450 -4.000 794.010 2.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1064.050 1072.940 1064.370 1073.000 ;
        RECT 1067.730 1072.940 1068.050 1073.000 ;
        RECT 1064.050 1072.800 1068.050 1072.940 ;
        RECT 1064.050 1072.740 1064.370 1072.800 ;
        RECT 1067.730 1072.740 1068.050 1072.800 ;
        RECT 639.010 23.360 639.330 23.420 ;
        RECT 1064.050 23.360 1064.370 23.420 ;
        RECT 639.010 23.220 1064.370 23.360 ;
        RECT 639.010 23.160 639.330 23.220 ;
        RECT 1064.050 23.160 1064.370 23.220 ;
      LAYER via ;
        RECT 1064.080 1072.740 1064.340 1073.000 ;
        RECT 1067.760 1072.740 1068.020 1073.000 ;
        RECT 639.040 23.160 639.300 23.420 ;
        RECT 1064.080 23.160 1064.340 23.420 ;
      LAYER met2 ;
        RECT 1069.050 1100.650 1069.330 1104.000 ;
        RECT 1067.820 1100.510 1069.330 1100.650 ;
        RECT 1067.820 1073.030 1067.960 1100.510 ;
        RECT 1069.050 1100.000 1069.330 1100.510 ;
        RECT 1064.080 1072.710 1064.340 1073.030 ;
        RECT 1067.760 1072.710 1068.020 1073.030 ;
        RECT 1064.140 23.450 1064.280 1072.710 ;
        RECT 639.040 23.130 639.300 23.450 ;
        RECT 1064.080 23.130 1064.340 23.450 ;
        RECT 639.100 2.000 639.240 23.130 ;
        RECT 638.890 -4.000 639.450 2.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1682.290 61.100 1682.610 61.160 ;
        RECT 2421.970 61.100 2422.290 61.160 ;
        RECT 1682.290 60.960 2422.290 61.100 ;
        RECT 1682.290 60.900 1682.610 60.960 ;
        RECT 2421.970 60.900 2422.290 60.960 ;
      LAYER via ;
        RECT 1682.320 60.900 1682.580 61.160 ;
        RECT 2422.000 60.900 2422.260 61.160 ;
      LAYER met2 ;
        RECT 1681.310 1100.650 1681.590 1104.000 ;
        RECT 1681.310 1100.510 1682.520 1100.650 ;
        RECT 1681.310 1100.000 1681.590 1100.510 ;
        RECT 1682.380 61.190 1682.520 1100.510 ;
        RECT 1682.320 60.870 1682.580 61.190 ;
        RECT 2422.000 60.870 2422.260 61.190 ;
        RECT 2422.060 2.450 2422.200 60.870 ;
        RECT 2422.060 2.310 2423.120 2.450 ;
        RECT 2422.980 2.000 2423.120 2.310 ;
        RECT 2422.770 -4.000 2423.330 2.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1687.810 1088.580 1688.130 1088.640 ;
        RECT 1689.650 1088.580 1689.970 1088.640 ;
        RECT 1687.810 1088.440 1689.970 1088.580 ;
        RECT 1687.810 1088.380 1688.130 1088.440 ;
        RECT 1689.650 1088.380 1689.970 1088.440 ;
        RECT 1689.650 60.760 1689.970 60.820 ;
        RECT 2435.770 60.760 2436.090 60.820 ;
        RECT 1689.650 60.620 2436.090 60.760 ;
        RECT 1689.650 60.560 1689.970 60.620 ;
        RECT 2435.770 60.560 2436.090 60.620 ;
        RECT 2435.770 2.620 2436.090 2.680 ;
        RECT 2440.830 2.620 2441.150 2.680 ;
        RECT 2435.770 2.480 2441.150 2.620 ;
        RECT 2435.770 2.420 2436.090 2.480 ;
        RECT 2440.830 2.420 2441.150 2.480 ;
      LAYER via ;
        RECT 1687.840 1088.380 1688.100 1088.640 ;
        RECT 1689.680 1088.380 1689.940 1088.640 ;
        RECT 1689.680 60.560 1689.940 60.820 ;
        RECT 2435.800 60.560 2436.060 60.820 ;
        RECT 2435.800 2.420 2436.060 2.680 ;
        RECT 2440.860 2.420 2441.120 2.680 ;
      LAYER met2 ;
        RECT 1687.750 1100.580 1688.030 1104.000 ;
        RECT 1687.750 1100.000 1688.040 1100.580 ;
        RECT 1687.900 1088.670 1688.040 1100.000 ;
        RECT 1687.840 1088.350 1688.100 1088.670 ;
        RECT 1689.680 1088.350 1689.940 1088.670 ;
        RECT 1689.740 60.850 1689.880 1088.350 ;
        RECT 1689.680 60.530 1689.940 60.850 ;
        RECT 2435.800 60.530 2436.060 60.850 ;
        RECT 2435.860 2.710 2436.000 60.530 ;
        RECT 2435.800 2.390 2436.060 2.710 ;
        RECT 2440.860 2.390 2441.120 2.710 ;
        RECT 2440.920 2.000 2441.060 2.390 ;
        RECT 2440.710 -4.000 2441.270 2.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1693.790 1086.880 1694.110 1086.940 ;
        RECT 1696.550 1086.880 1696.870 1086.940 ;
        RECT 1693.790 1086.740 1696.870 1086.880 ;
        RECT 1693.790 1086.680 1694.110 1086.740 ;
        RECT 1696.550 1086.680 1696.870 1086.740 ;
        RECT 1696.550 60.420 1696.870 60.480 ;
        RECT 2456.470 60.420 2456.790 60.480 ;
        RECT 1696.550 60.280 2456.790 60.420 ;
        RECT 1696.550 60.220 1696.870 60.280 ;
        RECT 2456.470 60.220 2456.790 60.280 ;
      LAYER via ;
        RECT 1693.820 1086.680 1694.080 1086.940 ;
        RECT 1696.580 1086.680 1696.840 1086.940 ;
        RECT 1696.580 60.220 1696.840 60.480 ;
        RECT 2456.500 60.220 2456.760 60.480 ;
      LAYER met2 ;
        RECT 1693.730 1100.580 1694.010 1104.000 ;
        RECT 1693.730 1100.000 1694.020 1100.580 ;
        RECT 1693.880 1086.970 1694.020 1100.000 ;
        RECT 1693.820 1086.650 1694.080 1086.970 ;
        RECT 1696.580 1086.650 1696.840 1086.970 ;
        RECT 1696.640 60.510 1696.780 1086.650 ;
        RECT 1696.580 60.190 1696.840 60.510 ;
        RECT 2456.500 60.190 2456.760 60.510 ;
        RECT 2456.560 2.450 2456.700 60.190 ;
        RECT 2456.560 2.310 2459.000 2.450 ;
        RECT 2458.860 2.000 2459.000 2.310 ;
        RECT 2458.650 -4.000 2459.210 2.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1699.770 1087.220 1700.090 1087.280 ;
        RECT 1702.990 1087.220 1703.310 1087.280 ;
        RECT 1699.770 1087.080 1703.310 1087.220 ;
        RECT 1699.770 1087.020 1700.090 1087.080 ;
        RECT 1702.990 1087.020 1703.310 1087.080 ;
        RECT 1702.990 60.080 1703.310 60.140 ;
        RECT 2470.270 60.080 2470.590 60.140 ;
        RECT 1702.990 59.940 2470.590 60.080 ;
        RECT 1702.990 59.880 1703.310 59.940 ;
        RECT 2470.270 59.880 2470.590 59.940 ;
        RECT 2470.270 16.900 2470.590 16.960 ;
        RECT 2476.710 16.900 2477.030 16.960 ;
        RECT 2470.270 16.760 2477.030 16.900 ;
        RECT 2470.270 16.700 2470.590 16.760 ;
        RECT 2476.710 16.700 2477.030 16.760 ;
      LAYER via ;
        RECT 1699.800 1087.020 1700.060 1087.280 ;
        RECT 1703.020 1087.020 1703.280 1087.280 ;
        RECT 1703.020 59.880 1703.280 60.140 ;
        RECT 2470.300 59.880 2470.560 60.140 ;
        RECT 2470.300 16.700 2470.560 16.960 ;
        RECT 2476.740 16.700 2477.000 16.960 ;
      LAYER met2 ;
        RECT 1699.710 1100.580 1699.990 1104.000 ;
        RECT 1699.710 1100.000 1700.000 1100.580 ;
        RECT 1699.860 1087.310 1700.000 1100.000 ;
        RECT 1699.800 1086.990 1700.060 1087.310 ;
        RECT 1703.020 1086.990 1703.280 1087.310 ;
        RECT 1703.080 60.170 1703.220 1086.990 ;
        RECT 1703.020 59.850 1703.280 60.170 ;
        RECT 2470.300 59.850 2470.560 60.170 ;
        RECT 2470.360 16.990 2470.500 59.850 ;
        RECT 2470.300 16.670 2470.560 16.990 ;
        RECT 2476.740 16.670 2477.000 16.990 ;
        RECT 2476.800 2.000 2476.940 16.670 ;
        RECT 2476.590 -4.000 2477.150 2.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1705.750 1088.580 1706.070 1088.640 ;
        RECT 1710.350 1088.580 1710.670 1088.640 ;
        RECT 1705.750 1088.440 1710.670 1088.580 ;
        RECT 1705.750 1088.380 1706.070 1088.440 ;
        RECT 1710.350 1088.380 1710.670 1088.440 ;
        RECT 1710.350 59.740 1710.670 59.800 ;
        RECT 2490.970 59.740 2491.290 59.800 ;
        RECT 1710.350 59.600 2491.290 59.740 ;
        RECT 1710.350 59.540 1710.670 59.600 ;
        RECT 2490.970 59.540 2491.290 59.600 ;
      LAYER via ;
        RECT 1705.780 1088.380 1706.040 1088.640 ;
        RECT 1710.380 1088.380 1710.640 1088.640 ;
        RECT 1710.380 59.540 1710.640 59.800 ;
        RECT 2491.000 59.540 2491.260 59.800 ;
      LAYER met2 ;
        RECT 1705.690 1100.580 1705.970 1104.000 ;
        RECT 1705.690 1100.000 1705.980 1100.580 ;
        RECT 1705.840 1088.670 1705.980 1100.000 ;
        RECT 1705.780 1088.350 1706.040 1088.670 ;
        RECT 1710.380 1088.350 1710.640 1088.670 ;
        RECT 1710.440 59.830 1710.580 1088.350 ;
        RECT 1710.380 59.510 1710.640 59.830 ;
        RECT 2491.000 59.510 2491.260 59.830 ;
        RECT 2491.060 2.450 2491.200 59.510 ;
        RECT 2491.060 2.310 2494.880 2.450 ;
        RECT 2494.740 2.000 2494.880 2.310 ;
        RECT 2494.530 -4.000 2495.090 2.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1712.190 1088.580 1712.510 1088.640 ;
        RECT 1717.250 1088.580 1717.570 1088.640 ;
        RECT 1712.190 1088.440 1717.570 1088.580 ;
        RECT 1712.190 1088.380 1712.510 1088.440 ;
        RECT 1717.250 1088.380 1717.570 1088.440 ;
        RECT 1717.250 59.400 1717.570 59.460 ;
        RECT 2512.130 59.400 2512.450 59.460 ;
        RECT 1717.250 59.260 2512.450 59.400 ;
        RECT 1717.250 59.200 1717.570 59.260 ;
        RECT 2512.130 59.200 2512.450 59.260 ;
      LAYER via ;
        RECT 1712.220 1088.380 1712.480 1088.640 ;
        RECT 1717.280 1088.380 1717.540 1088.640 ;
        RECT 1717.280 59.200 1717.540 59.460 ;
        RECT 2512.160 59.200 2512.420 59.460 ;
      LAYER met2 ;
        RECT 1712.130 1100.580 1712.410 1104.000 ;
        RECT 1712.130 1100.000 1712.420 1100.580 ;
        RECT 1712.280 1088.670 1712.420 1100.000 ;
        RECT 1712.220 1088.350 1712.480 1088.670 ;
        RECT 1717.280 1088.350 1717.540 1088.670 ;
        RECT 1717.340 59.490 1717.480 1088.350 ;
        RECT 1717.280 59.170 1717.540 59.490 ;
        RECT 2512.160 59.170 2512.420 59.490 ;
        RECT 2512.220 2.000 2512.360 59.170 ;
        RECT 2512.010 -4.000 2512.570 2.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1718.170 1083.820 1718.490 1083.880 ;
        RECT 1723.690 1083.820 1724.010 1083.880 ;
        RECT 1718.170 1083.680 1724.010 1083.820 ;
        RECT 1718.170 1083.620 1718.490 1083.680 ;
        RECT 1723.690 1083.620 1724.010 1083.680 ;
        RECT 1723.690 59.060 1724.010 59.120 ;
        RECT 2525.470 59.060 2525.790 59.120 ;
        RECT 1723.690 58.920 2525.790 59.060 ;
        RECT 1723.690 58.860 1724.010 58.920 ;
        RECT 2525.470 58.860 2525.790 58.920 ;
      LAYER via ;
        RECT 1718.200 1083.620 1718.460 1083.880 ;
        RECT 1723.720 1083.620 1723.980 1083.880 ;
        RECT 1723.720 58.860 1723.980 59.120 ;
        RECT 2525.500 58.860 2525.760 59.120 ;
      LAYER met2 ;
        RECT 1718.110 1100.580 1718.390 1104.000 ;
        RECT 1718.110 1100.000 1718.400 1100.580 ;
        RECT 1718.260 1083.910 1718.400 1100.000 ;
        RECT 1718.200 1083.590 1718.460 1083.910 ;
        RECT 1723.720 1083.590 1723.980 1083.910 ;
        RECT 1723.780 59.150 1723.920 1083.590 ;
        RECT 1723.720 58.830 1723.980 59.150 ;
        RECT 2525.500 58.830 2525.760 59.150 ;
        RECT 2525.560 16.730 2525.700 58.830 ;
        RECT 2525.560 16.590 2530.300 16.730 ;
        RECT 2530.160 2.000 2530.300 16.590 ;
        RECT 2529.950 -4.000 2530.510 2.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1724.610 34.920 1724.930 34.980 ;
        RECT 2548.010 34.920 2548.330 34.980 ;
        RECT 1724.610 34.780 2548.330 34.920 ;
        RECT 1724.610 34.720 1724.930 34.780 ;
        RECT 2548.010 34.720 2548.330 34.780 ;
      LAYER via ;
        RECT 1724.640 34.720 1724.900 34.980 ;
        RECT 2548.040 34.720 2548.300 34.980 ;
      LAYER met2 ;
        RECT 1724.090 1100.650 1724.370 1104.000 ;
        RECT 1724.090 1100.510 1724.840 1100.650 ;
        RECT 1724.090 1100.000 1724.370 1100.510 ;
        RECT 1724.700 35.010 1724.840 1100.510 ;
        RECT 1724.640 34.690 1724.900 35.010 ;
        RECT 2548.040 34.690 2548.300 35.010 ;
        RECT 2548.100 2.000 2548.240 34.690 ;
        RECT 2547.890 -4.000 2548.450 2.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1731.050 35.260 1731.370 35.320 ;
        RECT 2565.950 35.260 2566.270 35.320 ;
        RECT 1731.050 35.120 2566.270 35.260 ;
        RECT 1731.050 35.060 1731.370 35.120 ;
        RECT 2565.950 35.060 2566.270 35.120 ;
      LAYER via ;
        RECT 1731.080 35.060 1731.340 35.320 ;
        RECT 2565.980 35.060 2566.240 35.320 ;
      LAYER met2 ;
        RECT 1730.530 1100.650 1730.810 1104.000 ;
        RECT 1730.530 1100.510 1731.280 1100.650 ;
        RECT 1730.530 1100.000 1730.810 1100.510 ;
        RECT 1731.140 35.350 1731.280 1100.510 ;
        RECT 1731.080 35.030 1731.340 35.350 ;
        RECT 2565.980 35.030 2566.240 35.350 ;
        RECT 2566.040 2.000 2566.180 35.030 ;
        RECT 2565.830 -4.000 2566.390 2.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1737.950 35.600 1738.270 35.660 ;
        RECT 2583.890 35.600 2584.210 35.660 ;
        RECT 1737.950 35.460 2584.210 35.600 ;
        RECT 1737.950 35.400 1738.270 35.460 ;
        RECT 2583.890 35.400 2584.210 35.460 ;
      LAYER via ;
        RECT 1737.980 35.400 1738.240 35.660 ;
        RECT 2583.920 35.400 2584.180 35.660 ;
      LAYER met2 ;
        RECT 1736.510 1100.650 1736.790 1104.000 ;
        RECT 1736.510 1100.510 1738.180 1100.650 ;
        RECT 1736.510 1100.000 1736.790 1100.510 ;
        RECT 1738.040 35.690 1738.180 1100.510 ;
        RECT 1737.980 35.370 1738.240 35.690 ;
        RECT 2583.920 35.370 2584.180 35.690 ;
        RECT 2583.980 2.000 2584.120 35.370 ;
        RECT 2583.770 -4.000 2584.330 2.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1124.770 1052.200 1125.090 1052.260 ;
        RECT 1128.910 1052.200 1129.230 1052.260 ;
        RECT 1124.770 1052.060 1129.230 1052.200 ;
        RECT 1124.770 1052.000 1125.090 1052.060 ;
        RECT 1128.910 1052.000 1129.230 1052.060 ;
        RECT 817.490 21.320 817.810 21.380 ;
        RECT 1124.770 21.320 1125.090 21.380 ;
        RECT 817.490 21.180 1125.090 21.320 ;
        RECT 817.490 21.120 817.810 21.180 ;
        RECT 1124.770 21.120 1125.090 21.180 ;
      LAYER via ;
        RECT 1124.800 1052.000 1125.060 1052.260 ;
        RECT 1128.940 1052.000 1129.200 1052.260 ;
        RECT 817.520 21.120 817.780 21.380 ;
        RECT 1124.800 21.120 1125.060 21.380 ;
      LAYER met2 ;
        RECT 1130.230 1100.650 1130.510 1104.000 ;
        RECT 1129.000 1100.510 1130.510 1100.650 ;
        RECT 1129.000 1052.290 1129.140 1100.510 ;
        RECT 1130.230 1100.000 1130.510 1100.510 ;
        RECT 1124.800 1051.970 1125.060 1052.290 ;
        RECT 1128.940 1051.970 1129.200 1052.290 ;
        RECT 1124.860 21.410 1125.000 1051.970 ;
        RECT 817.520 21.090 817.780 21.410 ;
        RECT 1124.800 21.090 1125.060 21.410 ;
        RECT 817.580 2.000 817.720 21.090 ;
        RECT 817.370 -4.000 817.930 2.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1742.550 1088.580 1742.870 1088.640 ;
        RECT 1744.850 1088.580 1745.170 1088.640 ;
        RECT 1742.550 1088.440 1745.170 1088.580 ;
        RECT 1742.550 1088.380 1742.870 1088.440 ;
        RECT 1744.850 1088.380 1745.170 1088.440 ;
        RECT 1743.930 35.940 1744.250 36.000 ;
        RECT 2601.830 35.940 2602.150 36.000 ;
        RECT 1743.930 35.800 2602.150 35.940 ;
        RECT 1743.930 35.740 1744.250 35.800 ;
        RECT 2601.830 35.740 2602.150 35.800 ;
      LAYER via ;
        RECT 1742.580 1088.380 1742.840 1088.640 ;
        RECT 1744.880 1088.380 1745.140 1088.640 ;
        RECT 1743.960 35.740 1744.220 36.000 ;
        RECT 2601.860 35.740 2602.120 36.000 ;
      LAYER met2 ;
        RECT 1742.490 1100.580 1742.770 1104.000 ;
        RECT 1742.490 1100.000 1742.780 1100.580 ;
        RECT 1742.640 1088.670 1742.780 1100.000 ;
        RECT 1742.580 1088.350 1742.840 1088.670 ;
        RECT 1744.880 1088.350 1745.140 1088.670 ;
        RECT 1744.940 49.370 1745.080 1088.350 ;
        RECT 1744.020 49.230 1745.080 49.370 ;
        RECT 1744.020 36.030 1744.160 49.230 ;
        RECT 1743.960 35.710 1744.220 36.030 ;
        RECT 2601.860 35.710 2602.120 36.030 ;
        RECT 2601.920 17.410 2602.060 35.710 ;
        RECT 2601.460 17.270 2602.060 17.410 ;
        RECT 2601.460 2.000 2601.600 17.270 ;
        RECT 2601.250 -4.000 2601.810 2.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1748.990 1088.580 1749.310 1088.640 ;
        RECT 1751.750 1088.580 1752.070 1088.640 ;
        RECT 1748.990 1088.440 1752.070 1088.580 ;
        RECT 1748.990 1088.380 1749.310 1088.440 ;
        RECT 1751.750 1088.380 1752.070 1088.440 ;
        RECT 1751.750 36.280 1752.070 36.340 ;
        RECT 2619.310 36.280 2619.630 36.340 ;
        RECT 1751.750 36.140 2619.630 36.280 ;
        RECT 1751.750 36.080 1752.070 36.140 ;
        RECT 2619.310 36.080 2619.630 36.140 ;
      LAYER via ;
        RECT 1749.020 1088.380 1749.280 1088.640 ;
        RECT 1751.780 1088.380 1752.040 1088.640 ;
        RECT 1751.780 36.080 1752.040 36.340 ;
        RECT 2619.340 36.080 2619.600 36.340 ;
      LAYER met2 ;
        RECT 1748.930 1100.580 1749.210 1104.000 ;
        RECT 1748.930 1100.000 1749.220 1100.580 ;
        RECT 1749.080 1088.670 1749.220 1100.000 ;
        RECT 1749.020 1088.350 1749.280 1088.670 ;
        RECT 1751.780 1088.350 1752.040 1088.670 ;
        RECT 1751.840 36.370 1751.980 1088.350 ;
        RECT 1751.780 36.050 1752.040 36.370 ;
        RECT 2619.340 36.050 2619.600 36.370 ;
        RECT 2619.400 2.000 2619.540 36.050 ;
        RECT 2619.190 -4.000 2619.750 2.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1754.970 1088.580 1755.290 1088.640 ;
        RECT 1758.190 1088.580 1758.510 1088.640 ;
        RECT 1754.970 1088.440 1758.510 1088.580 ;
        RECT 1754.970 1088.380 1755.290 1088.440 ;
        RECT 1758.190 1088.380 1758.510 1088.440 ;
        RECT 1758.190 36.620 1758.510 36.680 ;
        RECT 2637.250 36.620 2637.570 36.680 ;
        RECT 1758.190 36.480 2637.570 36.620 ;
        RECT 1758.190 36.420 1758.510 36.480 ;
        RECT 2637.250 36.420 2637.570 36.480 ;
      LAYER via ;
        RECT 1755.000 1088.380 1755.260 1088.640 ;
        RECT 1758.220 1088.380 1758.480 1088.640 ;
        RECT 1758.220 36.420 1758.480 36.680 ;
        RECT 2637.280 36.420 2637.540 36.680 ;
      LAYER met2 ;
        RECT 1754.910 1100.580 1755.190 1104.000 ;
        RECT 1754.910 1100.000 1755.200 1100.580 ;
        RECT 1755.060 1088.670 1755.200 1100.000 ;
        RECT 1755.000 1088.350 1755.260 1088.670 ;
        RECT 1758.220 1088.350 1758.480 1088.670 ;
        RECT 1758.280 36.710 1758.420 1088.350 ;
        RECT 1758.220 36.390 1758.480 36.710 ;
        RECT 2637.280 36.390 2637.540 36.710 ;
        RECT 2637.340 2.000 2637.480 36.390 ;
        RECT 2637.130 -4.000 2637.690 2.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1760.950 1088.580 1761.270 1088.640 ;
        RECT 1765.550 1088.580 1765.870 1088.640 ;
        RECT 1760.950 1088.440 1765.870 1088.580 ;
        RECT 1760.950 1088.380 1761.270 1088.440 ;
        RECT 1765.550 1088.380 1765.870 1088.440 ;
        RECT 1765.550 36.960 1765.870 37.020 ;
        RECT 2655.190 36.960 2655.510 37.020 ;
        RECT 1765.550 36.820 2655.510 36.960 ;
        RECT 1765.550 36.760 1765.870 36.820 ;
        RECT 2655.190 36.760 2655.510 36.820 ;
      LAYER via ;
        RECT 1760.980 1088.380 1761.240 1088.640 ;
        RECT 1765.580 1088.380 1765.840 1088.640 ;
        RECT 1765.580 36.760 1765.840 37.020 ;
        RECT 2655.220 36.760 2655.480 37.020 ;
      LAYER met2 ;
        RECT 1760.890 1100.580 1761.170 1104.000 ;
        RECT 1760.890 1100.000 1761.180 1100.580 ;
        RECT 1761.040 1088.670 1761.180 1100.000 ;
        RECT 1760.980 1088.350 1761.240 1088.670 ;
        RECT 1765.580 1088.350 1765.840 1088.670 ;
        RECT 1765.640 37.050 1765.780 1088.350 ;
        RECT 1765.580 36.730 1765.840 37.050 ;
        RECT 2655.220 36.730 2655.480 37.050 ;
        RECT 2655.280 2.000 2655.420 36.730 ;
        RECT 2655.070 -4.000 2655.630 2.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1767.390 1088.580 1767.710 1088.640 ;
        RECT 1772.450 1088.580 1772.770 1088.640 ;
        RECT 1767.390 1088.440 1772.770 1088.580 ;
        RECT 1767.390 1088.380 1767.710 1088.440 ;
        RECT 1772.450 1088.380 1772.770 1088.440 ;
        RECT 1772.450 37.300 1772.770 37.360 ;
        RECT 2672.670 37.300 2672.990 37.360 ;
        RECT 1772.450 37.160 2672.990 37.300 ;
        RECT 1772.450 37.100 1772.770 37.160 ;
        RECT 2672.670 37.100 2672.990 37.160 ;
      LAYER via ;
        RECT 1767.420 1088.380 1767.680 1088.640 ;
        RECT 1772.480 1088.380 1772.740 1088.640 ;
        RECT 1772.480 37.100 1772.740 37.360 ;
        RECT 2672.700 37.100 2672.960 37.360 ;
      LAYER met2 ;
        RECT 1767.330 1100.580 1767.610 1104.000 ;
        RECT 1767.330 1100.000 1767.620 1100.580 ;
        RECT 1767.480 1088.670 1767.620 1100.000 ;
        RECT 1767.420 1088.350 1767.680 1088.670 ;
        RECT 1772.480 1088.350 1772.740 1088.670 ;
        RECT 1772.540 37.390 1772.680 1088.350 ;
        RECT 1772.480 37.070 1772.740 37.390 ;
        RECT 2672.700 37.070 2672.960 37.390 ;
        RECT 2672.760 2.000 2672.900 37.070 ;
        RECT 2672.550 -4.000 2673.110 2.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1773.370 1088.920 1773.690 1088.980 ;
        RECT 1779.350 1088.920 1779.670 1088.980 ;
        RECT 1773.370 1088.780 1779.670 1088.920 ;
        RECT 1773.370 1088.720 1773.690 1088.780 ;
        RECT 1779.350 1088.720 1779.670 1088.780 ;
        RECT 1779.350 378.800 1779.670 379.060 ;
        RECT 1779.440 378.380 1779.580 378.800 ;
        RECT 1779.350 378.120 1779.670 378.380 ;
        RECT 1779.350 37.640 1779.670 37.700 ;
        RECT 2690.610 37.640 2690.930 37.700 ;
        RECT 1779.350 37.500 2690.930 37.640 ;
        RECT 1779.350 37.440 1779.670 37.500 ;
        RECT 2690.610 37.440 2690.930 37.500 ;
      LAYER via ;
        RECT 1773.400 1088.720 1773.660 1088.980 ;
        RECT 1779.380 1088.720 1779.640 1088.980 ;
        RECT 1779.380 378.800 1779.640 379.060 ;
        RECT 1779.380 378.120 1779.640 378.380 ;
        RECT 1779.380 37.440 1779.640 37.700 ;
        RECT 2690.640 37.440 2690.900 37.700 ;
      LAYER met2 ;
        RECT 1773.310 1100.580 1773.590 1104.000 ;
        RECT 1773.310 1100.000 1773.600 1100.580 ;
        RECT 1773.460 1089.010 1773.600 1100.000 ;
        RECT 1773.400 1088.690 1773.660 1089.010 ;
        RECT 1779.380 1088.690 1779.640 1089.010 ;
        RECT 1779.440 379.090 1779.580 1088.690 ;
        RECT 1779.380 378.770 1779.640 379.090 ;
        RECT 1779.380 378.090 1779.640 378.410 ;
        RECT 1779.440 37.730 1779.580 378.090 ;
        RECT 1779.380 37.410 1779.640 37.730 ;
        RECT 2690.640 37.410 2690.900 37.730 ;
        RECT 2690.700 2.000 2690.840 37.410 ;
        RECT 2690.490 -4.000 2691.050 2.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1778.890 627.680 1779.210 627.940 ;
        RECT 1778.980 627.260 1779.120 627.680 ;
        RECT 1778.890 627.000 1779.210 627.260 ;
        RECT 1778.890 378.460 1779.210 378.720 ;
        RECT 1778.980 378.040 1779.120 378.460 ;
        RECT 1778.890 377.780 1779.210 378.040 ;
        RECT 1778.890 41.380 1779.210 41.440 ;
        RECT 2708.550 41.380 2708.870 41.440 ;
        RECT 1778.890 41.240 2708.870 41.380 ;
        RECT 1778.890 41.180 1779.210 41.240 ;
        RECT 2708.550 41.180 2708.870 41.240 ;
      LAYER via ;
        RECT 1778.920 627.680 1779.180 627.940 ;
        RECT 1778.920 627.000 1779.180 627.260 ;
        RECT 1778.920 378.460 1779.180 378.720 ;
        RECT 1778.920 377.780 1779.180 378.040 ;
        RECT 1778.920 41.180 1779.180 41.440 ;
        RECT 2708.580 41.180 2708.840 41.440 ;
      LAYER met2 ;
        RECT 1779.290 1100.650 1779.570 1104.000 ;
        RECT 1778.980 1100.510 1779.570 1100.650 ;
        RECT 1778.980 627.970 1779.120 1100.510 ;
        RECT 1779.290 1100.000 1779.570 1100.510 ;
        RECT 1778.920 627.650 1779.180 627.970 ;
        RECT 1778.920 626.970 1779.180 627.290 ;
        RECT 1778.980 378.750 1779.120 626.970 ;
        RECT 1778.920 378.430 1779.180 378.750 ;
        RECT 1778.920 377.750 1779.180 378.070 ;
        RECT 1778.980 41.470 1779.120 377.750 ;
        RECT 1778.920 41.150 1779.180 41.470 ;
        RECT 2708.580 41.150 2708.840 41.470 ;
        RECT 2708.640 2.000 2708.780 41.150 ;
        RECT 2708.430 -4.000 2708.990 2.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1786.250 41.040 1786.570 41.100 ;
        RECT 2726.490 41.040 2726.810 41.100 ;
        RECT 1786.250 40.900 2726.810 41.040 ;
        RECT 1786.250 40.840 1786.570 40.900 ;
        RECT 2726.490 40.840 2726.810 40.900 ;
      LAYER via ;
        RECT 1786.280 40.840 1786.540 41.100 ;
        RECT 2726.520 40.840 2726.780 41.100 ;
      LAYER met2 ;
        RECT 1785.730 1100.650 1786.010 1104.000 ;
        RECT 1785.730 1100.510 1786.480 1100.650 ;
        RECT 1785.730 1100.000 1786.010 1100.510 ;
        RECT 1786.340 41.130 1786.480 1100.510 ;
        RECT 1786.280 40.810 1786.540 41.130 ;
        RECT 2726.520 40.810 2726.780 41.130 ;
        RECT 2726.580 2.000 2726.720 40.810 ;
        RECT 2726.370 -4.000 2726.930 2.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1793.150 40.700 1793.470 40.760 ;
        RECT 2744.430 40.700 2744.750 40.760 ;
        RECT 1793.150 40.560 2744.750 40.700 ;
        RECT 1793.150 40.500 1793.470 40.560 ;
        RECT 2744.430 40.500 2744.750 40.560 ;
      LAYER via ;
        RECT 1793.180 40.500 1793.440 40.760 ;
        RECT 2744.460 40.500 2744.720 40.760 ;
      LAYER met2 ;
        RECT 1791.710 1100.650 1791.990 1104.000 ;
        RECT 1791.710 1100.510 1793.380 1100.650 ;
        RECT 1791.710 1100.000 1791.990 1100.510 ;
        RECT 1793.240 40.790 1793.380 1100.510 ;
        RECT 1793.180 40.470 1793.440 40.790 ;
        RECT 2744.460 40.470 2744.720 40.790 ;
        RECT 2744.520 2.000 2744.660 40.470 ;
        RECT 2744.310 -4.000 2744.870 2.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1799.590 40.360 1799.910 40.420 ;
        RECT 2761.910 40.360 2762.230 40.420 ;
        RECT 1799.590 40.220 2762.230 40.360 ;
        RECT 1799.590 40.160 1799.910 40.220 ;
        RECT 2761.910 40.160 2762.230 40.220 ;
      LAYER via ;
        RECT 1799.620 40.160 1799.880 40.420 ;
        RECT 2761.940 40.160 2762.200 40.420 ;
      LAYER met2 ;
        RECT 1797.690 1100.650 1797.970 1104.000 ;
        RECT 1797.690 1100.510 1799.820 1100.650 ;
        RECT 1797.690 1100.000 1797.970 1100.510 ;
        RECT 1799.680 40.450 1799.820 1100.510 ;
        RECT 1799.620 40.130 1799.880 40.450 ;
        RECT 2761.940 40.130 2762.200 40.450 ;
        RECT 2762.000 2.000 2762.140 40.130 ;
        RECT 2761.790 -4.000 2762.350 2.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1131.670 1052.200 1131.990 1052.260 ;
        RECT 1135.350 1052.200 1135.670 1052.260 ;
        RECT 1131.670 1052.060 1135.670 1052.200 ;
        RECT 1131.670 1052.000 1131.990 1052.060 ;
        RECT 1135.350 1052.000 1135.670 1052.060 ;
        RECT 835.430 20.980 835.750 21.040 ;
        RECT 1131.670 20.980 1131.990 21.040 ;
        RECT 835.430 20.840 1131.990 20.980 ;
        RECT 835.430 20.780 835.750 20.840 ;
        RECT 1131.670 20.780 1131.990 20.840 ;
      LAYER via ;
        RECT 1131.700 1052.000 1131.960 1052.260 ;
        RECT 1135.380 1052.000 1135.640 1052.260 ;
        RECT 835.460 20.780 835.720 21.040 ;
        RECT 1131.700 20.780 1131.960 21.040 ;
      LAYER met2 ;
        RECT 1136.670 1100.650 1136.950 1104.000 ;
        RECT 1135.440 1100.510 1136.950 1100.650 ;
        RECT 1135.440 1052.290 1135.580 1100.510 ;
        RECT 1136.670 1100.000 1136.950 1100.510 ;
        RECT 1131.700 1051.970 1131.960 1052.290 ;
        RECT 1135.380 1051.970 1135.640 1052.290 ;
        RECT 1131.760 21.070 1131.900 1051.970 ;
        RECT 835.460 20.750 835.720 21.070 ;
        RECT 1131.700 20.750 1131.960 21.070 ;
        RECT 835.520 2.000 835.660 20.750 ;
        RECT 835.310 -4.000 835.870 2.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1806.105 752.505 1806.275 800.275 ;
        RECT 1807.025 662.405 1807.195 710.515 ;
        RECT 1806.105 427.465 1806.275 469.115 ;
        RECT 1806.565 396.525 1806.735 420.835 ;
        RECT 1806.565 144.925 1806.735 159.035 ;
        RECT 1806.105 89.845 1806.275 137.955 ;
      LAYER mcon ;
        RECT 1806.105 800.105 1806.275 800.275 ;
        RECT 1807.025 710.345 1807.195 710.515 ;
        RECT 1806.105 468.945 1806.275 469.115 ;
        RECT 1806.565 420.665 1806.735 420.835 ;
        RECT 1806.565 158.865 1806.735 159.035 ;
        RECT 1806.105 137.785 1806.275 137.955 ;
      LAYER met1 ;
        RECT 1803.730 1062.740 1804.050 1062.800 ;
        RECT 1806.490 1062.740 1806.810 1062.800 ;
        RECT 1803.730 1062.600 1806.810 1062.740 ;
        RECT 1803.730 1062.540 1804.050 1062.600 ;
        RECT 1806.490 1062.540 1806.810 1062.600 ;
        RECT 1804.650 910.760 1804.970 910.820 ;
        RECT 1806.030 910.760 1806.350 910.820 ;
        RECT 1804.650 910.620 1806.350 910.760 ;
        RECT 1804.650 910.560 1804.970 910.620 ;
        RECT 1806.030 910.560 1806.350 910.620 ;
        RECT 1805.570 862.480 1805.890 862.540 ;
        RECT 1806.950 862.480 1807.270 862.540 ;
        RECT 1805.570 862.340 1807.270 862.480 ;
        RECT 1805.570 862.280 1805.890 862.340 ;
        RECT 1806.950 862.280 1807.270 862.340 ;
        RECT 1806.030 800.260 1806.350 800.320 ;
        RECT 1805.835 800.120 1806.350 800.260 ;
        RECT 1806.030 800.060 1806.350 800.120 ;
        RECT 1806.045 752.660 1806.335 752.705 ;
        RECT 1806.045 752.520 1806.720 752.660 ;
        RECT 1806.045 752.475 1806.335 752.520 ;
        RECT 1806.580 752.380 1806.720 752.520 ;
        RECT 1806.490 752.120 1806.810 752.380 ;
        RECT 1806.950 710.500 1807.270 710.560 ;
        RECT 1806.755 710.360 1807.270 710.500 ;
        RECT 1806.950 710.300 1807.270 710.360 ;
        RECT 1806.950 662.560 1807.270 662.620 ;
        RECT 1806.755 662.420 1807.270 662.560 ;
        RECT 1806.950 662.360 1807.270 662.420 ;
        RECT 1806.490 621.080 1806.810 621.140 ;
        RECT 1806.950 621.080 1807.270 621.140 ;
        RECT 1806.490 620.940 1807.270 621.080 ;
        RECT 1806.490 620.880 1806.810 620.940 ;
        RECT 1806.950 620.880 1807.270 620.940 ;
        RECT 1806.030 579.940 1806.350 580.000 ;
        RECT 1806.490 579.940 1806.810 580.000 ;
        RECT 1806.030 579.800 1806.810 579.940 ;
        RECT 1806.030 579.740 1806.350 579.800 ;
        RECT 1806.490 579.740 1806.810 579.800 ;
        RECT 1806.030 469.100 1806.350 469.160 ;
        RECT 1805.835 468.960 1806.350 469.100 ;
        RECT 1806.030 468.900 1806.350 468.960 ;
        RECT 1806.030 427.620 1806.350 427.680 ;
        RECT 1805.835 427.480 1806.350 427.620 ;
        RECT 1806.030 427.420 1806.350 427.480 ;
        RECT 1806.490 420.820 1806.810 420.880 ;
        RECT 1806.295 420.680 1806.810 420.820 ;
        RECT 1806.490 420.620 1806.810 420.680 ;
        RECT 1806.505 396.680 1806.795 396.725 ;
        RECT 1806.950 396.680 1807.270 396.740 ;
        RECT 1806.505 396.540 1807.270 396.680 ;
        RECT 1806.505 396.495 1806.795 396.540 ;
        RECT 1806.950 396.480 1807.270 396.540 ;
        RECT 1806.505 159.020 1806.795 159.065 ;
        RECT 1806.950 159.020 1807.270 159.080 ;
        RECT 1806.505 158.880 1807.270 159.020 ;
        RECT 1806.505 158.835 1806.795 158.880 ;
        RECT 1806.950 158.820 1807.270 158.880 ;
        RECT 1806.490 145.080 1806.810 145.140 ;
        RECT 1806.295 144.940 1806.810 145.080 ;
        RECT 1806.490 144.880 1806.810 144.940 ;
        RECT 1806.045 137.940 1806.335 137.985 ;
        RECT 1806.490 137.940 1806.810 138.000 ;
        RECT 1806.045 137.800 1806.810 137.940 ;
        RECT 1806.045 137.755 1806.335 137.800 ;
        RECT 1806.490 137.740 1806.810 137.800 ;
        RECT 1806.030 90.000 1806.350 90.060 ;
        RECT 1805.835 89.860 1806.350 90.000 ;
        RECT 1806.030 89.800 1806.350 89.860 ;
        RECT 1806.490 40.020 1806.810 40.080 ;
        RECT 2779.850 40.020 2780.170 40.080 ;
        RECT 1806.490 39.880 2780.170 40.020 ;
        RECT 1806.490 39.820 1806.810 39.880 ;
        RECT 2779.850 39.820 2780.170 39.880 ;
      LAYER via ;
        RECT 1803.760 1062.540 1804.020 1062.800 ;
        RECT 1806.520 1062.540 1806.780 1062.800 ;
        RECT 1804.680 910.560 1804.940 910.820 ;
        RECT 1806.060 910.560 1806.320 910.820 ;
        RECT 1805.600 862.280 1805.860 862.540 ;
        RECT 1806.980 862.280 1807.240 862.540 ;
        RECT 1806.060 800.060 1806.320 800.320 ;
        RECT 1806.520 752.120 1806.780 752.380 ;
        RECT 1806.980 710.300 1807.240 710.560 ;
        RECT 1806.980 662.360 1807.240 662.620 ;
        RECT 1806.520 620.880 1806.780 621.140 ;
        RECT 1806.980 620.880 1807.240 621.140 ;
        RECT 1806.060 579.740 1806.320 580.000 ;
        RECT 1806.520 579.740 1806.780 580.000 ;
        RECT 1806.060 468.900 1806.320 469.160 ;
        RECT 1806.060 427.420 1806.320 427.680 ;
        RECT 1806.520 420.620 1806.780 420.880 ;
        RECT 1806.980 396.480 1807.240 396.740 ;
        RECT 1806.980 158.820 1807.240 159.080 ;
        RECT 1806.520 144.880 1806.780 145.140 ;
        RECT 1806.520 137.740 1806.780 138.000 ;
        RECT 1806.060 89.800 1806.320 90.060 ;
        RECT 1806.520 39.820 1806.780 40.080 ;
        RECT 2779.880 39.820 2780.140 40.080 ;
      LAYER met2 ;
        RECT 1803.670 1100.580 1803.950 1104.000 ;
        RECT 1803.670 1100.000 1803.960 1100.580 ;
        RECT 1803.820 1062.830 1803.960 1100.000 ;
        RECT 1803.760 1062.510 1804.020 1062.830 ;
        RECT 1806.520 1062.510 1806.780 1062.830 ;
        RECT 1806.580 980.290 1806.720 1062.510 ;
        RECT 1806.120 980.150 1806.720 980.290 ;
        RECT 1806.120 930.650 1806.260 980.150 ;
        RECT 1806.120 930.510 1806.720 930.650 ;
        RECT 1806.580 917.730 1806.720 930.510 ;
        RECT 1806.120 917.590 1806.720 917.730 ;
        RECT 1806.120 910.850 1806.260 917.590 ;
        RECT 1804.680 910.530 1804.940 910.850 ;
        RECT 1806.060 910.530 1806.320 910.850 ;
        RECT 1804.740 862.765 1804.880 910.530 ;
        RECT 1804.670 862.395 1804.950 862.765 ;
        RECT 1805.590 862.395 1805.870 862.765 ;
        RECT 1805.600 862.250 1805.860 862.395 ;
        RECT 1806.980 862.250 1807.240 862.570 ;
        RECT 1807.040 807.570 1807.180 862.250 ;
        RECT 1806.120 807.430 1807.180 807.570 ;
        RECT 1806.120 800.350 1806.260 807.430 ;
        RECT 1806.060 800.030 1806.320 800.350 ;
        RECT 1806.520 752.090 1806.780 752.410 ;
        RECT 1806.580 717.130 1806.720 752.090 ;
        RECT 1806.580 716.990 1807.180 717.130 ;
        RECT 1807.040 710.590 1807.180 716.990 ;
        RECT 1806.980 710.270 1807.240 710.590 ;
        RECT 1806.980 662.330 1807.240 662.650 ;
        RECT 1807.040 621.170 1807.180 662.330 ;
        RECT 1806.520 620.850 1806.780 621.170 ;
        RECT 1806.980 620.850 1807.240 621.170 ;
        RECT 1806.580 580.030 1806.720 620.850 ;
        RECT 1806.060 579.710 1806.320 580.030 ;
        RECT 1806.520 579.710 1806.780 580.030 ;
        RECT 1806.120 532.285 1806.260 579.710 ;
        RECT 1806.050 531.915 1806.330 532.285 ;
        RECT 1806.510 531.235 1806.790 531.605 ;
        RECT 1806.580 499.530 1806.720 531.235 ;
        RECT 1806.120 499.390 1806.720 499.530 ;
        RECT 1806.120 469.190 1806.260 499.390 ;
        RECT 1806.060 468.870 1806.320 469.190 ;
        RECT 1806.060 427.390 1806.320 427.710 ;
        RECT 1806.120 421.330 1806.260 427.390 ;
        RECT 1806.120 421.190 1806.720 421.330 ;
        RECT 1806.580 420.910 1806.720 421.190 ;
        RECT 1806.520 420.590 1806.780 420.910 ;
        RECT 1806.980 396.450 1807.240 396.770 ;
        RECT 1807.040 351.290 1807.180 396.450 ;
        RECT 1806.580 351.150 1807.180 351.290 ;
        RECT 1806.580 290.090 1806.720 351.150 ;
        RECT 1806.120 289.950 1806.720 290.090 ;
        RECT 1806.120 265.610 1806.260 289.950 ;
        RECT 1806.120 265.470 1807.180 265.610 ;
        RECT 1807.040 254.730 1807.180 265.470 ;
        RECT 1806.580 254.590 1807.180 254.730 ;
        RECT 1806.580 207.130 1806.720 254.590 ;
        RECT 1806.580 206.990 1807.180 207.130 ;
        RECT 1807.040 159.110 1807.180 206.990 ;
        RECT 1806.980 158.790 1807.240 159.110 ;
        RECT 1806.520 144.850 1806.780 145.170 ;
        RECT 1806.580 138.030 1806.720 144.850 ;
        RECT 1806.520 137.710 1806.780 138.030 ;
        RECT 1806.060 89.770 1806.320 90.090 ;
        RECT 1806.120 61.610 1806.260 89.770 ;
        RECT 1806.120 61.470 1806.720 61.610 ;
        RECT 1806.580 40.110 1806.720 61.470 ;
        RECT 1806.520 39.790 1806.780 40.110 ;
        RECT 2779.880 39.790 2780.140 40.110 ;
        RECT 2779.940 2.000 2780.080 39.790 ;
        RECT 2779.730 -4.000 2780.290 2.000 ;
      LAYER via2 ;
        RECT 1804.670 862.440 1804.950 862.720 ;
        RECT 1805.590 862.440 1805.870 862.720 ;
        RECT 1806.050 531.960 1806.330 532.240 ;
        RECT 1806.510 531.280 1806.790 531.560 ;
      LAYER met3 ;
        RECT 1804.645 862.730 1804.975 862.745 ;
        RECT 1805.565 862.730 1805.895 862.745 ;
        RECT 1804.645 862.430 1805.895 862.730 ;
        RECT 1804.645 862.415 1804.975 862.430 ;
        RECT 1805.565 862.415 1805.895 862.430 ;
        RECT 1806.025 532.250 1806.355 532.265 ;
        RECT 1806.025 531.950 1807.490 532.250 ;
        RECT 1806.025 531.935 1806.355 531.950 ;
        RECT 1806.485 531.570 1806.815 531.585 ;
        RECT 1807.190 531.570 1807.490 531.950 ;
        RECT 1806.485 531.270 1807.490 531.570 ;
        RECT 1806.485 531.255 1806.815 531.270 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1812.545 959.225 1812.715 1007.335 ;
        RECT 1812.085 855.865 1812.255 910.775 ;
        RECT 1812.085 807.245 1812.255 855.355 ;
        RECT 1812.085 724.285 1812.255 783.275 ;
        RECT 1811.625 579.445 1811.795 607.155 ;
        RECT 1811.625 338.045 1811.795 420.835 ;
        RECT 1811.625 241.485 1811.795 289.595 ;
        RECT 1812.085 144.925 1812.255 159.375 ;
        RECT 1812.545 48.365 1812.715 96.475 ;
      LAYER mcon ;
        RECT 1812.545 1007.165 1812.715 1007.335 ;
        RECT 1812.085 910.605 1812.255 910.775 ;
        RECT 1812.085 855.185 1812.255 855.355 ;
        RECT 1812.085 783.105 1812.255 783.275 ;
        RECT 1811.625 606.985 1811.795 607.155 ;
        RECT 1811.625 420.665 1811.795 420.835 ;
        RECT 1811.625 289.425 1811.795 289.595 ;
        RECT 1812.085 159.205 1812.255 159.375 ;
        RECT 1812.545 96.305 1812.715 96.475 ;
      LAYER met1 ;
        RECT 1810.170 1089.260 1810.490 1089.320 ;
        RECT 1812.930 1089.260 1813.250 1089.320 ;
        RECT 1810.170 1089.120 1813.250 1089.260 ;
        RECT 1810.170 1089.060 1810.490 1089.120 ;
        RECT 1812.930 1089.060 1813.250 1089.120 ;
        RECT 1812.485 1007.320 1812.775 1007.365 ;
        RECT 1812.930 1007.320 1813.250 1007.380 ;
        RECT 1812.485 1007.180 1813.250 1007.320 ;
        RECT 1812.485 1007.135 1812.775 1007.180 ;
        RECT 1812.930 1007.120 1813.250 1007.180 ;
        RECT 1812.470 959.380 1812.790 959.440 ;
        RECT 1812.275 959.240 1812.790 959.380 ;
        RECT 1812.470 959.180 1812.790 959.240 ;
        RECT 1812.025 910.760 1812.315 910.805 ;
        RECT 1812.930 910.760 1813.250 910.820 ;
        RECT 1812.025 910.620 1813.250 910.760 ;
        RECT 1812.025 910.575 1812.315 910.620 ;
        RECT 1812.930 910.560 1813.250 910.620 ;
        RECT 1811.550 856.020 1811.870 856.080 ;
        RECT 1812.025 856.020 1812.315 856.065 ;
        RECT 1811.550 855.880 1812.315 856.020 ;
        RECT 1811.550 855.820 1811.870 855.880 ;
        RECT 1812.025 855.835 1812.315 855.880 ;
        RECT 1812.010 855.340 1812.330 855.400 ;
        RECT 1811.815 855.200 1812.330 855.340 ;
        RECT 1812.010 855.140 1812.330 855.200 ;
        RECT 1812.010 807.400 1812.330 807.460 ;
        RECT 1811.815 807.260 1812.330 807.400 ;
        RECT 1812.010 807.200 1812.330 807.260 ;
        RECT 1812.010 783.260 1812.330 783.320 ;
        RECT 1811.815 783.120 1812.330 783.260 ;
        RECT 1812.010 783.060 1812.330 783.120 ;
        RECT 1812.010 724.440 1812.330 724.500 ;
        RECT 1811.815 724.300 1812.330 724.440 ;
        RECT 1812.010 724.240 1812.330 724.300 ;
        RECT 1811.550 638.420 1811.870 638.480 ;
        RECT 1812.930 638.420 1813.250 638.480 ;
        RECT 1811.550 638.280 1813.250 638.420 ;
        RECT 1811.550 638.220 1811.870 638.280 ;
        RECT 1812.930 638.220 1813.250 638.280 ;
        RECT 1811.550 607.140 1811.870 607.200 ;
        RECT 1811.355 607.000 1811.870 607.140 ;
        RECT 1811.550 606.940 1811.870 607.000 ;
        RECT 1811.550 579.600 1811.870 579.660 ;
        RECT 1811.355 579.460 1811.870 579.600 ;
        RECT 1811.550 579.400 1811.870 579.460 ;
        RECT 1811.550 427.960 1811.870 428.020 ;
        RECT 1812.470 427.960 1812.790 428.020 ;
        RECT 1811.550 427.820 1812.790 427.960 ;
        RECT 1811.550 427.760 1811.870 427.820 ;
        RECT 1812.470 427.760 1812.790 427.820 ;
        RECT 1811.565 420.820 1811.855 420.865 ;
        RECT 1812.470 420.820 1812.790 420.880 ;
        RECT 1811.565 420.680 1812.790 420.820 ;
        RECT 1811.565 420.635 1811.855 420.680 ;
        RECT 1812.470 420.620 1812.790 420.680 ;
        RECT 1811.550 338.200 1811.870 338.260 ;
        RECT 1811.355 338.060 1811.870 338.200 ;
        RECT 1811.550 338.000 1811.870 338.060 ;
        RECT 1811.090 337.520 1811.410 337.580 ;
        RECT 1811.550 337.520 1811.870 337.580 ;
        RECT 1811.090 337.380 1811.870 337.520 ;
        RECT 1811.090 337.320 1811.410 337.380 ;
        RECT 1811.550 337.320 1811.870 337.380 ;
        RECT 1811.550 289.580 1811.870 289.640 ;
        RECT 1811.355 289.440 1811.870 289.580 ;
        RECT 1811.550 289.380 1811.870 289.440 ;
        RECT 1811.565 241.640 1811.855 241.685 ;
        RECT 1812.470 241.640 1812.790 241.700 ;
        RECT 1811.565 241.500 1812.790 241.640 ;
        RECT 1811.565 241.455 1811.855 241.500 ;
        RECT 1812.470 241.440 1812.790 241.500 ;
        RECT 1812.025 159.360 1812.315 159.405 ;
        RECT 1812.930 159.360 1813.250 159.420 ;
        RECT 1812.025 159.220 1813.250 159.360 ;
        RECT 1812.025 159.175 1812.315 159.220 ;
        RECT 1812.930 159.160 1813.250 159.220 ;
        RECT 1812.010 145.080 1812.330 145.140 ;
        RECT 1811.815 144.940 1812.330 145.080 ;
        RECT 1812.010 144.880 1812.330 144.940 ;
        RECT 1812.485 96.460 1812.775 96.505 ;
        RECT 1812.930 96.460 1813.250 96.520 ;
        RECT 1812.485 96.320 1813.250 96.460 ;
        RECT 1812.485 96.275 1812.775 96.320 ;
        RECT 1812.930 96.260 1813.250 96.320 ;
        RECT 1812.470 48.520 1812.790 48.580 ;
        RECT 1812.275 48.380 1812.790 48.520 ;
        RECT 1812.470 48.320 1812.790 48.380 ;
        RECT 1817.990 39.680 1818.310 39.740 ;
        RECT 2797.790 39.680 2798.110 39.740 ;
        RECT 1817.990 39.540 2798.110 39.680 ;
        RECT 1817.990 39.480 1818.310 39.540 ;
        RECT 2797.790 39.480 2798.110 39.540 ;
      LAYER via ;
        RECT 1810.200 1089.060 1810.460 1089.320 ;
        RECT 1812.960 1089.060 1813.220 1089.320 ;
        RECT 1812.960 1007.120 1813.220 1007.380 ;
        RECT 1812.500 959.180 1812.760 959.440 ;
        RECT 1812.960 910.560 1813.220 910.820 ;
        RECT 1811.580 855.820 1811.840 856.080 ;
        RECT 1812.040 855.140 1812.300 855.400 ;
        RECT 1812.040 807.200 1812.300 807.460 ;
        RECT 1812.040 783.060 1812.300 783.320 ;
        RECT 1812.040 724.240 1812.300 724.500 ;
        RECT 1811.580 638.220 1811.840 638.480 ;
        RECT 1812.960 638.220 1813.220 638.480 ;
        RECT 1811.580 606.940 1811.840 607.200 ;
        RECT 1811.580 579.400 1811.840 579.660 ;
        RECT 1811.580 427.760 1811.840 428.020 ;
        RECT 1812.500 427.760 1812.760 428.020 ;
        RECT 1812.500 420.620 1812.760 420.880 ;
        RECT 1811.580 338.000 1811.840 338.260 ;
        RECT 1811.120 337.320 1811.380 337.580 ;
        RECT 1811.580 337.320 1811.840 337.580 ;
        RECT 1811.580 289.380 1811.840 289.640 ;
        RECT 1812.500 241.440 1812.760 241.700 ;
        RECT 1812.960 159.160 1813.220 159.420 ;
        RECT 1812.040 144.880 1812.300 145.140 ;
        RECT 1812.960 96.260 1813.220 96.520 ;
        RECT 1812.500 48.320 1812.760 48.580 ;
        RECT 1818.020 39.480 1818.280 39.740 ;
        RECT 2797.820 39.480 2798.080 39.740 ;
      LAYER met2 ;
        RECT 1810.110 1100.580 1810.390 1104.000 ;
        RECT 1810.110 1100.000 1810.400 1100.580 ;
        RECT 1810.260 1089.350 1810.400 1100.000 ;
        RECT 1810.200 1089.030 1810.460 1089.350 ;
        RECT 1812.960 1089.030 1813.220 1089.350 ;
        RECT 1813.020 1007.410 1813.160 1089.030 ;
        RECT 1812.960 1007.090 1813.220 1007.410 ;
        RECT 1812.500 959.150 1812.760 959.470 ;
        RECT 1812.560 917.730 1812.700 959.150 ;
        RECT 1812.560 917.590 1813.160 917.730 ;
        RECT 1813.020 910.850 1813.160 917.590 ;
        RECT 1812.960 910.530 1813.220 910.850 ;
        RECT 1811.580 855.850 1811.840 856.110 ;
        RECT 1811.580 855.790 1812.240 855.850 ;
        RECT 1811.640 855.710 1812.240 855.790 ;
        RECT 1812.100 855.430 1812.240 855.710 ;
        RECT 1812.040 855.110 1812.300 855.430 ;
        RECT 1812.040 807.170 1812.300 807.490 ;
        RECT 1812.100 783.350 1812.240 807.170 ;
        RECT 1812.040 783.030 1812.300 783.350 ;
        RECT 1812.040 724.210 1812.300 724.530 ;
        RECT 1812.100 717.810 1812.240 724.210 ;
        RECT 1812.100 717.670 1812.700 717.810 ;
        RECT 1812.560 689.250 1812.700 717.670 ;
        RECT 1811.640 689.110 1812.700 689.250 ;
        RECT 1811.640 638.510 1811.780 689.110 ;
        RECT 1811.580 638.190 1811.840 638.510 ;
        RECT 1812.960 638.190 1813.220 638.510 ;
        RECT 1813.020 614.565 1813.160 638.190 ;
        RECT 1811.570 614.195 1811.850 614.565 ;
        RECT 1812.950 614.195 1813.230 614.565 ;
        RECT 1811.640 607.230 1811.780 614.195 ;
        RECT 1811.580 606.910 1811.840 607.230 ;
        RECT 1811.580 579.370 1811.840 579.690 ;
        RECT 1811.640 428.050 1811.780 579.370 ;
        RECT 1811.580 427.730 1811.840 428.050 ;
        RECT 1812.500 427.730 1812.760 428.050 ;
        RECT 1812.560 420.910 1812.700 427.730 ;
        RECT 1812.500 420.590 1812.760 420.910 ;
        RECT 1811.580 337.970 1811.840 338.290 ;
        RECT 1811.640 337.610 1811.780 337.970 ;
        RECT 1811.120 337.290 1811.380 337.610 ;
        RECT 1811.580 337.290 1811.840 337.610 ;
        RECT 1811.180 335.650 1811.320 337.290 ;
        RECT 1811.180 335.510 1811.780 335.650 ;
        RECT 1811.640 289.670 1811.780 335.510 ;
        RECT 1811.580 289.350 1811.840 289.670 ;
        RECT 1812.500 241.410 1812.760 241.730 ;
        RECT 1812.560 207.130 1812.700 241.410 ;
        RECT 1812.560 206.990 1813.160 207.130 ;
        RECT 1813.020 159.450 1813.160 206.990 ;
        RECT 1812.960 159.130 1813.220 159.450 ;
        RECT 1812.040 144.850 1812.300 145.170 ;
        RECT 1812.100 110.570 1812.240 144.850 ;
        RECT 1812.100 110.430 1813.160 110.570 ;
        RECT 1813.020 96.550 1813.160 110.430 ;
        RECT 1812.960 96.230 1813.220 96.550 ;
        RECT 1812.500 48.290 1812.760 48.610 ;
        RECT 1812.560 48.125 1812.700 48.290 ;
        RECT 1812.490 47.755 1812.770 48.125 ;
        RECT 1818.010 47.075 1818.290 47.445 ;
        RECT 1818.080 39.770 1818.220 47.075 ;
        RECT 1818.020 39.450 1818.280 39.770 ;
        RECT 2797.820 39.450 2798.080 39.770 ;
        RECT 2797.880 2.000 2798.020 39.450 ;
        RECT 2797.670 -4.000 2798.230 2.000 ;
      LAYER via2 ;
        RECT 1811.570 614.240 1811.850 614.520 ;
        RECT 1812.950 614.240 1813.230 614.520 ;
        RECT 1812.490 47.800 1812.770 48.080 ;
        RECT 1818.010 47.120 1818.290 47.400 ;
      LAYER met3 ;
        RECT 1811.545 614.530 1811.875 614.545 ;
        RECT 1812.925 614.530 1813.255 614.545 ;
        RECT 1811.545 614.230 1813.255 614.530 ;
        RECT 1811.545 614.215 1811.875 614.230 ;
        RECT 1812.925 614.215 1813.255 614.230 ;
        RECT 1812.465 48.090 1812.795 48.105 ;
        RECT 1812.465 47.775 1813.010 48.090 ;
        RECT 1812.710 47.410 1813.010 47.775 ;
        RECT 1817.985 47.410 1818.315 47.425 ;
        RECT 1812.710 47.110 1818.315 47.410 ;
        RECT 1817.985 47.095 1818.315 47.110 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1816.150 1088.580 1816.470 1088.640 ;
        RECT 1820.750 1088.580 1821.070 1088.640 ;
        RECT 1816.150 1088.440 1821.070 1088.580 ;
        RECT 1816.150 1088.380 1816.470 1088.440 ;
        RECT 1820.750 1088.380 1821.070 1088.440 ;
        RECT 1820.750 39.340 1821.070 39.400 ;
        RECT 2815.730 39.340 2816.050 39.400 ;
        RECT 1820.750 39.200 2816.050 39.340 ;
        RECT 1820.750 39.140 1821.070 39.200 ;
        RECT 2815.730 39.140 2816.050 39.200 ;
      LAYER via ;
        RECT 1816.180 1088.380 1816.440 1088.640 ;
        RECT 1820.780 1088.380 1821.040 1088.640 ;
        RECT 1820.780 39.140 1821.040 39.400 ;
        RECT 2815.760 39.140 2816.020 39.400 ;
      LAYER met2 ;
        RECT 1816.090 1100.580 1816.370 1104.000 ;
        RECT 1816.090 1100.000 1816.380 1100.580 ;
        RECT 1816.240 1088.670 1816.380 1100.000 ;
        RECT 1816.180 1088.350 1816.440 1088.670 ;
        RECT 1820.780 1088.350 1821.040 1088.670 ;
        RECT 1820.840 39.430 1820.980 1088.350 ;
        RECT 1820.780 39.110 1821.040 39.430 ;
        RECT 2815.760 39.110 2816.020 39.430 ;
        RECT 2815.820 2.000 2815.960 39.110 ;
        RECT 2815.610 -4.000 2816.170 2.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1822.130 1088.580 1822.450 1088.640 ;
        RECT 1827.190 1088.580 1827.510 1088.640 ;
        RECT 1822.130 1088.440 1827.510 1088.580 ;
        RECT 1822.130 1088.380 1822.450 1088.440 ;
        RECT 1827.190 1088.380 1827.510 1088.440 ;
        RECT 1827.190 39.000 1827.510 39.060 ;
        RECT 2833.670 39.000 2833.990 39.060 ;
        RECT 1827.190 38.860 2833.990 39.000 ;
        RECT 1827.190 38.800 1827.510 38.860 ;
        RECT 2833.670 38.800 2833.990 38.860 ;
      LAYER via ;
        RECT 1822.160 1088.380 1822.420 1088.640 ;
        RECT 1827.220 1088.380 1827.480 1088.640 ;
        RECT 1827.220 38.800 1827.480 39.060 ;
        RECT 2833.700 38.800 2833.960 39.060 ;
      LAYER met2 ;
        RECT 1822.070 1100.580 1822.350 1104.000 ;
        RECT 1822.070 1100.000 1822.360 1100.580 ;
        RECT 1822.220 1088.670 1822.360 1100.000 ;
        RECT 1822.160 1088.350 1822.420 1088.670 ;
        RECT 1827.220 1088.350 1827.480 1088.670 ;
        RECT 1827.280 39.090 1827.420 1088.350 ;
        RECT 1827.220 38.770 1827.480 39.090 ;
        RECT 2833.700 38.770 2833.960 39.090 ;
        RECT 2833.760 2.000 2833.900 38.770 ;
        RECT 2833.550 -4.000 2834.110 2.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1828.570 1088.920 1828.890 1088.980 ;
        RECT 1834.090 1088.920 1834.410 1088.980 ;
        RECT 1828.570 1088.780 1834.410 1088.920 ;
        RECT 1828.570 1088.720 1828.890 1088.780 ;
        RECT 1834.090 1088.720 1834.410 1088.780 ;
        RECT 1834.090 38.660 1834.410 38.720 ;
        RECT 2851.150 38.660 2851.470 38.720 ;
        RECT 1834.090 38.520 2851.470 38.660 ;
        RECT 1834.090 38.460 1834.410 38.520 ;
        RECT 2851.150 38.460 2851.470 38.520 ;
      LAYER via ;
        RECT 1828.600 1088.720 1828.860 1088.980 ;
        RECT 1834.120 1088.720 1834.380 1088.980 ;
        RECT 1834.120 38.460 1834.380 38.720 ;
        RECT 2851.180 38.460 2851.440 38.720 ;
      LAYER met2 ;
        RECT 1828.510 1100.580 1828.790 1104.000 ;
        RECT 1828.510 1100.000 1828.800 1100.580 ;
        RECT 1828.660 1089.010 1828.800 1100.000 ;
        RECT 1828.600 1088.690 1828.860 1089.010 ;
        RECT 1834.120 1088.690 1834.380 1089.010 ;
        RECT 1834.180 38.750 1834.320 1088.690 ;
        RECT 1834.120 38.430 1834.380 38.750 ;
        RECT 2851.180 38.430 2851.440 38.750 ;
        RECT 2851.240 2.000 2851.380 38.430 ;
        RECT 2851.030 -4.000 2851.590 2.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1835.010 38.320 1835.330 38.380 ;
        RECT 2869.090 38.320 2869.410 38.380 ;
        RECT 1835.010 38.180 2869.410 38.320 ;
        RECT 1835.010 38.120 1835.330 38.180 ;
        RECT 2869.090 38.120 2869.410 38.180 ;
      LAYER via ;
        RECT 1835.040 38.120 1835.300 38.380 ;
        RECT 2869.120 38.120 2869.380 38.380 ;
      LAYER met2 ;
        RECT 1834.490 1100.580 1834.770 1104.000 ;
        RECT 1834.490 1100.000 1834.780 1100.580 ;
        RECT 1834.640 50.050 1834.780 1100.000 ;
        RECT 1834.640 49.910 1835.240 50.050 ;
        RECT 1835.100 38.410 1835.240 49.910 ;
        RECT 1835.040 38.090 1835.300 38.410 ;
        RECT 2869.120 38.090 2869.380 38.410 ;
        RECT 2869.180 2.000 2869.320 38.090 ;
        RECT 2868.970 -4.000 2869.530 2.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1840.990 37.980 1841.310 38.040 ;
        RECT 2887.030 37.980 2887.350 38.040 ;
        RECT 1840.990 37.840 2887.350 37.980 ;
        RECT 1840.990 37.780 1841.310 37.840 ;
        RECT 2887.030 37.780 2887.350 37.840 ;
      LAYER via ;
        RECT 1841.020 37.780 1841.280 38.040 ;
        RECT 2887.060 37.780 2887.320 38.040 ;
      LAYER met2 ;
        RECT 1840.470 1100.650 1840.750 1104.000 ;
        RECT 1840.470 1100.510 1841.220 1100.650 ;
        RECT 1840.470 1100.000 1840.750 1100.510 ;
        RECT 1841.080 38.070 1841.220 1100.510 ;
        RECT 1841.020 37.750 1841.280 38.070 ;
        RECT 2887.060 37.750 2887.320 38.070 ;
        RECT 2887.120 2.000 2887.260 37.750 ;
        RECT 2886.910 -4.000 2887.470 2.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1846.910 1100.650 1847.190 1104.000 ;
        RECT 1846.910 1100.510 1848.120 1100.650 ;
        RECT 1846.910 1100.000 1847.190 1100.510 ;
        RECT 1847.980 37.925 1848.120 1100.510 ;
        RECT 1847.910 37.555 1848.190 37.925 ;
        RECT 2904.990 37.555 2905.270 37.925 ;
        RECT 2905.060 2.000 2905.200 37.555 ;
        RECT 2904.850 -4.000 2905.410 2.000 ;
      LAYER via2 ;
        RECT 1847.910 37.600 1848.190 37.880 ;
        RECT 2904.990 37.600 2905.270 37.880 ;
      LAYER met3 ;
        RECT 1847.885 37.890 1848.215 37.905 ;
        RECT 2904.965 37.890 2905.295 37.905 ;
        RECT 1847.885 37.590 2905.295 37.890 ;
        RECT 1847.885 37.575 1848.215 37.590 ;
        RECT 2904.965 37.575 2905.295 37.590 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1140.945 697.085 1141.115 786.675 ;
        RECT 1140.945 234.345 1141.115 275.995 ;
      LAYER mcon ;
        RECT 1140.945 786.505 1141.115 786.675 ;
        RECT 1140.945 275.825 1141.115 275.995 ;
      LAYER met1 ;
        RECT 1141.330 910.760 1141.650 910.820 ;
        RECT 1141.790 910.760 1142.110 910.820 ;
        RECT 1141.330 910.620 1142.110 910.760 ;
        RECT 1141.330 910.560 1141.650 910.620 ;
        RECT 1141.790 910.560 1142.110 910.620 ;
        RECT 1141.790 793.460 1142.110 793.520 ;
        RECT 1142.710 793.460 1143.030 793.520 ;
        RECT 1141.790 793.320 1143.030 793.460 ;
        RECT 1141.790 793.260 1142.110 793.320 ;
        RECT 1142.710 793.260 1143.030 793.320 ;
        RECT 1140.885 786.660 1141.175 786.705 ;
        RECT 1142.710 786.660 1143.030 786.720 ;
        RECT 1140.885 786.520 1143.030 786.660 ;
        RECT 1140.885 786.475 1141.175 786.520 ;
        RECT 1142.710 786.460 1143.030 786.520 ;
        RECT 1140.870 697.240 1141.190 697.300 ;
        RECT 1140.675 697.100 1141.190 697.240 ;
        RECT 1140.870 697.040 1141.190 697.100 ;
        RECT 1141.330 669.020 1141.650 669.080 ;
        RECT 1142.250 669.020 1142.570 669.080 ;
        RECT 1141.330 668.880 1142.570 669.020 ;
        RECT 1141.330 668.820 1141.650 668.880 ;
        RECT 1142.250 668.820 1142.570 668.880 ;
        RECT 1140.870 434.760 1141.190 434.820 ;
        RECT 1141.330 434.760 1141.650 434.820 ;
        RECT 1140.870 434.620 1141.650 434.760 ;
        RECT 1140.870 434.560 1141.190 434.620 ;
        RECT 1141.330 434.560 1141.650 434.620 ;
        RECT 1140.870 427.620 1141.190 427.680 ;
        RECT 1141.330 427.620 1141.650 427.680 ;
        RECT 1140.870 427.480 1141.650 427.620 ;
        RECT 1140.870 427.420 1141.190 427.480 ;
        RECT 1141.330 427.420 1141.650 427.480 ;
        RECT 1140.870 275.980 1141.190 276.040 ;
        RECT 1140.675 275.840 1141.190 275.980 ;
        RECT 1140.870 275.780 1141.190 275.840 ;
        RECT 1140.885 234.500 1141.175 234.545 ;
        RECT 1141.330 234.500 1141.650 234.560 ;
        RECT 1140.885 234.360 1141.650 234.500 ;
        RECT 1140.885 234.315 1141.175 234.360 ;
        RECT 1141.330 234.300 1141.650 234.360 ;
        RECT 1140.870 227.700 1141.190 227.760 ;
        RECT 1141.330 227.700 1141.650 227.760 ;
        RECT 1140.870 227.560 1141.650 227.700 ;
        RECT 1140.870 227.500 1141.190 227.560 ;
        RECT 1141.330 227.500 1141.650 227.560 ;
        RECT 852.910 24.040 853.230 24.100 ;
        RECT 1140.870 24.040 1141.190 24.100 ;
        RECT 852.910 23.900 1141.190 24.040 ;
        RECT 852.910 23.840 853.230 23.900 ;
        RECT 1140.870 23.840 1141.190 23.900 ;
      LAYER via ;
        RECT 1141.360 910.560 1141.620 910.820 ;
        RECT 1141.820 910.560 1142.080 910.820 ;
        RECT 1141.820 793.260 1142.080 793.520 ;
        RECT 1142.740 793.260 1143.000 793.520 ;
        RECT 1142.740 786.460 1143.000 786.720 ;
        RECT 1140.900 697.040 1141.160 697.300 ;
        RECT 1141.360 668.820 1141.620 669.080 ;
        RECT 1142.280 668.820 1142.540 669.080 ;
        RECT 1140.900 434.560 1141.160 434.820 ;
        RECT 1141.360 434.560 1141.620 434.820 ;
        RECT 1140.900 427.420 1141.160 427.680 ;
        RECT 1141.360 427.420 1141.620 427.680 ;
        RECT 1140.900 275.780 1141.160 276.040 ;
        RECT 1141.360 234.300 1141.620 234.560 ;
        RECT 1140.900 227.500 1141.160 227.760 ;
        RECT 1141.360 227.500 1141.620 227.760 ;
        RECT 852.940 23.840 853.200 24.100 ;
        RECT 1140.900 23.840 1141.160 24.100 ;
      LAYER met2 ;
        RECT 1142.650 1101.330 1142.930 1104.000 ;
        RECT 1141.420 1101.190 1142.930 1101.330 ;
        RECT 1141.420 910.850 1141.560 1101.190 ;
        RECT 1142.650 1100.000 1142.930 1101.190 ;
        RECT 1141.360 910.530 1141.620 910.850 ;
        RECT 1141.820 910.530 1142.080 910.850 ;
        RECT 1141.880 793.550 1142.020 910.530 ;
        RECT 1141.820 793.230 1142.080 793.550 ;
        RECT 1142.740 793.230 1143.000 793.550 ;
        RECT 1142.800 786.750 1142.940 793.230 ;
        RECT 1142.740 786.430 1143.000 786.750 ;
        RECT 1140.900 697.010 1141.160 697.330 ;
        RECT 1140.960 696.730 1141.100 697.010 ;
        RECT 1141.350 696.730 1141.630 696.845 ;
        RECT 1140.960 696.590 1141.630 696.730 ;
        RECT 1141.350 696.475 1141.630 696.590 ;
        RECT 1142.270 696.475 1142.550 696.845 ;
        RECT 1142.340 669.110 1142.480 696.475 ;
        RECT 1141.360 668.790 1141.620 669.110 ;
        RECT 1142.280 668.790 1142.540 669.110 ;
        RECT 1141.420 613.770 1141.560 668.790 ;
        RECT 1141.420 613.630 1142.020 613.770 ;
        RECT 1141.880 554.610 1142.020 613.630 ;
        RECT 1141.420 554.470 1142.020 554.610 ;
        RECT 1141.420 498.170 1141.560 554.470 ;
        RECT 1141.420 498.030 1142.020 498.170 ;
        RECT 1141.880 496.810 1142.020 498.030 ;
        RECT 1141.420 496.670 1142.020 496.810 ;
        RECT 1141.420 434.850 1141.560 496.670 ;
        RECT 1140.900 434.530 1141.160 434.850 ;
        RECT 1141.360 434.530 1141.620 434.850 ;
        RECT 1140.960 427.710 1141.100 434.530 ;
        RECT 1140.900 427.390 1141.160 427.710 ;
        RECT 1141.360 427.390 1141.620 427.710 ;
        RECT 1141.420 379.850 1141.560 427.390 ;
        RECT 1140.960 379.710 1141.560 379.850 ;
        RECT 1140.960 276.070 1141.100 379.710 ;
        RECT 1140.900 275.750 1141.160 276.070 ;
        RECT 1141.360 234.270 1141.620 234.590 ;
        RECT 1141.420 227.790 1141.560 234.270 ;
        RECT 1140.900 227.470 1141.160 227.790 ;
        RECT 1141.360 227.470 1141.620 227.790 ;
        RECT 1140.960 89.490 1141.100 227.470 ;
        RECT 1140.960 89.350 1141.560 89.490 ;
        RECT 1141.420 42.570 1141.560 89.350 ;
        RECT 1140.960 42.430 1141.560 42.570 ;
        RECT 1140.960 24.130 1141.100 42.430 ;
        RECT 852.940 23.810 853.200 24.130 ;
        RECT 1140.900 23.810 1141.160 24.130 ;
        RECT 853.000 2.000 853.140 23.810 ;
        RECT 852.790 -4.000 853.350 2.000 ;
      LAYER via2 ;
        RECT 1141.350 696.520 1141.630 696.800 ;
        RECT 1142.270 696.520 1142.550 696.800 ;
      LAYER met3 ;
        RECT 1141.325 696.810 1141.655 696.825 ;
        RECT 1142.245 696.810 1142.575 696.825 ;
        RECT 1141.325 696.510 1142.575 696.810 ;
        RECT 1141.325 696.495 1141.655 696.510 ;
        RECT 1142.245 696.495 1142.575 696.510 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1145.470 1052.200 1145.790 1052.260 ;
        RECT 1147.310 1052.200 1147.630 1052.260 ;
        RECT 1145.470 1052.060 1147.630 1052.200 ;
        RECT 1145.470 1052.000 1145.790 1052.060 ;
        RECT 1147.310 1052.000 1147.630 1052.060 ;
        RECT 870.850 24.380 871.170 24.440 ;
        RECT 1145.470 24.380 1145.790 24.440 ;
        RECT 870.850 24.240 1145.790 24.380 ;
        RECT 870.850 24.180 871.170 24.240 ;
        RECT 1145.470 24.180 1145.790 24.240 ;
      LAYER via ;
        RECT 1145.500 1052.000 1145.760 1052.260 ;
        RECT 1147.340 1052.000 1147.600 1052.260 ;
        RECT 870.880 24.180 871.140 24.440 ;
        RECT 1145.500 24.180 1145.760 24.440 ;
      LAYER met2 ;
        RECT 1148.630 1100.650 1148.910 1104.000 ;
        RECT 1147.400 1100.510 1148.910 1100.650 ;
        RECT 1147.400 1052.290 1147.540 1100.510 ;
        RECT 1148.630 1100.000 1148.910 1100.510 ;
        RECT 1145.500 1051.970 1145.760 1052.290 ;
        RECT 1147.340 1051.970 1147.600 1052.290 ;
        RECT 1145.560 24.470 1145.700 1051.970 ;
        RECT 870.880 24.150 871.140 24.470 ;
        RECT 1145.500 24.150 1145.760 24.470 ;
        RECT 870.940 2.000 871.080 24.150 ;
        RECT 870.730 -4.000 871.290 2.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1153.290 1029.420 1153.610 1029.480 ;
        RECT 1154.210 1029.420 1154.530 1029.480 ;
        RECT 1153.290 1029.280 1154.530 1029.420 ;
        RECT 1153.290 1029.220 1153.610 1029.280 ;
        RECT 1154.210 1029.220 1154.530 1029.280 ;
        RECT 888.790 45.120 889.110 45.180 ;
        RECT 1153.290 45.120 1153.610 45.180 ;
        RECT 888.790 44.980 1153.610 45.120 ;
        RECT 888.790 44.920 889.110 44.980 ;
        RECT 1153.290 44.920 1153.610 44.980 ;
      LAYER via ;
        RECT 1153.320 1029.220 1153.580 1029.480 ;
        RECT 1154.240 1029.220 1154.500 1029.480 ;
        RECT 888.820 44.920 889.080 45.180 ;
        RECT 1153.320 44.920 1153.580 45.180 ;
      LAYER met2 ;
        RECT 1155.070 1100.650 1155.350 1104.000 ;
        RECT 1154.300 1100.510 1155.350 1100.650 ;
        RECT 1154.300 1029.510 1154.440 1100.510 ;
        RECT 1155.070 1100.000 1155.350 1100.510 ;
        RECT 1153.320 1029.190 1153.580 1029.510 ;
        RECT 1154.240 1029.190 1154.500 1029.510 ;
        RECT 1153.380 45.210 1153.520 1029.190 ;
        RECT 888.820 44.890 889.080 45.210 ;
        RECT 1153.320 44.890 1153.580 45.210 ;
        RECT 888.880 2.000 889.020 44.890 ;
        RECT 888.670 -4.000 889.230 2.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 906.730 17.240 907.050 17.300 ;
        RECT 906.730 17.100 1132.360 17.240 ;
        RECT 906.730 17.040 907.050 17.100 ;
        RECT 1132.220 16.900 1132.360 17.100 ;
        RECT 1159.730 16.900 1160.050 16.960 ;
        RECT 1132.220 16.760 1160.050 16.900 ;
        RECT 1159.730 16.700 1160.050 16.760 ;
      LAYER via ;
        RECT 906.760 17.040 907.020 17.300 ;
        RECT 1159.760 16.700 1160.020 16.960 ;
      LAYER met2 ;
        RECT 1161.050 1100.650 1161.330 1104.000 ;
        RECT 1159.820 1100.510 1161.330 1100.650 ;
        RECT 906.760 17.010 907.020 17.330 ;
        RECT 906.820 2.000 906.960 17.010 ;
        RECT 1159.820 16.990 1159.960 1100.510 ;
        RECT 1161.050 1100.000 1161.330 1100.510 ;
        RECT 1159.760 16.670 1160.020 16.990 ;
        RECT 906.610 -4.000 907.170 2.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1125.305 16.745 1125.475 17.595 ;
        RECT 1131.745 16.745 1131.915 19.635 ;
      LAYER mcon ;
        RECT 1131.745 19.465 1131.915 19.635 ;
        RECT 1125.305 17.425 1125.475 17.595 ;
      LAYER met1 ;
        RECT 1131.685 19.620 1131.975 19.665 ;
        RECT 1166.170 19.620 1166.490 19.680 ;
        RECT 1131.685 19.480 1166.490 19.620 ;
        RECT 1131.685 19.435 1131.975 19.480 ;
        RECT 1166.170 19.420 1166.490 19.480 ;
        RECT 924.210 17.580 924.530 17.640 ;
        RECT 1125.245 17.580 1125.535 17.625 ;
        RECT 924.210 17.440 1125.535 17.580 ;
        RECT 924.210 17.380 924.530 17.440 ;
        RECT 1125.245 17.395 1125.535 17.440 ;
        RECT 1125.245 16.900 1125.535 16.945 ;
        RECT 1131.685 16.900 1131.975 16.945 ;
        RECT 1125.245 16.760 1131.975 16.900 ;
        RECT 1125.245 16.715 1125.535 16.760 ;
        RECT 1131.685 16.715 1131.975 16.760 ;
      LAYER via ;
        RECT 1166.200 19.420 1166.460 19.680 ;
        RECT 924.240 17.380 924.500 17.640 ;
      LAYER met2 ;
        RECT 1167.030 1100.650 1167.310 1104.000 ;
        RECT 1166.260 1100.510 1167.310 1100.650 ;
        RECT 1166.260 19.710 1166.400 1100.510 ;
        RECT 1167.030 1100.000 1167.310 1100.510 ;
        RECT 1166.200 19.390 1166.460 19.710 ;
        RECT 924.240 17.350 924.500 17.670 ;
        RECT 924.300 2.000 924.440 17.350 ;
        RECT 924.090 -4.000 924.650 2.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1173.990 1028.540 1174.310 1028.800 ;
        RECT 1174.080 1028.120 1174.220 1028.540 ;
        RECT 1173.990 1027.860 1174.310 1028.120 ;
        RECT 1173.990 989.980 1174.310 990.040 ;
        RECT 1175.830 989.980 1176.150 990.040 ;
        RECT 1173.990 989.840 1176.150 989.980 ;
        RECT 1173.990 989.780 1174.310 989.840 ;
        RECT 1175.830 989.780 1176.150 989.840 ;
        RECT 1175.370 820.800 1175.690 821.060 ;
        RECT 1175.460 820.660 1175.600 820.800 ;
        RECT 1175.830 820.660 1176.150 820.720 ;
        RECT 1175.460 820.520 1176.150 820.660 ;
        RECT 1175.830 820.460 1176.150 820.520 ;
        RECT 1174.910 772.720 1175.230 772.780 ;
        RECT 1175.830 772.720 1176.150 772.780 ;
        RECT 1174.910 772.580 1176.150 772.720 ;
        RECT 1174.910 772.520 1175.230 772.580 ;
        RECT 1175.830 772.520 1176.150 772.580 ;
        RECT 1175.370 710.300 1175.690 710.560 ;
        RECT 1175.460 710.160 1175.600 710.300 ;
        RECT 1175.830 710.160 1176.150 710.220 ;
        RECT 1175.460 710.020 1176.150 710.160 ;
        RECT 1175.830 709.960 1176.150 710.020 ;
        RECT 1175.370 627.680 1175.690 627.940 ;
        RECT 1175.460 627.540 1175.600 627.680 ;
        RECT 1175.830 627.540 1176.150 627.600 ;
        RECT 1175.460 627.400 1176.150 627.540 ;
        RECT 1175.830 627.340 1176.150 627.400 ;
        RECT 1175.370 531.120 1175.690 531.380 ;
        RECT 1175.460 530.980 1175.600 531.120 ;
        RECT 1175.830 530.980 1176.150 531.040 ;
        RECT 1175.460 530.840 1176.150 530.980 ;
        RECT 1175.830 530.780 1176.150 530.840 ;
        RECT 1175.830 483.040 1176.150 483.100 ;
        RECT 1176.750 483.040 1177.070 483.100 ;
        RECT 1175.830 482.900 1177.070 483.040 ;
        RECT 1175.830 482.840 1176.150 482.900 ;
        RECT 1176.750 482.840 1177.070 482.900 ;
        RECT 1175.370 434.560 1175.690 434.820 ;
        RECT 1175.460 434.420 1175.600 434.560 ;
        RECT 1175.830 434.420 1176.150 434.480 ;
        RECT 1175.460 434.280 1176.150 434.420 ;
        RECT 1175.830 434.220 1176.150 434.280 ;
        RECT 1175.830 338.540 1176.150 338.600 ;
        RECT 1175.460 338.400 1176.150 338.540 ;
        RECT 1175.460 338.260 1175.600 338.400 ;
        RECT 1175.830 338.340 1176.150 338.400 ;
        RECT 1175.370 338.000 1175.690 338.260 ;
        RECT 1175.370 330.860 1175.690 331.120 ;
        RECT 1175.460 330.720 1175.600 330.860 ;
        RECT 1175.830 330.720 1176.150 330.780 ;
        RECT 1175.460 330.580 1176.150 330.720 ;
        RECT 1175.830 330.520 1176.150 330.580 ;
        RECT 1175.830 241.980 1176.150 242.040 ;
        RECT 1175.460 241.840 1176.150 241.980 ;
        RECT 1175.460 241.700 1175.600 241.840 ;
        RECT 1175.830 241.780 1176.150 241.840 ;
        RECT 1175.370 241.440 1175.690 241.700 ;
        RECT 1173.990 207.300 1174.310 207.360 ;
        RECT 1175.370 207.300 1175.690 207.360 ;
        RECT 1173.990 207.160 1175.690 207.300 ;
        RECT 1173.990 207.100 1174.310 207.160 ;
        RECT 1175.370 207.100 1175.690 207.160 ;
        RECT 1173.990 159.020 1174.310 159.080 ;
        RECT 1173.620 158.880 1174.310 159.020 ;
        RECT 1173.620 158.740 1173.760 158.880 ;
        RECT 1173.990 158.820 1174.310 158.880 ;
        RECT 1173.530 158.480 1173.850 158.740 ;
        RECT 1173.530 125.700 1173.850 125.760 ;
        RECT 1175.830 125.700 1176.150 125.760 ;
        RECT 1173.530 125.560 1176.150 125.700 ;
        RECT 1173.530 125.500 1173.850 125.560 ;
        RECT 1175.830 125.500 1176.150 125.560 ;
        RECT 1173.530 62.460 1173.850 62.520 ;
        RECT 1175.830 62.460 1176.150 62.520 ;
        RECT 1173.530 62.320 1176.150 62.460 ;
        RECT 1173.530 62.260 1173.850 62.320 ;
        RECT 1175.830 62.260 1176.150 62.320 ;
        RECT 942.150 18.260 942.470 18.320 ;
        RECT 1173.530 18.260 1173.850 18.320 ;
        RECT 942.150 18.120 1173.850 18.260 ;
        RECT 942.150 18.060 942.470 18.120 ;
        RECT 1173.530 18.060 1173.850 18.120 ;
      LAYER via ;
        RECT 1174.020 1028.540 1174.280 1028.800 ;
        RECT 1174.020 1027.860 1174.280 1028.120 ;
        RECT 1174.020 989.780 1174.280 990.040 ;
        RECT 1175.860 989.780 1176.120 990.040 ;
        RECT 1175.400 820.800 1175.660 821.060 ;
        RECT 1175.860 820.460 1176.120 820.720 ;
        RECT 1174.940 772.520 1175.200 772.780 ;
        RECT 1175.860 772.520 1176.120 772.780 ;
        RECT 1175.400 710.300 1175.660 710.560 ;
        RECT 1175.860 709.960 1176.120 710.220 ;
        RECT 1175.400 627.680 1175.660 627.940 ;
        RECT 1175.860 627.340 1176.120 627.600 ;
        RECT 1175.400 531.120 1175.660 531.380 ;
        RECT 1175.860 530.780 1176.120 531.040 ;
        RECT 1175.860 482.840 1176.120 483.100 ;
        RECT 1176.780 482.840 1177.040 483.100 ;
        RECT 1175.400 434.560 1175.660 434.820 ;
        RECT 1175.860 434.220 1176.120 434.480 ;
        RECT 1175.860 338.340 1176.120 338.600 ;
        RECT 1175.400 338.000 1175.660 338.260 ;
        RECT 1175.400 330.860 1175.660 331.120 ;
        RECT 1175.860 330.520 1176.120 330.780 ;
        RECT 1175.860 241.780 1176.120 242.040 ;
        RECT 1175.400 241.440 1175.660 241.700 ;
        RECT 1174.020 207.100 1174.280 207.360 ;
        RECT 1175.400 207.100 1175.660 207.360 ;
        RECT 1174.020 158.820 1174.280 159.080 ;
        RECT 1173.560 158.480 1173.820 158.740 ;
        RECT 1173.560 125.500 1173.820 125.760 ;
        RECT 1175.860 125.500 1176.120 125.760 ;
        RECT 1173.560 62.260 1173.820 62.520 ;
        RECT 1175.860 62.260 1176.120 62.520 ;
        RECT 942.180 18.060 942.440 18.320 ;
        RECT 1173.560 18.060 1173.820 18.320 ;
      LAYER met2 ;
        RECT 1173.470 1100.650 1173.750 1104.000 ;
        RECT 1173.470 1100.510 1174.220 1100.650 ;
        RECT 1173.470 1100.000 1173.750 1100.510 ;
        RECT 1174.080 1028.830 1174.220 1100.510 ;
        RECT 1174.020 1028.510 1174.280 1028.830 ;
        RECT 1174.020 1027.830 1174.280 1028.150 ;
        RECT 1174.080 990.070 1174.220 1027.830 ;
        RECT 1174.020 989.750 1174.280 990.070 ;
        RECT 1175.860 989.750 1176.120 990.070 ;
        RECT 1175.920 821.965 1176.060 989.750 ;
        RECT 1175.850 821.595 1176.130 821.965 ;
        RECT 1175.390 820.915 1175.670 821.285 ;
        RECT 1175.400 820.770 1175.660 820.915 ;
        RECT 1175.860 820.430 1176.120 820.750 ;
        RECT 1175.920 772.810 1176.060 820.430 ;
        RECT 1174.940 772.490 1175.200 772.810 ;
        RECT 1175.860 772.490 1176.120 772.810 ;
        RECT 1175.000 725.290 1175.140 772.490 ;
        RECT 1175.000 725.150 1175.600 725.290 ;
        RECT 1175.460 710.590 1175.600 725.150 ;
        RECT 1175.400 710.270 1175.660 710.590 ;
        RECT 1175.860 709.930 1176.120 710.250 ;
        RECT 1175.920 628.845 1176.060 709.930 ;
        RECT 1175.850 628.475 1176.130 628.845 ;
        RECT 1175.390 627.795 1175.670 628.165 ;
        RECT 1175.400 627.650 1175.660 627.795 ;
        RECT 1175.860 627.310 1176.120 627.630 ;
        RECT 1175.920 532.285 1176.060 627.310 ;
        RECT 1175.850 531.915 1176.130 532.285 ;
        RECT 1175.390 531.235 1175.670 531.605 ;
        RECT 1175.400 531.090 1175.660 531.235 ;
        RECT 1175.860 530.750 1176.120 531.070 ;
        RECT 1175.920 483.130 1176.060 530.750 ;
        RECT 1175.860 482.810 1176.120 483.130 ;
        RECT 1176.780 482.810 1177.040 483.130 ;
        RECT 1176.840 435.045 1176.980 482.810 ;
        RECT 1175.390 434.675 1175.670 435.045 ;
        RECT 1176.770 434.675 1177.050 435.045 ;
        RECT 1175.400 434.530 1175.660 434.675 ;
        RECT 1175.860 434.190 1176.120 434.510 ;
        RECT 1175.920 338.630 1176.060 434.190 ;
        RECT 1175.860 338.310 1176.120 338.630 ;
        RECT 1175.400 337.970 1175.660 338.290 ;
        RECT 1175.460 331.150 1175.600 337.970 ;
        RECT 1175.400 330.830 1175.660 331.150 ;
        RECT 1175.860 330.490 1176.120 330.810 ;
        RECT 1175.920 242.070 1176.060 330.490 ;
        RECT 1175.860 241.750 1176.120 242.070 ;
        RECT 1175.400 241.410 1175.660 241.730 ;
        RECT 1175.460 207.390 1175.600 241.410 ;
        RECT 1174.020 207.070 1174.280 207.390 ;
        RECT 1175.400 207.070 1175.660 207.390 ;
        RECT 1174.080 159.110 1174.220 207.070 ;
        RECT 1174.020 158.790 1174.280 159.110 ;
        RECT 1173.560 158.450 1173.820 158.770 ;
        RECT 1173.620 125.790 1173.760 158.450 ;
        RECT 1173.560 125.470 1173.820 125.790 ;
        RECT 1175.860 125.470 1176.120 125.790 ;
        RECT 1175.920 62.550 1176.060 125.470 ;
        RECT 1173.560 62.230 1173.820 62.550 ;
        RECT 1175.860 62.230 1176.120 62.550 ;
        RECT 1173.620 18.350 1173.760 62.230 ;
        RECT 942.180 18.030 942.440 18.350 ;
        RECT 1173.560 18.030 1173.820 18.350 ;
        RECT 942.240 2.000 942.380 18.030 ;
        RECT 942.030 -4.000 942.590 2.000 ;
      LAYER via2 ;
        RECT 1175.850 821.640 1176.130 821.920 ;
        RECT 1175.390 820.960 1175.670 821.240 ;
        RECT 1175.850 628.520 1176.130 628.800 ;
        RECT 1175.390 627.840 1175.670 628.120 ;
        RECT 1175.850 531.960 1176.130 532.240 ;
        RECT 1175.390 531.280 1175.670 531.560 ;
        RECT 1175.390 434.720 1175.670 435.000 ;
        RECT 1176.770 434.720 1177.050 435.000 ;
      LAYER met3 ;
        RECT 1175.825 821.930 1176.155 821.945 ;
        RECT 1175.150 821.630 1176.155 821.930 ;
        RECT 1175.150 821.265 1175.450 821.630 ;
        RECT 1175.825 821.615 1176.155 821.630 ;
        RECT 1175.150 820.950 1175.695 821.265 ;
        RECT 1175.365 820.935 1175.695 820.950 ;
        RECT 1175.825 628.810 1176.155 628.825 ;
        RECT 1175.150 628.510 1176.155 628.810 ;
        RECT 1175.150 628.145 1175.450 628.510 ;
        RECT 1175.825 628.495 1176.155 628.510 ;
        RECT 1175.150 627.830 1175.695 628.145 ;
        RECT 1175.365 627.815 1175.695 627.830 ;
        RECT 1175.825 532.250 1176.155 532.265 ;
        RECT 1175.150 531.950 1176.155 532.250 ;
        RECT 1175.150 531.585 1175.450 531.950 ;
        RECT 1175.825 531.935 1176.155 531.950 ;
        RECT 1175.150 531.270 1175.695 531.585 ;
        RECT 1175.365 531.255 1175.695 531.270 ;
        RECT 1175.365 435.010 1175.695 435.025 ;
        RECT 1176.745 435.010 1177.075 435.025 ;
        RECT 1175.365 434.710 1177.075 435.010 ;
        RECT 1175.365 434.695 1175.695 434.710 ;
        RECT 1176.745 434.695 1177.075 434.710 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1176.365 579.785 1176.535 593.555 ;
        RECT 1176.365 483.225 1176.535 496.995 ;
        RECT 1176.365 386.325 1176.535 400.435 ;
      LAYER mcon ;
        RECT 1176.365 593.385 1176.535 593.555 ;
        RECT 1176.365 496.825 1176.535 496.995 ;
        RECT 1176.365 400.265 1176.535 400.435 ;
      LAYER met1 ;
        RECT 1174.910 990.320 1175.230 990.380 ;
        RECT 1178.130 990.320 1178.450 990.380 ;
        RECT 1174.910 990.180 1178.450 990.320 ;
        RECT 1174.910 990.120 1175.230 990.180 ;
        RECT 1178.130 990.120 1178.450 990.180 ;
        RECT 1174.910 917.900 1175.230 917.960 ;
        RECT 1175.370 917.900 1175.690 917.960 ;
        RECT 1174.910 917.760 1175.690 917.900 ;
        RECT 1174.910 917.700 1175.230 917.760 ;
        RECT 1175.370 917.700 1175.690 917.760 ;
        RECT 1176.290 821.340 1176.610 821.400 ;
        RECT 1176.750 821.340 1177.070 821.400 ;
        RECT 1176.290 821.200 1177.070 821.340 ;
        RECT 1176.290 821.140 1176.610 821.200 ;
        RECT 1176.750 821.140 1177.070 821.200 ;
        RECT 1174.910 714.240 1175.230 714.300 ;
        RECT 1176.290 714.240 1176.610 714.300 ;
        RECT 1174.910 714.100 1176.610 714.240 ;
        RECT 1174.910 714.040 1175.230 714.100 ;
        RECT 1176.290 714.040 1176.610 714.100 ;
        RECT 1176.290 593.540 1176.610 593.600 ;
        RECT 1176.095 593.400 1176.610 593.540 ;
        RECT 1176.290 593.340 1176.610 593.400 ;
        RECT 1176.290 579.940 1176.610 580.000 ;
        RECT 1176.095 579.800 1176.610 579.940 ;
        RECT 1176.290 579.740 1176.610 579.800 ;
        RECT 1176.290 496.980 1176.610 497.040 ;
        RECT 1176.095 496.840 1176.610 496.980 ;
        RECT 1176.290 496.780 1176.610 496.840 ;
        RECT 1176.290 483.380 1176.610 483.440 ;
        RECT 1176.095 483.240 1176.610 483.380 ;
        RECT 1176.290 483.180 1176.610 483.240 ;
        RECT 1176.290 400.420 1176.610 400.480 ;
        RECT 1176.095 400.280 1176.610 400.420 ;
        RECT 1176.290 400.220 1176.610 400.280 ;
        RECT 1176.290 386.480 1176.610 386.540 ;
        RECT 1176.095 386.340 1176.610 386.480 ;
        RECT 1176.290 386.280 1176.610 386.340 ;
        RECT 1174.910 327.660 1175.230 327.720 ;
        RECT 1176.290 327.660 1176.610 327.720 ;
        RECT 1174.910 327.520 1176.610 327.660 ;
        RECT 1174.910 327.460 1175.230 327.520 ;
        RECT 1176.290 327.460 1176.610 327.520 ;
        RECT 1174.910 303.180 1175.230 303.240 ;
        RECT 1176.290 303.180 1176.610 303.240 ;
        RECT 1174.910 303.040 1176.610 303.180 ;
        RECT 1174.910 302.980 1175.230 303.040 ;
        RECT 1176.290 302.980 1176.610 303.040 ;
        RECT 1176.290 255.380 1176.610 255.640 ;
        RECT 1176.380 255.240 1176.520 255.380 ;
        RECT 1176.750 255.240 1177.070 255.300 ;
        RECT 1176.380 255.100 1177.070 255.240 ;
        RECT 1176.750 255.040 1177.070 255.100 ;
        RECT 1175.370 193.020 1175.690 193.080 ;
        RECT 1176.290 193.020 1176.610 193.080 ;
        RECT 1175.370 192.880 1176.610 193.020 ;
        RECT 1175.370 192.820 1175.690 192.880 ;
        RECT 1176.290 192.820 1176.610 192.880 ;
        RECT 960.090 19.280 960.410 19.340 ;
        RECT 1176.290 19.280 1176.610 19.340 ;
        RECT 960.090 19.140 1176.610 19.280 ;
        RECT 960.090 19.080 960.410 19.140 ;
        RECT 1176.290 19.080 1176.610 19.140 ;
      LAYER via ;
        RECT 1174.940 990.120 1175.200 990.380 ;
        RECT 1178.160 990.120 1178.420 990.380 ;
        RECT 1174.940 917.700 1175.200 917.960 ;
        RECT 1175.400 917.700 1175.660 917.960 ;
        RECT 1176.320 821.140 1176.580 821.400 ;
        RECT 1176.780 821.140 1177.040 821.400 ;
        RECT 1174.940 714.040 1175.200 714.300 ;
        RECT 1176.320 714.040 1176.580 714.300 ;
        RECT 1176.320 593.340 1176.580 593.600 ;
        RECT 1176.320 579.740 1176.580 580.000 ;
        RECT 1176.320 496.780 1176.580 497.040 ;
        RECT 1176.320 483.180 1176.580 483.440 ;
        RECT 1176.320 400.220 1176.580 400.480 ;
        RECT 1176.320 386.280 1176.580 386.540 ;
        RECT 1174.940 327.460 1175.200 327.720 ;
        RECT 1176.320 327.460 1176.580 327.720 ;
        RECT 1174.940 302.980 1175.200 303.240 ;
        RECT 1176.320 302.980 1176.580 303.240 ;
        RECT 1176.320 255.380 1176.580 255.640 ;
        RECT 1176.780 255.040 1177.040 255.300 ;
        RECT 1175.400 192.820 1175.660 193.080 ;
        RECT 1176.320 192.820 1176.580 193.080 ;
        RECT 960.120 19.080 960.380 19.340 ;
        RECT 1176.320 19.080 1176.580 19.340 ;
      LAYER met2 ;
        RECT 1179.450 1101.330 1179.730 1104.000 ;
        RECT 1177.760 1101.190 1179.730 1101.330 ;
        RECT 1177.760 1062.570 1177.900 1101.190 ;
        RECT 1179.450 1100.000 1179.730 1101.190 ;
        RECT 1177.760 1062.430 1178.360 1062.570 ;
        RECT 1178.220 990.410 1178.360 1062.430 ;
        RECT 1174.940 990.090 1175.200 990.410 ;
        RECT 1178.160 990.090 1178.420 990.410 ;
        RECT 1175.000 917.990 1175.140 990.090 ;
        RECT 1174.940 917.670 1175.200 917.990 ;
        RECT 1175.400 917.845 1175.660 917.990 ;
        RECT 1175.390 917.475 1175.670 917.845 ;
        RECT 1176.770 917.475 1177.050 917.845 ;
        RECT 1176.840 821.430 1176.980 917.475 ;
        RECT 1176.320 821.110 1176.580 821.430 ;
        RECT 1176.780 821.110 1177.040 821.430 ;
        RECT 1176.380 714.330 1176.520 821.110 ;
        RECT 1174.940 714.010 1175.200 714.330 ;
        RECT 1176.320 714.010 1176.580 714.330 ;
        RECT 1175.000 690.045 1175.140 714.010 ;
        RECT 1174.930 689.675 1175.210 690.045 ;
        RECT 1176.310 689.675 1176.590 690.045 ;
        RECT 1176.380 593.630 1176.520 689.675 ;
        RECT 1176.320 593.310 1176.580 593.630 ;
        RECT 1176.320 579.710 1176.580 580.030 ;
        RECT 1176.380 497.070 1176.520 579.710 ;
        RECT 1176.320 496.750 1176.580 497.070 ;
        RECT 1176.320 483.150 1176.580 483.470 ;
        RECT 1176.380 400.510 1176.520 483.150 ;
        RECT 1176.320 400.190 1176.580 400.510 ;
        RECT 1176.320 386.250 1176.580 386.570 ;
        RECT 1176.380 327.750 1176.520 386.250 ;
        RECT 1174.940 327.430 1175.200 327.750 ;
        RECT 1176.320 327.430 1176.580 327.750 ;
        RECT 1175.000 303.270 1175.140 327.430 ;
        RECT 1174.940 302.950 1175.200 303.270 ;
        RECT 1176.320 302.950 1176.580 303.270 ;
        RECT 1176.380 255.670 1176.520 302.950 ;
        RECT 1176.320 255.350 1176.580 255.670 ;
        RECT 1176.780 255.010 1177.040 255.330 ;
        RECT 1176.840 207.245 1176.980 255.010 ;
        RECT 1174.930 206.875 1175.210 207.245 ;
        RECT 1176.770 206.875 1177.050 207.245 ;
        RECT 1175.000 206.450 1175.140 206.875 ;
        RECT 1175.000 206.310 1175.600 206.450 ;
        RECT 1175.460 193.110 1175.600 206.310 ;
        RECT 1175.400 192.790 1175.660 193.110 ;
        RECT 1176.320 192.790 1176.580 193.110 ;
        RECT 1176.380 19.370 1176.520 192.790 ;
        RECT 960.120 19.050 960.380 19.370 ;
        RECT 1176.320 19.050 1176.580 19.370 ;
        RECT 960.180 2.000 960.320 19.050 ;
        RECT 959.970 -4.000 960.530 2.000 ;
      LAYER via2 ;
        RECT 1175.390 917.520 1175.670 917.800 ;
        RECT 1176.770 917.520 1177.050 917.800 ;
        RECT 1174.930 689.720 1175.210 690.000 ;
        RECT 1176.310 689.720 1176.590 690.000 ;
        RECT 1174.930 206.920 1175.210 207.200 ;
        RECT 1176.770 206.920 1177.050 207.200 ;
      LAYER met3 ;
        RECT 1175.365 917.810 1175.695 917.825 ;
        RECT 1176.745 917.810 1177.075 917.825 ;
        RECT 1175.365 917.510 1177.075 917.810 ;
        RECT 1175.365 917.495 1175.695 917.510 ;
        RECT 1176.745 917.495 1177.075 917.510 ;
        RECT 1174.905 690.010 1175.235 690.025 ;
        RECT 1176.285 690.010 1176.615 690.025 ;
        RECT 1174.905 689.710 1176.615 690.010 ;
        RECT 1174.905 689.695 1175.235 689.710 ;
        RECT 1176.285 689.695 1176.615 689.710 ;
        RECT 1174.905 207.210 1175.235 207.225 ;
        RECT 1176.745 207.210 1177.075 207.225 ;
        RECT 1174.905 206.910 1177.075 207.210 ;
        RECT 1174.905 206.895 1175.235 206.910 ;
        RECT 1176.745 206.895 1177.075 206.910 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1126.225 18.785 1126.395 19.635 ;
      LAYER mcon ;
        RECT 1126.225 19.465 1126.395 19.635 ;
      LAYER met1 ;
        RECT 1179.970 1052.200 1180.290 1052.260 ;
        RECT 1184.110 1052.200 1184.430 1052.260 ;
        RECT 1179.970 1052.060 1184.430 1052.200 ;
        RECT 1179.970 1052.000 1180.290 1052.060 ;
        RECT 1184.110 1052.000 1184.430 1052.060 ;
        RECT 978.030 19.620 978.350 19.680 ;
        RECT 1126.165 19.620 1126.455 19.665 ;
        RECT 978.030 19.480 1126.455 19.620 ;
        RECT 978.030 19.420 978.350 19.480 ;
        RECT 1126.165 19.435 1126.455 19.480 ;
        RECT 1126.165 18.940 1126.455 18.985 ;
        RECT 1179.970 18.940 1180.290 19.000 ;
        RECT 1126.165 18.800 1180.290 18.940 ;
        RECT 1126.165 18.755 1126.455 18.800 ;
        RECT 1179.970 18.740 1180.290 18.800 ;
      LAYER via ;
        RECT 1180.000 1052.000 1180.260 1052.260 ;
        RECT 1184.140 1052.000 1184.400 1052.260 ;
        RECT 978.060 19.420 978.320 19.680 ;
        RECT 1180.000 18.740 1180.260 19.000 ;
      LAYER met2 ;
        RECT 1185.430 1100.650 1185.710 1104.000 ;
        RECT 1184.200 1100.510 1185.710 1100.650 ;
        RECT 1184.200 1052.290 1184.340 1100.510 ;
        RECT 1185.430 1100.000 1185.710 1100.510 ;
        RECT 1180.000 1051.970 1180.260 1052.290 ;
        RECT 1184.140 1051.970 1184.400 1052.290 ;
        RECT 978.060 19.390 978.320 19.710 ;
        RECT 978.120 2.000 978.260 19.390 ;
        RECT 1180.060 19.030 1180.200 1051.970 ;
        RECT 1180.000 18.710 1180.260 19.030 ;
        RECT 977.910 -4.000 978.470 2.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1070.030 1072.940 1070.350 1073.000 ;
        RECT 1073.710 1072.940 1074.030 1073.000 ;
        RECT 1070.030 1072.800 1074.030 1072.940 ;
        RECT 1070.030 1072.740 1070.350 1072.800 ;
        RECT 1073.710 1072.740 1074.030 1072.800 ;
        RECT 656.950 47.160 657.270 47.220 ;
        RECT 1070.030 47.160 1070.350 47.220 ;
        RECT 656.950 47.020 1070.350 47.160 ;
        RECT 656.950 46.960 657.270 47.020 ;
        RECT 1070.030 46.960 1070.350 47.020 ;
      LAYER via ;
        RECT 1070.060 1072.740 1070.320 1073.000 ;
        RECT 1073.740 1072.740 1074.000 1073.000 ;
        RECT 656.980 46.960 657.240 47.220 ;
        RECT 1070.060 46.960 1070.320 47.220 ;
      LAYER met2 ;
        RECT 1075.490 1100.650 1075.770 1104.000 ;
        RECT 1073.800 1100.510 1075.770 1100.650 ;
        RECT 1073.800 1073.030 1073.940 1100.510 ;
        RECT 1075.490 1100.000 1075.770 1100.510 ;
        RECT 1070.060 1072.710 1070.320 1073.030 ;
        RECT 1073.740 1072.710 1074.000 1073.030 ;
        RECT 1070.120 47.250 1070.260 1072.710 ;
        RECT 656.980 46.930 657.240 47.250 ;
        RECT 1070.060 46.930 1070.320 47.250 ;
        RECT 657.040 2.000 657.180 46.930 ;
        RECT 656.830 -4.000 657.390 2.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1017.590 1087.220 1017.910 1087.280 ;
        RECT 1191.470 1087.220 1191.790 1087.280 ;
        RECT 1017.590 1087.080 1191.790 1087.220 ;
        RECT 1017.590 1087.020 1017.910 1087.080 ;
        RECT 1191.470 1087.020 1191.790 1087.080 ;
        RECT 995.970 20.640 996.290 20.700 ;
        RECT 1017.590 20.640 1017.910 20.700 ;
        RECT 995.970 20.500 1017.910 20.640 ;
        RECT 995.970 20.440 996.290 20.500 ;
        RECT 1017.590 20.440 1017.910 20.500 ;
      LAYER via ;
        RECT 1017.620 1087.020 1017.880 1087.280 ;
        RECT 1191.500 1087.020 1191.760 1087.280 ;
        RECT 996.000 20.440 996.260 20.700 ;
        RECT 1017.620 20.440 1017.880 20.700 ;
      LAYER met2 ;
        RECT 1191.410 1100.580 1191.690 1104.000 ;
        RECT 1191.410 1100.000 1191.700 1100.580 ;
        RECT 1191.560 1087.310 1191.700 1100.000 ;
        RECT 1017.620 1086.990 1017.880 1087.310 ;
        RECT 1191.500 1086.990 1191.760 1087.310 ;
        RECT 1017.680 20.730 1017.820 1086.990 ;
        RECT 996.000 20.410 996.260 20.730 ;
        RECT 1017.620 20.410 1017.880 20.730 ;
        RECT 996.060 2.000 996.200 20.410 ;
        RECT 995.850 -4.000 996.410 2.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1045.190 1088.920 1045.510 1088.980 ;
        RECT 1197.910 1088.920 1198.230 1088.980 ;
        RECT 1045.190 1088.780 1198.230 1088.920 ;
        RECT 1045.190 1088.720 1045.510 1088.780 ;
        RECT 1197.910 1088.720 1198.230 1088.780 ;
        RECT 1013.450 15.540 1013.770 15.600 ;
        RECT 1045.190 15.540 1045.510 15.600 ;
        RECT 1013.450 15.400 1045.510 15.540 ;
        RECT 1013.450 15.340 1013.770 15.400 ;
        RECT 1045.190 15.340 1045.510 15.400 ;
      LAYER via ;
        RECT 1045.220 1088.720 1045.480 1088.980 ;
        RECT 1197.940 1088.720 1198.200 1088.980 ;
        RECT 1013.480 15.340 1013.740 15.600 ;
        RECT 1045.220 15.340 1045.480 15.600 ;
      LAYER met2 ;
        RECT 1197.850 1100.580 1198.130 1104.000 ;
        RECT 1197.850 1100.000 1198.140 1100.580 ;
        RECT 1198.000 1089.010 1198.140 1100.000 ;
        RECT 1045.220 1088.690 1045.480 1089.010 ;
        RECT 1197.940 1088.690 1198.200 1089.010 ;
        RECT 1045.280 15.630 1045.420 1088.690 ;
        RECT 1013.480 15.310 1013.740 15.630 ;
        RECT 1045.220 15.310 1045.480 15.630 ;
        RECT 1013.540 2.000 1013.680 15.310 ;
        RECT 1013.330 -4.000 1013.890 2.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1059.525 1014.305 1059.695 1062.415 ;
        RECT 1059.525 772.905 1059.695 855.355 ;
        RECT 1059.525 676.345 1059.695 724.455 ;
        RECT 1059.525 579.785 1059.695 627.895 ;
        RECT 1059.525 500.225 1059.695 531.335 ;
      LAYER mcon ;
        RECT 1059.525 1062.245 1059.695 1062.415 ;
        RECT 1059.525 855.185 1059.695 855.355 ;
        RECT 1059.525 724.285 1059.695 724.455 ;
        RECT 1059.525 627.725 1059.695 627.895 ;
        RECT 1059.525 531.165 1059.695 531.335 ;
      LAYER met1 ;
        RECT 1061.750 1089.260 1062.070 1089.320 ;
        RECT 1203.890 1089.260 1204.210 1089.320 ;
        RECT 1061.750 1089.120 1204.210 1089.260 ;
        RECT 1061.750 1089.060 1062.070 1089.120 ;
        RECT 1203.890 1089.060 1204.210 1089.120 ;
        RECT 1059.450 1062.400 1059.770 1062.460 ;
        RECT 1059.255 1062.260 1059.770 1062.400 ;
        RECT 1059.450 1062.200 1059.770 1062.260 ;
        RECT 1059.465 1014.460 1059.755 1014.505 ;
        RECT 1059.910 1014.460 1060.230 1014.520 ;
        RECT 1059.465 1014.320 1060.230 1014.460 ;
        RECT 1059.465 1014.275 1059.755 1014.320 ;
        RECT 1059.910 1014.260 1060.230 1014.320 ;
        RECT 1058.530 883.560 1058.850 883.620 ;
        RECT 1059.910 883.560 1060.230 883.620 ;
        RECT 1058.530 883.420 1060.230 883.560 ;
        RECT 1058.530 883.360 1058.850 883.420 ;
        RECT 1059.910 883.360 1060.230 883.420 ;
        RECT 1058.530 855.340 1058.850 855.400 ;
        RECT 1059.465 855.340 1059.755 855.385 ;
        RECT 1058.530 855.200 1059.755 855.340 ;
        RECT 1058.530 855.140 1058.850 855.200 ;
        RECT 1059.465 855.155 1059.755 855.200 ;
        RECT 1059.450 773.060 1059.770 773.120 ;
        RECT 1059.255 772.920 1059.770 773.060 ;
        RECT 1059.450 772.860 1059.770 772.920 ;
        RECT 1059.450 738.180 1059.770 738.440 ;
        RECT 1059.540 738.040 1059.680 738.180 ;
        RECT 1059.910 738.040 1060.230 738.100 ;
        RECT 1059.540 737.900 1060.230 738.040 ;
        RECT 1059.910 737.840 1060.230 737.900 ;
        RECT 1059.465 724.440 1059.755 724.485 ;
        RECT 1059.910 724.440 1060.230 724.500 ;
        RECT 1059.465 724.300 1060.230 724.440 ;
        RECT 1059.465 724.255 1059.755 724.300 ;
        RECT 1059.910 724.240 1060.230 724.300 ;
        RECT 1059.450 676.500 1059.770 676.560 ;
        RECT 1059.255 676.360 1059.770 676.500 ;
        RECT 1059.450 676.300 1059.770 676.360 ;
        RECT 1059.450 641.620 1059.770 641.880 ;
        RECT 1059.540 641.480 1059.680 641.620 ;
        RECT 1059.910 641.480 1060.230 641.540 ;
        RECT 1059.540 641.340 1060.230 641.480 ;
        RECT 1059.910 641.280 1060.230 641.340 ;
        RECT 1059.465 627.880 1059.755 627.925 ;
        RECT 1059.910 627.880 1060.230 627.940 ;
        RECT 1059.465 627.740 1060.230 627.880 ;
        RECT 1059.465 627.695 1059.755 627.740 ;
        RECT 1059.910 627.680 1060.230 627.740 ;
        RECT 1059.450 579.940 1059.770 580.000 ;
        RECT 1059.255 579.800 1059.770 579.940 ;
        RECT 1059.450 579.740 1059.770 579.800 ;
        RECT 1059.450 545.060 1059.770 545.320 ;
        RECT 1059.540 544.920 1059.680 545.060 ;
        RECT 1059.910 544.920 1060.230 544.980 ;
        RECT 1059.540 544.780 1060.230 544.920 ;
        RECT 1059.910 544.720 1060.230 544.780 ;
        RECT 1059.465 531.320 1059.755 531.365 ;
        RECT 1059.910 531.320 1060.230 531.380 ;
        RECT 1059.465 531.180 1060.230 531.320 ;
        RECT 1059.465 531.135 1059.755 531.180 ;
        RECT 1059.910 531.120 1060.230 531.180 ;
        RECT 1059.465 500.380 1059.755 500.425 ;
        RECT 1059.910 500.380 1060.230 500.440 ;
        RECT 1059.465 500.240 1060.230 500.380 ;
        RECT 1059.465 500.195 1059.755 500.240 ;
        RECT 1059.910 500.180 1060.230 500.240 ;
        RECT 1059.450 434.760 1059.770 434.820 ;
        RECT 1059.910 434.760 1060.230 434.820 ;
        RECT 1059.450 434.620 1060.230 434.760 ;
        RECT 1059.450 434.560 1059.770 434.620 ;
        RECT 1059.910 434.560 1060.230 434.620 ;
        RECT 1059.450 352.280 1059.770 352.540 ;
        RECT 1059.540 351.860 1059.680 352.280 ;
        RECT 1059.450 351.600 1059.770 351.860 ;
        RECT 1059.450 241.300 1059.770 241.360 ;
        RECT 1059.910 241.300 1060.230 241.360 ;
        RECT 1059.450 241.160 1060.230 241.300 ;
        RECT 1059.450 241.100 1059.770 241.160 ;
        RECT 1059.910 241.100 1060.230 241.160 ;
        RECT 1059.450 193.020 1059.770 193.080 ;
        RECT 1059.910 193.020 1060.230 193.080 ;
        RECT 1059.450 192.880 1060.230 193.020 ;
        RECT 1059.450 192.820 1059.770 192.880 ;
        RECT 1059.910 192.820 1060.230 192.880 ;
        RECT 1060.370 137.940 1060.690 138.000 ;
        RECT 1060.830 137.940 1061.150 138.000 ;
        RECT 1060.370 137.800 1061.150 137.940 ;
        RECT 1060.370 137.740 1060.690 137.800 ;
        RECT 1060.830 137.740 1061.150 137.800 ;
        RECT 1059.450 62.120 1059.770 62.180 ;
        RECT 1060.830 62.120 1061.150 62.180 ;
        RECT 1059.450 61.980 1061.150 62.120 ;
        RECT 1059.450 61.920 1059.770 61.980 ;
        RECT 1060.830 61.920 1061.150 61.980 ;
        RECT 1031.390 20.300 1031.710 20.360 ;
        RECT 1059.450 20.300 1059.770 20.360 ;
        RECT 1031.390 20.160 1059.770 20.300 ;
        RECT 1031.390 20.100 1031.710 20.160 ;
        RECT 1059.450 20.100 1059.770 20.160 ;
      LAYER via ;
        RECT 1061.780 1089.060 1062.040 1089.320 ;
        RECT 1203.920 1089.060 1204.180 1089.320 ;
        RECT 1059.480 1062.200 1059.740 1062.460 ;
        RECT 1059.940 1014.260 1060.200 1014.520 ;
        RECT 1058.560 883.360 1058.820 883.620 ;
        RECT 1059.940 883.360 1060.200 883.620 ;
        RECT 1058.560 855.140 1058.820 855.400 ;
        RECT 1059.480 772.860 1059.740 773.120 ;
        RECT 1059.480 738.180 1059.740 738.440 ;
        RECT 1059.940 737.840 1060.200 738.100 ;
        RECT 1059.940 724.240 1060.200 724.500 ;
        RECT 1059.480 676.300 1059.740 676.560 ;
        RECT 1059.480 641.620 1059.740 641.880 ;
        RECT 1059.940 641.280 1060.200 641.540 ;
        RECT 1059.940 627.680 1060.200 627.940 ;
        RECT 1059.480 579.740 1059.740 580.000 ;
        RECT 1059.480 545.060 1059.740 545.320 ;
        RECT 1059.940 544.720 1060.200 544.980 ;
        RECT 1059.940 531.120 1060.200 531.380 ;
        RECT 1059.940 500.180 1060.200 500.440 ;
        RECT 1059.480 434.560 1059.740 434.820 ;
        RECT 1059.940 434.560 1060.200 434.820 ;
        RECT 1059.480 352.280 1059.740 352.540 ;
        RECT 1059.480 351.600 1059.740 351.860 ;
        RECT 1059.480 241.100 1059.740 241.360 ;
        RECT 1059.940 241.100 1060.200 241.360 ;
        RECT 1059.480 192.820 1059.740 193.080 ;
        RECT 1059.940 192.820 1060.200 193.080 ;
        RECT 1060.400 137.740 1060.660 138.000 ;
        RECT 1060.860 137.740 1061.120 138.000 ;
        RECT 1059.480 61.920 1059.740 62.180 ;
        RECT 1060.860 61.920 1061.120 62.180 ;
        RECT 1031.420 20.100 1031.680 20.360 ;
        RECT 1059.480 20.100 1059.740 20.360 ;
      LAYER met2 ;
        RECT 1203.830 1100.580 1204.110 1104.000 ;
        RECT 1203.830 1100.000 1204.120 1100.580 ;
        RECT 1203.980 1089.350 1204.120 1100.000 ;
        RECT 1061.780 1089.030 1062.040 1089.350 ;
        RECT 1203.920 1089.030 1204.180 1089.350 ;
        RECT 1061.840 1063.365 1061.980 1089.030 ;
        RECT 1061.770 1062.995 1062.050 1063.365 ;
        RECT 1059.470 1062.485 1059.750 1062.855 ;
        RECT 1059.480 1062.170 1059.740 1062.485 ;
        RECT 1059.940 1014.230 1060.200 1014.550 ;
        RECT 1060.000 978.930 1060.140 1014.230 ;
        RECT 1059.540 978.790 1060.140 978.930 ;
        RECT 1059.540 910.930 1059.680 978.790 ;
        RECT 1059.540 910.790 1060.140 910.930 ;
        RECT 1060.000 883.650 1060.140 910.790 ;
        RECT 1058.560 883.330 1058.820 883.650 ;
        RECT 1059.940 883.330 1060.200 883.650 ;
        RECT 1058.620 855.430 1058.760 883.330 ;
        RECT 1058.560 855.110 1058.820 855.430 ;
        RECT 1059.480 772.830 1059.740 773.150 ;
        RECT 1059.540 738.470 1059.680 772.830 ;
        RECT 1059.480 738.150 1059.740 738.470 ;
        RECT 1059.940 737.810 1060.200 738.130 ;
        RECT 1060.000 724.530 1060.140 737.810 ;
        RECT 1059.940 724.210 1060.200 724.530 ;
        RECT 1059.480 676.270 1059.740 676.590 ;
        RECT 1059.540 641.910 1059.680 676.270 ;
        RECT 1059.480 641.590 1059.740 641.910 ;
        RECT 1059.940 641.250 1060.200 641.570 ;
        RECT 1060.000 627.970 1060.140 641.250 ;
        RECT 1059.940 627.650 1060.200 627.970 ;
        RECT 1059.480 579.710 1059.740 580.030 ;
        RECT 1059.540 545.350 1059.680 579.710 ;
        RECT 1059.480 545.030 1059.740 545.350 ;
        RECT 1059.940 544.690 1060.200 545.010 ;
        RECT 1060.000 531.410 1060.140 544.690 ;
        RECT 1059.940 531.090 1060.200 531.410 ;
        RECT 1059.940 500.150 1060.200 500.470 ;
        RECT 1060.000 434.850 1060.140 500.150 ;
        RECT 1059.480 434.530 1059.740 434.850 ;
        RECT 1059.940 434.530 1060.200 434.850 ;
        RECT 1059.540 352.570 1059.680 434.530 ;
        RECT 1059.480 352.250 1059.740 352.570 ;
        RECT 1059.480 351.570 1059.740 351.890 ;
        RECT 1059.540 290.885 1059.680 351.570 ;
        RECT 1059.470 290.515 1059.750 290.885 ;
        RECT 1059.930 289.155 1060.210 289.525 ;
        RECT 1060.000 241.390 1060.140 289.155 ;
        RECT 1059.480 241.070 1059.740 241.390 ;
        RECT 1059.940 241.070 1060.200 241.390 ;
        RECT 1059.540 193.110 1059.680 241.070 ;
        RECT 1059.480 192.790 1059.740 193.110 ;
        RECT 1059.940 192.790 1060.200 193.110 ;
        RECT 1060.000 168.370 1060.140 192.790 ;
        RECT 1060.000 168.230 1060.600 168.370 ;
        RECT 1060.460 138.030 1060.600 168.230 ;
        RECT 1060.400 137.710 1060.660 138.030 ;
        RECT 1060.860 137.710 1061.120 138.030 ;
        RECT 1060.920 62.210 1061.060 137.710 ;
        RECT 1059.480 61.890 1059.740 62.210 ;
        RECT 1060.860 61.890 1061.120 62.210 ;
        RECT 1059.540 20.390 1059.680 61.890 ;
        RECT 1031.420 20.070 1031.680 20.390 ;
        RECT 1059.480 20.070 1059.740 20.390 ;
        RECT 1031.480 2.000 1031.620 20.070 ;
        RECT 1031.270 -4.000 1031.830 2.000 ;
      LAYER via2 ;
        RECT 1061.770 1063.040 1062.050 1063.320 ;
        RECT 1059.470 1062.530 1059.750 1062.810 ;
        RECT 1059.470 290.560 1059.750 290.840 ;
        RECT 1059.930 289.200 1060.210 289.480 ;
      LAYER met3 ;
        RECT 1061.745 1063.330 1062.075 1063.345 ;
        RECT 1060.150 1063.030 1062.075 1063.330 ;
        RECT 1059.445 1062.820 1059.775 1062.835 ;
        RECT 1060.150 1062.820 1060.450 1063.030 ;
        RECT 1061.745 1063.015 1062.075 1063.030 ;
        RECT 1059.445 1062.520 1060.450 1062.820 ;
        RECT 1059.445 1062.505 1059.775 1062.520 ;
        RECT 1059.445 290.850 1059.775 290.865 ;
        RECT 1059.230 290.535 1059.775 290.850 ;
        RECT 1059.230 289.490 1059.530 290.535 ;
        RECT 1059.905 289.490 1060.235 289.505 ;
        RECT 1059.230 289.190 1060.235 289.490 ;
        RECT 1059.905 289.175 1060.235 289.190 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1124.845 16.235 1125.015 16.915 ;
        RECT 1124.845 16.065 1125.475 16.235 ;
        RECT 1143.705 16.065 1143.875 17.255 ;
      LAYER mcon ;
        RECT 1143.705 17.085 1143.875 17.255 ;
        RECT 1124.845 16.745 1125.015 16.915 ;
        RECT 1125.305 16.065 1125.475 16.235 ;
      LAYER met1 ;
        RECT 1162.490 1084.160 1162.810 1084.220 ;
        RECT 1209.870 1084.160 1210.190 1084.220 ;
        RECT 1162.490 1084.020 1210.190 1084.160 ;
        RECT 1162.490 1083.960 1162.810 1084.020 ;
        RECT 1209.870 1083.960 1210.190 1084.020 ;
        RECT 1143.645 17.240 1143.935 17.285 ;
        RECT 1162.030 17.240 1162.350 17.300 ;
        RECT 1143.645 17.100 1162.350 17.240 ;
        RECT 1143.645 17.055 1143.935 17.100 ;
        RECT 1162.030 17.040 1162.350 17.100 ;
        RECT 1124.785 16.900 1125.075 16.945 ;
        RECT 1124.400 16.760 1125.075 16.900 ;
        RECT 1049.330 16.220 1049.650 16.280 ;
        RECT 1124.400 16.220 1124.540 16.760 ;
        RECT 1124.785 16.715 1125.075 16.760 ;
        RECT 1049.330 16.080 1124.540 16.220 ;
        RECT 1125.245 16.220 1125.535 16.265 ;
        RECT 1143.645 16.220 1143.935 16.265 ;
        RECT 1125.245 16.080 1143.935 16.220 ;
        RECT 1049.330 16.020 1049.650 16.080 ;
        RECT 1125.245 16.035 1125.535 16.080 ;
        RECT 1143.645 16.035 1143.935 16.080 ;
      LAYER via ;
        RECT 1162.520 1083.960 1162.780 1084.220 ;
        RECT 1209.900 1083.960 1210.160 1084.220 ;
        RECT 1162.060 17.040 1162.320 17.300 ;
        RECT 1049.360 16.020 1049.620 16.280 ;
      LAYER met2 ;
        RECT 1209.810 1100.580 1210.090 1104.000 ;
        RECT 1209.810 1100.000 1210.100 1100.580 ;
        RECT 1209.960 1084.250 1210.100 1100.000 ;
        RECT 1162.520 1083.930 1162.780 1084.250 ;
        RECT 1209.900 1083.930 1210.160 1084.250 ;
        RECT 1162.580 18.090 1162.720 1083.930 ;
        RECT 1162.120 17.950 1162.720 18.090 ;
        RECT 1162.120 17.330 1162.260 17.950 ;
        RECT 1162.060 17.010 1162.320 17.330 ;
        RECT 1049.360 15.990 1049.620 16.310 ;
        RECT 1049.420 2.000 1049.560 15.990 ;
        RECT 1049.210 -4.000 1049.770 2.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1173.605 19.805 1174.235 19.975 ;
        RECT 1174.065 18.445 1174.235 19.805 ;
      LAYER met1 ;
        RECT 1067.270 19.960 1067.590 20.020 ;
        RECT 1173.545 19.960 1173.835 20.005 ;
        RECT 1067.270 19.820 1173.835 19.960 ;
        RECT 1067.270 19.760 1067.590 19.820 ;
        RECT 1173.545 19.775 1173.835 19.820 ;
        RECT 1174.005 18.600 1174.295 18.645 ;
        RECT 1215.390 18.600 1215.710 18.660 ;
        RECT 1174.005 18.460 1215.710 18.600 ;
        RECT 1174.005 18.415 1174.295 18.460 ;
        RECT 1215.390 18.400 1215.710 18.460 ;
      LAYER via ;
        RECT 1067.300 19.760 1067.560 20.020 ;
        RECT 1215.420 18.400 1215.680 18.660 ;
      LAYER met2 ;
        RECT 1216.250 1100.650 1216.530 1104.000 ;
        RECT 1215.480 1100.510 1216.530 1100.650 ;
        RECT 1067.300 19.730 1067.560 20.050 ;
        RECT 1067.360 2.000 1067.500 19.730 ;
        RECT 1215.480 18.690 1215.620 1100.510 ;
        RECT 1216.250 1100.000 1216.530 1100.510 ;
        RECT 1215.420 18.370 1215.680 18.690 ;
        RECT 1067.150 -4.000 1067.710 2.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1119.800 1090.140 1123.620 1090.280 ;
        RECT 1093.490 1089.940 1093.810 1090.000 ;
        RECT 1119.800 1089.940 1119.940 1090.140 ;
        RECT 1093.490 1089.800 1119.940 1089.940 ;
        RECT 1123.480 1089.940 1123.620 1090.140 ;
        RECT 1222.290 1089.940 1222.610 1090.000 ;
        RECT 1123.480 1089.800 1222.610 1089.940 ;
        RECT 1093.490 1089.740 1093.810 1089.800 ;
        RECT 1222.290 1089.740 1222.610 1089.800 ;
        RECT 1085.210 20.640 1085.530 20.700 ;
        RECT 1093.490 20.640 1093.810 20.700 ;
        RECT 1085.210 20.500 1093.810 20.640 ;
        RECT 1085.210 20.440 1085.530 20.500 ;
        RECT 1093.490 20.440 1093.810 20.500 ;
      LAYER via ;
        RECT 1093.520 1089.740 1093.780 1090.000 ;
        RECT 1222.320 1089.740 1222.580 1090.000 ;
        RECT 1085.240 20.440 1085.500 20.700 ;
        RECT 1093.520 20.440 1093.780 20.700 ;
      LAYER met2 ;
        RECT 1222.230 1100.580 1222.510 1104.000 ;
        RECT 1222.230 1100.000 1222.520 1100.580 ;
        RECT 1222.380 1090.030 1222.520 1100.000 ;
        RECT 1093.520 1089.710 1093.780 1090.030 ;
        RECT 1222.320 1089.710 1222.580 1090.030 ;
        RECT 1093.580 20.730 1093.720 1089.710 ;
        RECT 1085.240 20.410 1085.500 20.730 ;
        RECT 1093.520 20.410 1093.780 20.730 ;
        RECT 1085.300 2.000 1085.440 20.410 ;
        RECT 1085.090 -4.000 1085.650 2.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1190.090 1087.560 1190.410 1087.620 ;
        RECT 1228.270 1087.560 1228.590 1087.620 ;
        RECT 1190.090 1087.420 1228.590 1087.560 ;
        RECT 1190.090 1087.360 1190.410 1087.420 ;
        RECT 1228.270 1087.360 1228.590 1087.420 ;
        RECT 1190.090 15.540 1190.410 15.600 ;
        RECT 1149.240 15.400 1190.410 15.540 ;
        RECT 1102.690 14.520 1103.010 14.580 ;
        RECT 1149.240 14.520 1149.380 15.400 ;
        RECT 1190.090 15.340 1190.410 15.400 ;
        RECT 1102.690 14.380 1149.380 14.520 ;
        RECT 1102.690 14.320 1103.010 14.380 ;
      LAYER via ;
        RECT 1190.120 1087.360 1190.380 1087.620 ;
        RECT 1228.300 1087.360 1228.560 1087.620 ;
        RECT 1102.720 14.320 1102.980 14.580 ;
        RECT 1190.120 15.340 1190.380 15.600 ;
      LAYER met2 ;
        RECT 1228.210 1100.580 1228.490 1104.000 ;
        RECT 1228.210 1100.000 1228.500 1100.580 ;
        RECT 1228.360 1087.650 1228.500 1100.000 ;
        RECT 1190.120 1087.330 1190.380 1087.650 ;
        RECT 1228.300 1087.330 1228.560 1087.650 ;
        RECT 1190.180 15.630 1190.320 1087.330 ;
        RECT 1190.120 15.310 1190.380 15.630 ;
        RECT 1102.720 14.290 1102.980 14.610 ;
        RECT 1102.780 2.000 1102.920 14.290 ;
        RECT 1102.570 -4.000 1103.130 2.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1217.690 1084.160 1218.010 1084.220 ;
        RECT 1234.710 1084.160 1235.030 1084.220 ;
        RECT 1217.690 1084.020 1235.030 1084.160 ;
        RECT 1217.690 1083.960 1218.010 1084.020 ;
        RECT 1234.710 1083.960 1235.030 1084.020 ;
        RECT 1217.690 16.220 1218.010 16.280 ;
        RECT 1144.180 16.080 1218.010 16.220 ;
        RECT 1120.630 15.540 1120.950 15.600 ;
        RECT 1144.180 15.540 1144.320 16.080 ;
        RECT 1217.690 16.020 1218.010 16.080 ;
        RECT 1120.630 15.400 1144.320 15.540 ;
        RECT 1120.630 15.340 1120.950 15.400 ;
      LAYER via ;
        RECT 1217.720 1083.960 1217.980 1084.220 ;
        RECT 1234.740 1083.960 1235.000 1084.220 ;
        RECT 1120.660 15.340 1120.920 15.600 ;
        RECT 1217.720 16.020 1217.980 16.280 ;
      LAYER met2 ;
        RECT 1234.650 1100.580 1234.930 1104.000 ;
        RECT 1234.650 1100.000 1234.940 1100.580 ;
        RECT 1234.800 1084.250 1234.940 1100.000 ;
        RECT 1217.720 1083.930 1217.980 1084.250 ;
        RECT 1234.740 1083.930 1235.000 1084.250 ;
        RECT 1217.780 16.310 1217.920 1083.930 ;
        RECT 1217.720 15.990 1217.980 16.310 ;
        RECT 1120.660 15.310 1120.920 15.630 ;
        RECT 1120.720 2.000 1120.860 15.310 ;
        RECT 1120.510 -4.000 1121.070 2.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1224.590 1083.820 1224.910 1083.880 ;
        RECT 1240.690 1083.820 1241.010 1083.880 ;
        RECT 1224.590 1083.680 1241.010 1083.820 ;
        RECT 1224.590 1083.620 1224.910 1083.680 ;
        RECT 1240.690 1083.620 1241.010 1083.680 ;
        RECT 1224.590 14.860 1224.910 14.920 ;
        RECT 1149.700 14.720 1224.910 14.860 ;
        RECT 1138.570 14.180 1138.890 14.240 ;
        RECT 1149.700 14.180 1149.840 14.720 ;
        RECT 1224.590 14.660 1224.910 14.720 ;
        RECT 1138.570 14.040 1149.840 14.180 ;
        RECT 1138.570 13.980 1138.890 14.040 ;
      LAYER via ;
        RECT 1224.620 1083.620 1224.880 1083.880 ;
        RECT 1240.720 1083.620 1240.980 1083.880 ;
        RECT 1138.600 13.980 1138.860 14.240 ;
        RECT 1224.620 14.660 1224.880 14.920 ;
      LAYER met2 ;
        RECT 1240.630 1100.580 1240.910 1104.000 ;
        RECT 1240.630 1100.000 1240.920 1100.580 ;
        RECT 1240.780 1083.910 1240.920 1100.000 ;
        RECT 1224.620 1083.590 1224.880 1083.910 ;
        RECT 1240.720 1083.590 1240.980 1083.910 ;
        RECT 1224.680 14.950 1224.820 1083.590 ;
        RECT 1224.620 14.630 1224.880 14.950 ;
        RECT 1138.600 13.950 1138.860 14.270 ;
        RECT 1138.660 2.000 1138.800 13.950 ;
        RECT 1138.450 -4.000 1139.010 2.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1156.510 15.200 1156.830 15.260 ;
        RECT 1242.990 15.200 1243.310 15.260 ;
        RECT 1156.510 15.060 1243.310 15.200 ;
        RECT 1156.510 15.000 1156.830 15.060 ;
        RECT 1242.990 15.000 1243.310 15.060 ;
      LAYER via ;
        RECT 1156.540 15.000 1156.800 15.260 ;
        RECT 1243.020 15.000 1243.280 15.260 ;
      LAYER met2 ;
        RECT 1246.610 1100.650 1246.890 1104.000 ;
        RECT 1245.380 1100.510 1246.890 1100.650 ;
        RECT 1245.380 1072.770 1245.520 1100.510 ;
        RECT 1246.610 1100.000 1246.890 1100.510 ;
        RECT 1243.080 1072.630 1245.520 1072.770 ;
        RECT 1243.080 15.290 1243.220 1072.630 ;
        RECT 1156.540 14.970 1156.800 15.290 ;
        RECT 1243.020 14.970 1243.280 15.290 ;
        RECT 1156.600 2.000 1156.740 14.970 ;
        RECT 1156.390 -4.000 1156.950 2.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1076.930 1052.200 1077.250 1052.260 ;
        RECT 1080.150 1052.200 1080.470 1052.260 ;
        RECT 1076.930 1052.060 1080.470 1052.200 ;
        RECT 1076.930 1052.000 1077.250 1052.060 ;
        RECT 1080.150 1052.000 1080.470 1052.060 ;
        RECT 674.430 47.500 674.750 47.560 ;
        RECT 1076.930 47.500 1077.250 47.560 ;
        RECT 674.430 47.360 1077.250 47.500 ;
        RECT 674.430 47.300 674.750 47.360 ;
        RECT 1076.930 47.300 1077.250 47.360 ;
      LAYER via ;
        RECT 1076.960 1052.000 1077.220 1052.260 ;
        RECT 1080.180 1052.000 1080.440 1052.260 ;
        RECT 674.460 47.300 674.720 47.560 ;
        RECT 1076.960 47.300 1077.220 47.560 ;
      LAYER met2 ;
        RECT 1081.470 1100.650 1081.750 1104.000 ;
        RECT 1080.240 1100.510 1081.750 1100.650 ;
        RECT 1080.240 1052.290 1080.380 1100.510 ;
        RECT 1081.470 1100.000 1081.750 1100.510 ;
        RECT 1076.960 1051.970 1077.220 1052.290 ;
        RECT 1080.180 1051.970 1080.440 1052.290 ;
        RECT 1077.020 47.590 1077.160 1051.970 ;
        RECT 674.460 47.270 674.720 47.590 ;
        RECT 1076.960 47.270 1077.220 47.590 ;
        RECT 674.520 2.000 674.660 47.270 ;
        RECT 674.310 -4.000 674.870 2.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1238.850 1088.240 1239.170 1088.300 ;
        RECT 1253.110 1088.240 1253.430 1088.300 ;
        RECT 1238.850 1088.100 1253.430 1088.240 ;
        RECT 1238.850 1088.040 1239.170 1088.100 ;
        RECT 1253.110 1088.040 1253.430 1088.100 ;
        RECT 1173.990 19.960 1174.310 20.020 ;
        RECT 1238.850 19.960 1239.170 20.020 ;
        RECT 1173.990 19.820 1239.170 19.960 ;
        RECT 1173.990 19.760 1174.310 19.820 ;
        RECT 1238.850 19.760 1239.170 19.820 ;
      LAYER via ;
        RECT 1238.880 1088.040 1239.140 1088.300 ;
        RECT 1253.140 1088.040 1253.400 1088.300 ;
        RECT 1174.020 19.760 1174.280 20.020 ;
        RECT 1238.880 19.760 1239.140 20.020 ;
      LAYER met2 ;
        RECT 1253.050 1100.580 1253.330 1104.000 ;
        RECT 1253.050 1100.000 1253.340 1100.580 ;
        RECT 1253.200 1088.330 1253.340 1100.000 ;
        RECT 1238.880 1088.010 1239.140 1088.330 ;
        RECT 1253.140 1088.010 1253.400 1088.330 ;
        RECT 1238.940 20.050 1239.080 1088.010 ;
        RECT 1174.020 19.730 1174.280 20.050 ;
        RECT 1238.880 19.730 1239.140 20.050 ;
        RECT 1174.080 2.000 1174.220 19.730 ;
        RECT 1173.870 -4.000 1174.430 2.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1193.310 1087.220 1193.630 1087.280 ;
        RECT 1259.090 1087.220 1259.410 1087.280 ;
        RECT 1193.310 1087.080 1259.410 1087.220 ;
        RECT 1193.310 1087.020 1193.630 1087.080 ;
        RECT 1259.090 1087.020 1259.410 1087.080 ;
      LAYER via ;
        RECT 1193.340 1087.020 1193.600 1087.280 ;
        RECT 1259.120 1087.020 1259.380 1087.280 ;
      LAYER met2 ;
        RECT 1259.030 1100.580 1259.310 1104.000 ;
        RECT 1259.030 1100.000 1259.320 1100.580 ;
        RECT 1259.180 1087.310 1259.320 1100.000 ;
        RECT 1193.340 1086.990 1193.600 1087.310 ;
        RECT 1259.120 1086.990 1259.380 1087.310 ;
        RECT 1193.400 2.450 1193.540 1086.990 ;
        RECT 1192.020 2.310 1193.540 2.450 ;
        RECT 1192.020 2.000 1192.160 2.310 ;
        RECT 1191.810 -4.000 1192.370 2.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1246.670 1085.180 1246.990 1085.240 ;
        RECT 1265.070 1085.180 1265.390 1085.240 ;
        RECT 1246.670 1085.040 1265.390 1085.180 ;
        RECT 1246.670 1084.980 1246.990 1085.040 ;
        RECT 1265.070 1084.980 1265.390 1085.040 ;
        RECT 1209.870 19.620 1210.190 19.680 ;
        RECT 1245.750 19.620 1246.070 19.680 ;
        RECT 1209.870 19.480 1246.070 19.620 ;
        RECT 1209.870 19.420 1210.190 19.480 ;
        RECT 1245.750 19.420 1246.070 19.480 ;
      LAYER via ;
        RECT 1246.700 1084.980 1246.960 1085.240 ;
        RECT 1265.100 1084.980 1265.360 1085.240 ;
        RECT 1209.900 19.420 1210.160 19.680 ;
        RECT 1245.780 19.420 1246.040 19.680 ;
      LAYER met2 ;
        RECT 1265.010 1100.580 1265.290 1104.000 ;
        RECT 1265.010 1100.000 1265.300 1100.580 ;
        RECT 1265.160 1085.270 1265.300 1100.000 ;
        RECT 1246.700 1084.950 1246.960 1085.270 ;
        RECT 1265.100 1084.950 1265.360 1085.270 ;
        RECT 1246.760 1071.410 1246.900 1084.950 ;
        RECT 1245.840 1071.270 1246.900 1071.410 ;
        RECT 1245.840 19.710 1245.980 1071.270 ;
        RECT 1209.900 19.390 1210.160 19.710 ;
        RECT 1245.780 19.390 1246.040 19.710 ;
        RECT 1209.960 2.000 1210.100 19.390 ;
        RECT 1209.750 -4.000 1210.310 2.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1254.490 1084.160 1254.810 1084.220 ;
        RECT 1271.050 1084.160 1271.370 1084.220 ;
        RECT 1254.490 1084.020 1271.370 1084.160 ;
        RECT 1254.490 1083.960 1254.810 1084.020 ;
        RECT 1271.050 1083.960 1271.370 1084.020 ;
        RECT 1227.810 16.900 1228.130 16.960 ;
        RECT 1252.650 16.900 1252.970 16.960 ;
        RECT 1227.810 16.760 1252.970 16.900 ;
        RECT 1227.810 16.700 1228.130 16.760 ;
        RECT 1252.650 16.700 1252.970 16.760 ;
      LAYER via ;
        RECT 1254.520 1083.960 1254.780 1084.220 ;
        RECT 1271.080 1083.960 1271.340 1084.220 ;
        RECT 1227.840 16.700 1228.100 16.960 ;
        RECT 1252.680 16.700 1252.940 16.960 ;
      LAYER met2 ;
        RECT 1270.990 1100.580 1271.270 1104.000 ;
        RECT 1270.990 1100.000 1271.280 1100.580 ;
        RECT 1271.140 1084.250 1271.280 1100.000 ;
        RECT 1254.520 1083.930 1254.780 1084.250 ;
        RECT 1271.080 1083.930 1271.340 1084.250 ;
        RECT 1254.580 1071.410 1254.720 1083.930 ;
        RECT 1252.740 1071.270 1254.720 1071.410 ;
        RECT 1252.740 16.990 1252.880 1071.270 ;
        RECT 1227.840 16.670 1228.100 16.990 ;
        RECT 1252.680 16.670 1252.940 16.990 ;
        RECT 1227.900 2.000 1228.040 16.670 ;
        RECT 1227.690 -4.000 1228.250 2.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1259.550 1084.500 1259.870 1084.560 ;
        RECT 1277.490 1084.500 1277.810 1084.560 ;
        RECT 1259.550 1084.360 1277.810 1084.500 ;
        RECT 1259.550 1084.300 1259.870 1084.360 ;
        RECT 1277.490 1084.300 1277.810 1084.360 ;
        RECT 1245.750 17.240 1246.070 17.300 ;
        RECT 1259.550 17.240 1259.870 17.300 ;
        RECT 1245.750 17.100 1259.870 17.240 ;
        RECT 1245.750 17.040 1246.070 17.100 ;
        RECT 1259.550 17.040 1259.870 17.100 ;
      LAYER via ;
        RECT 1259.580 1084.300 1259.840 1084.560 ;
        RECT 1277.520 1084.300 1277.780 1084.560 ;
        RECT 1245.780 17.040 1246.040 17.300 ;
        RECT 1259.580 17.040 1259.840 17.300 ;
      LAYER met2 ;
        RECT 1277.430 1100.580 1277.710 1104.000 ;
        RECT 1277.430 1100.000 1277.720 1100.580 ;
        RECT 1277.580 1084.590 1277.720 1100.000 ;
        RECT 1259.580 1084.270 1259.840 1084.590 ;
        RECT 1277.520 1084.270 1277.780 1084.590 ;
        RECT 1259.640 17.330 1259.780 1084.270 ;
        RECT 1245.780 17.010 1246.040 17.330 ;
        RECT 1259.580 17.010 1259.840 17.330 ;
        RECT 1245.840 2.000 1245.980 17.010 ;
        RECT 1245.630 -4.000 1246.190 2.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1272.890 1084.160 1273.210 1084.220 ;
        RECT 1283.470 1084.160 1283.790 1084.220 ;
        RECT 1272.890 1084.020 1283.790 1084.160 ;
        RECT 1272.890 1083.960 1273.210 1084.020 ;
        RECT 1283.470 1083.960 1283.790 1084.020 ;
        RECT 1263.230 15.200 1263.550 15.260 ;
        RECT 1272.890 15.200 1273.210 15.260 ;
        RECT 1263.230 15.060 1273.210 15.200 ;
        RECT 1263.230 15.000 1263.550 15.060 ;
        RECT 1272.890 15.000 1273.210 15.060 ;
      LAYER via ;
        RECT 1272.920 1083.960 1273.180 1084.220 ;
        RECT 1283.500 1083.960 1283.760 1084.220 ;
        RECT 1263.260 15.000 1263.520 15.260 ;
        RECT 1272.920 15.000 1273.180 15.260 ;
      LAYER met2 ;
        RECT 1283.410 1100.580 1283.690 1104.000 ;
        RECT 1283.410 1100.000 1283.700 1100.580 ;
        RECT 1283.560 1084.250 1283.700 1100.000 ;
        RECT 1272.920 1083.930 1273.180 1084.250 ;
        RECT 1283.500 1083.930 1283.760 1084.250 ;
        RECT 1272.980 15.290 1273.120 1083.930 ;
        RECT 1263.260 14.970 1263.520 15.290 ;
        RECT 1272.920 14.970 1273.180 15.290 ;
        RECT 1263.320 2.000 1263.460 14.970 ;
        RECT 1263.110 -4.000 1263.670 2.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1283.010 1088.580 1283.330 1088.640 ;
        RECT 1289.450 1088.580 1289.770 1088.640 ;
        RECT 1283.010 1088.440 1289.770 1088.580 ;
        RECT 1283.010 1088.380 1283.330 1088.440 ;
        RECT 1289.450 1088.380 1289.770 1088.440 ;
      LAYER via ;
        RECT 1283.040 1088.380 1283.300 1088.640 ;
        RECT 1289.480 1088.380 1289.740 1088.640 ;
      LAYER met2 ;
        RECT 1289.390 1100.580 1289.670 1104.000 ;
        RECT 1289.390 1100.000 1289.680 1100.580 ;
        RECT 1289.540 1088.670 1289.680 1100.000 ;
        RECT 1283.040 1088.350 1283.300 1088.670 ;
        RECT 1289.480 1088.350 1289.740 1088.670 ;
        RECT 1283.100 2.450 1283.240 1088.350 ;
        RECT 1281.260 2.310 1283.240 2.450 ;
        RECT 1281.260 2.000 1281.400 2.310 ;
        RECT 1281.050 -4.000 1281.610 2.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1296.810 20.640 1297.130 20.700 ;
        RECT 1299.110 20.640 1299.430 20.700 ;
        RECT 1296.810 20.500 1299.430 20.640 ;
        RECT 1296.810 20.440 1297.130 20.500 ;
        RECT 1299.110 20.440 1299.430 20.500 ;
      LAYER via ;
        RECT 1296.840 20.440 1297.100 20.700 ;
        RECT 1299.140 20.440 1299.400 20.700 ;
      LAYER met2 ;
        RECT 1295.830 1100.650 1296.110 1104.000 ;
        RECT 1295.830 1100.510 1297.040 1100.650 ;
        RECT 1295.830 1100.000 1296.110 1100.510 ;
        RECT 1296.900 20.730 1297.040 1100.510 ;
        RECT 1296.840 20.410 1297.100 20.730 ;
        RECT 1299.140 20.410 1299.400 20.730 ;
        RECT 1299.200 2.000 1299.340 20.410 ;
        RECT 1298.990 -4.000 1299.550 2.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1312.985 1027.905 1313.155 1055.615 ;
        RECT 1312.525 931.345 1312.695 959.055 ;
        RECT 1312.985 862.665 1313.155 910.435 ;
        RECT 1311.605 386.325 1311.775 434.775 ;
        RECT 1312.525 241.485 1312.695 289.595 ;
      LAYER mcon ;
        RECT 1312.985 1055.445 1313.155 1055.615 ;
        RECT 1312.525 958.885 1312.695 959.055 ;
        RECT 1312.985 910.265 1313.155 910.435 ;
        RECT 1311.605 434.605 1311.775 434.775 ;
        RECT 1312.525 289.425 1312.695 289.595 ;
      LAYER met1 ;
        RECT 1301.870 1056.280 1302.190 1056.340 ;
        RECT 1312.910 1056.280 1313.230 1056.340 ;
        RECT 1301.870 1056.140 1313.230 1056.280 ;
        RECT 1301.870 1056.080 1302.190 1056.140 ;
        RECT 1312.910 1056.080 1313.230 1056.140 ;
        RECT 1312.910 1055.600 1313.230 1055.660 ;
        RECT 1312.715 1055.460 1313.230 1055.600 ;
        RECT 1312.910 1055.400 1313.230 1055.460 ;
        RECT 1312.910 1028.060 1313.230 1028.120 ;
        RECT 1312.715 1027.920 1313.230 1028.060 ;
        RECT 1312.910 1027.860 1313.230 1027.920 ;
        RECT 1311.990 983.180 1312.310 983.240 ;
        RECT 1313.370 983.180 1313.690 983.240 ;
        RECT 1311.990 983.040 1313.690 983.180 ;
        RECT 1311.990 982.980 1312.310 983.040 ;
        RECT 1313.370 982.980 1313.690 983.040 ;
        RECT 1312.450 959.040 1312.770 959.100 ;
        RECT 1312.255 958.900 1312.770 959.040 ;
        RECT 1312.450 958.840 1312.770 958.900 ;
        RECT 1312.450 931.500 1312.770 931.560 ;
        RECT 1312.255 931.360 1312.770 931.500 ;
        RECT 1312.450 931.300 1312.770 931.360 ;
        RECT 1312.910 910.420 1313.230 910.480 ;
        RECT 1312.715 910.280 1313.230 910.420 ;
        RECT 1312.910 910.220 1313.230 910.280 ;
        RECT 1312.910 862.820 1313.230 862.880 ;
        RECT 1312.715 862.680 1313.230 862.820 ;
        RECT 1312.910 862.620 1313.230 862.680 ;
        RECT 1311.530 821.000 1311.850 821.060 ;
        RECT 1312.450 821.000 1312.770 821.060 ;
        RECT 1311.530 820.860 1312.770 821.000 ;
        RECT 1311.530 820.800 1311.850 820.860 ;
        RECT 1312.450 820.800 1312.770 820.860 ;
        RECT 1311.545 434.760 1311.835 434.805 ;
        RECT 1311.990 434.760 1312.310 434.820 ;
        RECT 1311.545 434.620 1312.310 434.760 ;
        RECT 1311.545 434.575 1311.835 434.620 ;
        RECT 1311.990 434.560 1312.310 434.620 ;
        RECT 1311.530 386.480 1311.850 386.540 ;
        RECT 1311.335 386.340 1311.850 386.480 ;
        RECT 1311.530 386.280 1311.850 386.340 ;
        RECT 1311.990 303.520 1312.310 303.580 ;
        RECT 1312.910 303.520 1313.230 303.580 ;
        RECT 1311.990 303.380 1313.230 303.520 ;
        RECT 1311.990 303.320 1312.310 303.380 ;
        RECT 1312.910 303.320 1313.230 303.380 ;
        RECT 1312.465 289.580 1312.755 289.625 ;
        RECT 1312.910 289.580 1313.230 289.640 ;
        RECT 1312.465 289.440 1313.230 289.580 ;
        RECT 1312.465 289.395 1312.755 289.440 ;
        RECT 1312.910 289.380 1313.230 289.440 ;
        RECT 1312.450 241.640 1312.770 241.700 ;
        RECT 1312.255 241.500 1312.770 241.640 ;
        RECT 1312.450 241.440 1312.770 241.500 ;
        RECT 1311.990 206.960 1312.310 207.020 ;
        RECT 1312.910 206.960 1313.230 207.020 ;
        RECT 1311.990 206.820 1313.230 206.960 ;
        RECT 1311.990 206.760 1312.310 206.820 ;
        RECT 1312.910 206.760 1313.230 206.820 ;
        RECT 1311.990 110.400 1312.310 110.460 ;
        RECT 1312.910 110.400 1313.230 110.460 ;
        RECT 1311.990 110.260 1313.230 110.400 ;
        RECT 1311.990 110.200 1312.310 110.260 ;
        RECT 1312.910 110.200 1313.230 110.260 ;
      LAYER via ;
        RECT 1301.900 1056.080 1302.160 1056.340 ;
        RECT 1312.940 1056.080 1313.200 1056.340 ;
        RECT 1312.940 1055.400 1313.200 1055.660 ;
        RECT 1312.940 1027.860 1313.200 1028.120 ;
        RECT 1312.020 982.980 1312.280 983.240 ;
        RECT 1313.400 982.980 1313.660 983.240 ;
        RECT 1312.480 958.840 1312.740 959.100 ;
        RECT 1312.480 931.300 1312.740 931.560 ;
        RECT 1312.940 910.220 1313.200 910.480 ;
        RECT 1312.940 862.620 1313.200 862.880 ;
        RECT 1311.560 820.800 1311.820 821.060 ;
        RECT 1312.480 820.800 1312.740 821.060 ;
        RECT 1312.020 434.560 1312.280 434.820 ;
        RECT 1311.560 386.280 1311.820 386.540 ;
        RECT 1312.020 303.320 1312.280 303.580 ;
        RECT 1312.940 303.320 1313.200 303.580 ;
        RECT 1312.940 289.380 1313.200 289.640 ;
        RECT 1312.480 241.440 1312.740 241.700 ;
        RECT 1312.020 206.760 1312.280 207.020 ;
        RECT 1312.940 206.760 1313.200 207.020 ;
        RECT 1312.020 110.200 1312.280 110.460 ;
        RECT 1312.940 110.200 1313.200 110.460 ;
      LAYER met2 ;
        RECT 1301.810 1100.580 1302.090 1104.000 ;
        RECT 1301.810 1100.000 1302.100 1100.580 ;
        RECT 1301.960 1056.370 1302.100 1100.000 ;
        RECT 1301.900 1056.050 1302.160 1056.370 ;
        RECT 1312.940 1056.050 1313.200 1056.370 ;
        RECT 1313.000 1055.690 1313.140 1056.050 ;
        RECT 1312.940 1055.370 1313.200 1055.690 ;
        RECT 1312.940 1027.830 1313.200 1028.150 ;
        RECT 1313.000 1007.490 1313.140 1027.830 ;
        RECT 1313.000 1007.350 1313.600 1007.490 ;
        RECT 1313.460 983.270 1313.600 1007.350 ;
        RECT 1312.020 982.950 1312.280 983.270 ;
        RECT 1313.400 982.950 1313.660 983.270 ;
        RECT 1312.080 959.210 1312.220 982.950 ;
        RECT 1312.080 959.130 1312.680 959.210 ;
        RECT 1312.080 959.070 1312.740 959.130 ;
        RECT 1312.480 958.810 1312.740 959.070 ;
        RECT 1312.540 958.655 1312.680 958.810 ;
        RECT 1312.480 931.270 1312.740 931.590 ;
        RECT 1312.540 910.930 1312.680 931.270 ;
        RECT 1312.540 910.790 1313.140 910.930 ;
        RECT 1313.000 910.510 1313.140 910.790 ;
        RECT 1312.940 910.190 1313.200 910.510 ;
        RECT 1312.940 862.590 1313.200 862.910 ;
        RECT 1313.000 834.770 1313.140 862.590 ;
        RECT 1312.540 834.630 1313.140 834.770 ;
        RECT 1312.540 821.090 1312.680 834.630 ;
        RECT 1311.560 820.770 1311.820 821.090 ;
        RECT 1312.480 820.770 1312.740 821.090 ;
        RECT 1311.620 773.005 1311.760 820.770 ;
        RECT 1311.550 772.635 1311.830 773.005 ;
        RECT 1312.930 772.635 1313.210 773.005 ;
        RECT 1313.000 738.210 1313.140 772.635 ;
        RECT 1312.540 738.070 1313.140 738.210 ;
        RECT 1312.540 700.130 1312.680 738.070 ;
        RECT 1311.620 699.990 1312.680 700.130 ;
        RECT 1311.620 676.445 1311.760 699.990 ;
        RECT 1311.550 676.075 1311.830 676.445 ;
        RECT 1312.930 676.075 1313.210 676.445 ;
        RECT 1313.000 641.650 1313.140 676.075 ;
        RECT 1312.540 641.510 1313.140 641.650 ;
        RECT 1312.540 603.570 1312.680 641.510 ;
        RECT 1311.620 603.430 1312.680 603.570 ;
        RECT 1311.620 579.885 1311.760 603.430 ;
        RECT 1311.550 579.515 1311.830 579.885 ;
        RECT 1312.930 579.515 1313.210 579.885 ;
        RECT 1313.000 545.090 1313.140 579.515 ;
        RECT 1312.540 544.950 1313.140 545.090 ;
        RECT 1312.540 507.010 1312.680 544.950 ;
        RECT 1311.620 506.870 1312.680 507.010 ;
        RECT 1311.620 483.325 1311.760 506.870 ;
        RECT 1311.550 482.955 1311.830 483.325 ;
        RECT 1312.930 482.955 1313.210 483.325 ;
        RECT 1313.000 448.530 1313.140 482.955 ;
        RECT 1312.080 448.390 1313.140 448.530 ;
        RECT 1312.080 434.850 1312.220 448.390 ;
        RECT 1312.020 434.530 1312.280 434.850 ;
        RECT 1311.560 386.250 1311.820 386.570 ;
        RECT 1311.620 351.290 1311.760 386.250 ;
        RECT 1311.620 351.150 1312.220 351.290 ;
        RECT 1312.080 303.610 1312.220 351.150 ;
        RECT 1312.020 303.290 1312.280 303.610 ;
        RECT 1312.940 303.290 1313.200 303.610 ;
        RECT 1313.000 289.670 1313.140 303.290 ;
        RECT 1312.940 289.350 1313.200 289.670 ;
        RECT 1312.480 241.410 1312.740 241.730 ;
        RECT 1312.540 207.130 1312.680 241.410 ;
        RECT 1312.080 207.050 1312.680 207.130 ;
        RECT 1312.020 206.990 1312.680 207.050 ;
        RECT 1312.020 206.730 1312.280 206.990 ;
        RECT 1312.940 206.730 1313.200 207.050 ;
        RECT 1313.000 158.850 1313.140 206.730 ;
        RECT 1312.540 158.710 1313.140 158.850 ;
        RECT 1312.540 110.570 1312.680 158.710 ;
        RECT 1312.080 110.490 1312.680 110.570 ;
        RECT 1312.020 110.430 1312.680 110.490 ;
        RECT 1312.020 110.170 1312.280 110.430 ;
        RECT 1312.940 110.170 1313.200 110.490 ;
        RECT 1313.000 16.730 1313.140 110.170 ;
        RECT 1313.000 16.590 1317.280 16.730 ;
        RECT 1317.140 2.000 1317.280 16.590 ;
        RECT 1316.930 -4.000 1317.490 2.000 ;
      LAYER via2 ;
        RECT 1311.550 772.680 1311.830 772.960 ;
        RECT 1312.930 772.680 1313.210 772.960 ;
        RECT 1311.550 676.120 1311.830 676.400 ;
        RECT 1312.930 676.120 1313.210 676.400 ;
        RECT 1311.550 579.560 1311.830 579.840 ;
        RECT 1312.930 579.560 1313.210 579.840 ;
        RECT 1311.550 483.000 1311.830 483.280 ;
        RECT 1312.930 483.000 1313.210 483.280 ;
      LAYER met3 ;
        RECT 1311.525 772.970 1311.855 772.985 ;
        RECT 1312.905 772.970 1313.235 772.985 ;
        RECT 1311.525 772.670 1313.235 772.970 ;
        RECT 1311.525 772.655 1311.855 772.670 ;
        RECT 1312.905 772.655 1313.235 772.670 ;
        RECT 1311.525 676.410 1311.855 676.425 ;
        RECT 1312.905 676.410 1313.235 676.425 ;
        RECT 1311.525 676.110 1313.235 676.410 ;
        RECT 1311.525 676.095 1311.855 676.110 ;
        RECT 1312.905 676.095 1313.235 676.110 ;
        RECT 1311.525 579.850 1311.855 579.865 ;
        RECT 1312.905 579.850 1313.235 579.865 ;
        RECT 1311.525 579.550 1313.235 579.850 ;
        RECT 1311.525 579.535 1311.855 579.550 ;
        RECT 1312.905 579.535 1313.235 579.550 ;
        RECT 1311.525 483.290 1311.855 483.305 ;
        RECT 1312.905 483.290 1313.235 483.305 ;
        RECT 1311.525 482.990 1313.235 483.290 ;
        RECT 1311.525 482.975 1311.855 482.990 ;
        RECT 1312.905 482.975 1313.235 482.990 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1309.690 1059.680 1310.010 1059.740 ;
        RECT 1332.690 1059.680 1333.010 1059.740 ;
        RECT 1309.690 1059.540 1333.010 1059.680 ;
        RECT 1309.690 1059.480 1310.010 1059.540 ;
        RECT 1332.690 1059.480 1333.010 1059.540 ;
        RECT 1332.690 1055.600 1333.010 1055.660 ;
        RECT 1333.610 1055.600 1333.930 1055.660 ;
        RECT 1332.690 1055.460 1333.930 1055.600 ;
        RECT 1332.690 1055.400 1333.010 1055.460 ;
        RECT 1333.610 1055.400 1333.930 1055.460 ;
        RECT 1332.690 159.160 1333.010 159.420 ;
        RECT 1332.780 158.740 1332.920 159.160 ;
        RECT 1332.690 158.480 1333.010 158.740 ;
        RECT 1332.690 118.220 1333.010 118.280 ;
        RECT 1334.070 118.220 1334.390 118.280 ;
        RECT 1332.690 118.080 1334.390 118.220 ;
        RECT 1332.690 118.020 1333.010 118.080 ;
        RECT 1334.070 118.020 1334.390 118.080 ;
      LAYER via ;
        RECT 1309.720 1059.480 1309.980 1059.740 ;
        RECT 1332.720 1059.480 1332.980 1059.740 ;
        RECT 1332.720 1055.400 1332.980 1055.660 ;
        RECT 1333.640 1055.400 1333.900 1055.660 ;
        RECT 1332.720 159.160 1332.980 159.420 ;
        RECT 1332.720 158.480 1332.980 158.740 ;
        RECT 1332.720 118.020 1332.980 118.280 ;
        RECT 1334.100 118.020 1334.360 118.280 ;
      LAYER met2 ;
        RECT 1307.790 1100.650 1308.070 1104.000 ;
        RECT 1307.790 1100.510 1309.920 1100.650 ;
        RECT 1307.790 1100.000 1308.070 1100.510 ;
        RECT 1309.780 1059.770 1309.920 1100.510 ;
        RECT 1309.720 1059.450 1309.980 1059.770 ;
        RECT 1332.720 1059.450 1332.980 1059.770 ;
        RECT 1332.780 1055.690 1332.920 1059.450 ;
        RECT 1332.720 1055.370 1332.980 1055.690 ;
        RECT 1333.640 1055.370 1333.900 1055.690 ;
        RECT 1333.700 959.325 1333.840 1055.370 ;
        RECT 1332.710 958.955 1332.990 959.325 ;
        RECT 1333.630 958.955 1333.910 959.325 ;
        RECT 1332.780 835.450 1332.920 958.955 ;
        RECT 1332.320 835.310 1332.920 835.450 ;
        RECT 1332.320 834.770 1332.460 835.310 ;
        RECT 1332.320 834.630 1332.920 834.770 ;
        RECT 1332.780 738.890 1332.920 834.630 ;
        RECT 1332.320 738.750 1332.920 738.890 ;
        RECT 1332.320 738.210 1332.460 738.750 ;
        RECT 1332.320 738.070 1332.920 738.210 ;
        RECT 1332.780 642.330 1332.920 738.070 ;
        RECT 1332.320 642.190 1332.920 642.330 ;
        RECT 1332.320 641.650 1332.460 642.190 ;
        RECT 1332.320 641.510 1332.920 641.650 ;
        RECT 1332.780 545.770 1332.920 641.510 ;
        RECT 1332.320 545.630 1332.920 545.770 ;
        RECT 1332.320 545.090 1332.460 545.630 ;
        RECT 1332.320 544.950 1332.920 545.090 ;
        RECT 1332.780 449.210 1332.920 544.950 ;
        RECT 1332.320 449.070 1332.920 449.210 ;
        RECT 1332.320 448.530 1332.460 449.070 ;
        RECT 1332.320 448.390 1332.920 448.530 ;
        RECT 1332.780 351.970 1332.920 448.390 ;
        RECT 1332.320 351.830 1332.920 351.970 ;
        RECT 1332.320 351.290 1332.460 351.830 ;
        RECT 1332.320 351.150 1332.920 351.290 ;
        RECT 1332.780 255.410 1332.920 351.150 ;
        RECT 1332.320 255.270 1332.920 255.410 ;
        RECT 1332.320 254.730 1332.460 255.270 ;
        RECT 1332.320 254.590 1332.920 254.730 ;
        RECT 1332.780 159.450 1332.920 254.590 ;
        RECT 1332.720 159.130 1332.980 159.450 ;
        RECT 1332.720 158.450 1332.980 158.770 ;
        RECT 1332.780 118.310 1332.920 158.450 ;
        RECT 1332.720 117.990 1332.980 118.310 ;
        RECT 1334.100 117.990 1334.360 118.310 ;
        RECT 1334.160 96.290 1334.300 117.990 ;
        RECT 1334.160 96.150 1334.760 96.290 ;
        RECT 1334.620 16.050 1334.760 96.150 ;
        RECT 1334.620 15.910 1335.220 16.050 ;
        RECT 1335.080 2.000 1335.220 15.910 ;
        RECT 1334.870 -4.000 1335.430 2.000 ;
      LAYER via2 ;
        RECT 1332.710 959.000 1332.990 959.280 ;
        RECT 1333.630 959.000 1333.910 959.280 ;
      LAYER met3 ;
        RECT 1332.685 959.290 1333.015 959.305 ;
        RECT 1333.605 959.290 1333.935 959.305 ;
        RECT 1332.685 958.990 1333.935 959.290 ;
        RECT 1332.685 958.975 1333.015 958.990 ;
        RECT 1333.605 958.975 1333.935 958.990 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1084.290 1078.040 1084.610 1078.100 ;
        RECT 1087.510 1078.040 1087.830 1078.100 ;
        RECT 1084.290 1077.900 1087.830 1078.040 ;
        RECT 1084.290 1077.840 1084.610 1077.900 ;
        RECT 1087.510 1077.840 1087.830 1077.900 ;
        RECT 692.370 48.180 692.690 48.240 ;
        RECT 692.370 48.040 1084.520 48.180 ;
        RECT 692.370 47.980 692.690 48.040 ;
        RECT 1084.380 47.900 1084.520 48.040 ;
        RECT 1084.290 47.640 1084.610 47.900 ;
      LAYER via ;
        RECT 1084.320 1077.840 1084.580 1078.100 ;
        RECT 1087.540 1077.840 1087.800 1078.100 ;
        RECT 692.400 47.980 692.660 48.240 ;
        RECT 1084.320 47.640 1084.580 47.900 ;
      LAYER met2 ;
        RECT 1087.450 1100.580 1087.730 1104.000 ;
        RECT 1087.450 1100.000 1087.740 1100.580 ;
        RECT 1087.600 1078.130 1087.740 1100.000 ;
        RECT 1084.320 1077.810 1084.580 1078.130 ;
        RECT 1087.540 1077.810 1087.800 1078.130 ;
        RECT 692.400 47.950 692.660 48.270 ;
        RECT 692.460 2.000 692.600 47.950 ;
        RECT 1084.380 47.930 1084.520 1077.810 ;
        RECT 1084.320 47.610 1084.580 47.930 ;
        RECT 692.250 -4.000 692.810 2.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1314.290 1088.580 1314.610 1088.640 ;
        RECT 1317.510 1088.580 1317.830 1088.640 ;
        RECT 1314.290 1088.440 1317.830 1088.580 ;
        RECT 1314.290 1088.380 1314.610 1088.440 ;
        RECT 1317.510 1088.380 1317.830 1088.440 ;
        RECT 1317.510 20.300 1317.830 20.360 ;
        RECT 1352.470 20.300 1352.790 20.360 ;
        RECT 1317.510 20.160 1352.790 20.300 ;
        RECT 1317.510 20.100 1317.830 20.160 ;
        RECT 1352.470 20.100 1352.790 20.160 ;
      LAYER via ;
        RECT 1314.320 1088.380 1314.580 1088.640 ;
        RECT 1317.540 1088.380 1317.800 1088.640 ;
        RECT 1317.540 20.100 1317.800 20.360 ;
        RECT 1352.500 20.100 1352.760 20.360 ;
      LAYER met2 ;
        RECT 1314.230 1100.580 1314.510 1104.000 ;
        RECT 1314.230 1100.000 1314.520 1100.580 ;
        RECT 1314.380 1088.670 1314.520 1100.000 ;
        RECT 1314.320 1088.350 1314.580 1088.670 ;
        RECT 1317.540 1088.350 1317.800 1088.670 ;
        RECT 1317.600 20.390 1317.740 1088.350 ;
        RECT 1317.540 20.070 1317.800 20.390 ;
        RECT 1352.500 20.070 1352.760 20.390 ;
        RECT 1352.560 2.000 1352.700 20.070 ;
        RECT 1352.350 -4.000 1352.910 2.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1320.270 1086.880 1320.590 1086.940 ;
        RECT 1334.990 1086.880 1335.310 1086.940 ;
        RECT 1320.270 1086.740 1335.310 1086.880 ;
        RECT 1320.270 1086.680 1320.590 1086.740 ;
        RECT 1334.990 1086.680 1335.310 1086.740 ;
        RECT 1334.990 16.900 1335.310 16.960 ;
        RECT 1370.410 16.900 1370.730 16.960 ;
        RECT 1334.990 16.760 1370.730 16.900 ;
        RECT 1334.990 16.700 1335.310 16.760 ;
        RECT 1370.410 16.700 1370.730 16.760 ;
      LAYER via ;
        RECT 1320.300 1086.680 1320.560 1086.940 ;
        RECT 1335.020 1086.680 1335.280 1086.940 ;
        RECT 1335.020 16.700 1335.280 16.960 ;
        RECT 1370.440 16.700 1370.700 16.960 ;
      LAYER met2 ;
        RECT 1320.210 1100.580 1320.490 1104.000 ;
        RECT 1320.210 1100.000 1320.500 1100.580 ;
        RECT 1320.360 1086.970 1320.500 1100.000 ;
        RECT 1320.300 1086.650 1320.560 1086.970 ;
        RECT 1335.020 1086.650 1335.280 1086.970 ;
        RECT 1335.080 16.990 1335.220 1086.650 ;
        RECT 1335.020 16.670 1335.280 16.990 ;
        RECT 1370.440 16.670 1370.700 16.990 ;
        RECT 1370.500 2.000 1370.640 16.670 ;
        RECT 1370.290 -4.000 1370.850 2.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1326.250 1086.540 1326.570 1086.600 ;
        RECT 1383.290 1086.540 1383.610 1086.600 ;
        RECT 1326.250 1086.400 1383.610 1086.540 ;
        RECT 1326.250 1086.340 1326.570 1086.400 ;
        RECT 1383.290 1086.340 1383.610 1086.400 ;
        RECT 1383.290 20.640 1383.610 20.700 ;
        RECT 1388.350 20.640 1388.670 20.700 ;
        RECT 1383.290 20.500 1388.670 20.640 ;
        RECT 1383.290 20.440 1383.610 20.500 ;
        RECT 1388.350 20.440 1388.670 20.500 ;
      LAYER via ;
        RECT 1326.280 1086.340 1326.540 1086.600 ;
        RECT 1383.320 1086.340 1383.580 1086.600 ;
        RECT 1383.320 20.440 1383.580 20.700 ;
        RECT 1388.380 20.440 1388.640 20.700 ;
      LAYER met2 ;
        RECT 1326.190 1100.580 1326.470 1104.000 ;
        RECT 1326.190 1100.000 1326.480 1100.580 ;
        RECT 1326.340 1086.630 1326.480 1100.000 ;
        RECT 1326.280 1086.310 1326.540 1086.630 ;
        RECT 1383.320 1086.310 1383.580 1086.630 ;
        RECT 1383.380 20.730 1383.520 1086.310 ;
        RECT 1383.320 20.410 1383.580 20.730 ;
        RECT 1388.380 20.410 1388.640 20.730 ;
        RECT 1388.440 2.000 1388.580 20.410 ;
        RECT 1388.230 -4.000 1388.790 2.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1370.945 18.105 1371.115 18.955 ;
      LAYER mcon ;
        RECT 1370.945 18.785 1371.115 18.955 ;
      LAYER met1 ;
        RECT 1332.690 1085.180 1333.010 1085.240 ;
        RECT 1338.210 1085.180 1338.530 1085.240 ;
        RECT 1332.690 1085.040 1338.530 1085.180 ;
        RECT 1332.690 1084.980 1333.010 1085.040 ;
        RECT 1338.210 1084.980 1338.530 1085.040 ;
        RECT 1338.210 18.940 1338.530 19.000 ;
        RECT 1370.885 18.940 1371.175 18.985 ;
        RECT 1338.210 18.800 1371.175 18.940 ;
        RECT 1338.210 18.740 1338.530 18.800 ;
        RECT 1370.885 18.755 1371.175 18.800 ;
        RECT 1370.885 18.260 1371.175 18.305 ;
        RECT 1406.290 18.260 1406.610 18.320 ;
        RECT 1370.885 18.120 1406.610 18.260 ;
        RECT 1370.885 18.075 1371.175 18.120 ;
        RECT 1406.290 18.060 1406.610 18.120 ;
      LAYER via ;
        RECT 1332.720 1084.980 1332.980 1085.240 ;
        RECT 1338.240 1084.980 1338.500 1085.240 ;
        RECT 1338.240 18.740 1338.500 19.000 ;
        RECT 1406.320 18.060 1406.580 18.320 ;
      LAYER met2 ;
        RECT 1332.630 1100.580 1332.910 1104.000 ;
        RECT 1332.630 1100.000 1332.920 1100.580 ;
        RECT 1332.780 1085.270 1332.920 1100.000 ;
        RECT 1332.720 1084.950 1332.980 1085.270 ;
        RECT 1338.240 1084.950 1338.500 1085.270 ;
        RECT 1338.300 19.030 1338.440 1084.950 ;
        RECT 1338.240 18.710 1338.500 19.030 ;
        RECT 1406.320 18.030 1406.580 18.350 ;
        RECT 1406.380 2.000 1406.520 18.030 ;
        RECT 1406.170 -4.000 1406.730 2.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1338.670 1088.580 1338.990 1088.640 ;
        RECT 1344.650 1088.580 1344.970 1088.640 ;
        RECT 1338.670 1088.440 1344.970 1088.580 ;
        RECT 1338.670 1088.380 1338.990 1088.440 ;
        RECT 1344.650 1088.380 1344.970 1088.440 ;
        RECT 1344.650 14.180 1344.970 14.240 ;
        RECT 1423.770 14.180 1424.090 14.240 ;
        RECT 1344.650 14.040 1424.090 14.180 ;
        RECT 1344.650 13.980 1344.970 14.040 ;
        RECT 1423.770 13.980 1424.090 14.040 ;
      LAYER via ;
        RECT 1338.700 1088.380 1338.960 1088.640 ;
        RECT 1344.680 1088.380 1344.940 1088.640 ;
        RECT 1344.680 13.980 1344.940 14.240 ;
        RECT 1423.800 13.980 1424.060 14.240 ;
      LAYER met2 ;
        RECT 1338.610 1100.580 1338.890 1104.000 ;
        RECT 1338.610 1100.000 1338.900 1100.580 ;
        RECT 1338.760 1088.670 1338.900 1100.000 ;
        RECT 1338.700 1088.350 1338.960 1088.670 ;
        RECT 1344.680 1088.350 1344.940 1088.670 ;
        RECT 1344.740 14.270 1344.880 1088.350 ;
        RECT 1344.680 13.950 1344.940 14.270 ;
        RECT 1423.800 13.950 1424.060 14.270 ;
        RECT 1423.860 2.000 1424.000 13.950 ;
        RECT 1423.650 -4.000 1424.210 2.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1345.110 14.520 1345.430 14.580 ;
        RECT 1441.710 14.520 1442.030 14.580 ;
        RECT 1345.110 14.380 1442.030 14.520 ;
        RECT 1345.110 14.320 1345.430 14.380 ;
        RECT 1441.710 14.320 1442.030 14.380 ;
      LAYER via ;
        RECT 1345.140 14.320 1345.400 14.580 ;
        RECT 1441.740 14.320 1442.000 14.580 ;
      LAYER met2 ;
        RECT 1344.590 1100.650 1344.870 1104.000 ;
        RECT 1344.590 1100.510 1345.340 1100.650 ;
        RECT 1344.590 1100.000 1344.870 1100.510 ;
        RECT 1345.200 14.610 1345.340 1100.510 ;
        RECT 1345.140 14.290 1345.400 14.610 ;
        RECT 1441.740 14.290 1442.000 14.610 ;
        RECT 1441.800 2.000 1441.940 14.290 ;
        RECT 1441.590 -4.000 1442.150 2.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1390.265 17.425 1390.435 18.615 ;
      LAYER mcon ;
        RECT 1390.265 18.445 1390.435 18.615 ;
      LAYER met1 ;
        RECT 1352.010 18.600 1352.330 18.660 ;
        RECT 1390.205 18.600 1390.495 18.645 ;
        RECT 1352.010 18.460 1390.495 18.600 ;
        RECT 1352.010 18.400 1352.330 18.460 ;
        RECT 1390.205 18.415 1390.495 18.460 ;
        RECT 1390.205 17.580 1390.495 17.625 ;
        RECT 1459.650 17.580 1459.970 17.640 ;
        RECT 1390.205 17.440 1459.970 17.580 ;
        RECT 1390.205 17.395 1390.495 17.440 ;
        RECT 1459.650 17.380 1459.970 17.440 ;
      LAYER via ;
        RECT 1352.040 18.400 1352.300 18.660 ;
        RECT 1459.680 17.380 1459.940 17.640 ;
      LAYER met2 ;
        RECT 1351.030 1100.650 1351.310 1104.000 ;
        RECT 1351.030 1100.510 1352.240 1100.650 ;
        RECT 1351.030 1100.000 1351.310 1100.510 ;
        RECT 1352.100 18.690 1352.240 1100.510 ;
        RECT 1352.040 18.370 1352.300 18.690 ;
        RECT 1459.680 17.350 1459.940 17.670 ;
        RECT 1459.740 2.000 1459.880 17.350 ;
        RECT 1459.530 -4.000 1460.090 2.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1357.070 1084.160 1357.390 1084.220 ;
        RECT 1369.490 1084.160 1369.810 1084.220 ;
        RECT 1357.070 1084.020 1369.810 1084.160 ;
        RECT 1357.070 1083.960 1357.390 1084.020 ;
        RECT 1369.490 1083.960 1369.810 1084.020 ;
        RECT 1370.870 16.900 1371.190 16.960 ;
        RECT 1370.870 16.760 1372.480 16.900 ;
        RECT 1370.870 16.700 1371.190 16.760 ;
        RECT 1372.340 16.560 1372.480 16.760 ;
        RECT 1386.050 16.560 1386.370 16.620 ;
        RECT 1372.340 16.420 1386.370 16.560 ;
        RECT 1386.050 16.360 1386.370 16.420 ;
        RECT 1402.150 15.200 1402.470 15.260 ;
        RECT 1477.590 15.200 1477.910 15.260 ;
        RECT 1402.150 15.060 1477.910 15.200 ;
        RECT 1402.150 15.000 1402.470 15.060 ;
        RECT 1477.590 15.000 1477.910 15.060 ;
      LAYER via ;
        RECT 1357.100 1083.960 1357.360 1084.220 ;
        RECT 1369.520 1083.960 1369.780 1084.220 ;
        RECT 1370.900 16.700 1371.160 16.960 ;
        RECT 1386.080 16.360 1386.340 16.620 ;
        RECT 1402.180 15.000 1402.440 15.260 ;
        RECT 1477.620 15.000 1477.880 15.260 ;
      LAYER met2 ;
        RECT 1357.010 1100.580 1357.290 1104.000 ;
        RECT 1357.010 1100.000 1357.300 1100.580 ;
        RECT 1357.160 1084.250 1357.300 1100.000 ;
        RECT 1357.100 1083.930 1357.360 1084.250 ;
        RECT 1369.520 1083.930 1369.780 1084.250 ;
        RECT 1369.580 38.490 1369.720 1083.930 ;
        RECT 1369.580 38.350 1371.100 38.490 ;
        RECT 1370.960 16.990 1371.100 38.350 ;
        RECT 1370.900 16.670 1371.160 16.990 ;
        RECT 1386.080 16.330 1386.340 16.650 ;
        RECT 1386.140 15.485 1386.280 16.330 ;
        RECT 1386.070 15.115 1386.350 15.485 ;
        RECT 1402.170 15.115 1402.450 15.485 ;
        RECT 1402.180 14.970 1402.440 15.115 ;
        RECT 1477.620 14.970 1477.880 15.290 ;
        RECT 1477.680 2.000 1477.820 14.970 ;
        RECT 1477.470 -4.000 1478.030 2.000 ;
      LAYER via2 ;
        RECT 1386.070 15.160 1386.350 15.440 ;
        RECT 1402.170 15.160 1402.450 15.440 ;
      LAYER met3 ;
        RECT 1386.045 15.450 1386.375 15.465 ;
        RECT 1402.145 15.450 1402.475 15.465 ;
        RECT 1386.045 15.150 1402.475 15.450 ;
        RECT 1386.045 15.135 1386.375 15.150 ;
        RECT 1402.145 15.135 1402.475 15.150 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1365.425 531.505 1365.595 579.615 ;
        RECT 1365.425 185.725 1365.595 227.715 ;
        RECT 1389.805 15.555 1389.975 19.975 ;
        RECT 1389.805 15.385 1391.815 15.555 ;
      LAYER mcon ;
        RECT 1365.425 579.445 1365.595 579.615 ;
        RECT 1365.425 227.545 1365.595 227.715 ;
        RECT 1389.805 19.805 1389.975 19.975 ;
        RECT 1391.645 15.385 1391.815 15.555 ;
      LAYER met1 ;
        RECT 1365.350 835.620 1365.670 835.680 ;
        RECT 1364.980 835.480 1365.670 835.620 ;
        RECT 1364.980 834.660 1365.120 835.480 ;
        RECT 1365.350 835.420 1365.670 835.480 ;
        RECT 1364.890 834.400 1365.210 834.660 ;
        RECT 1364.890 790.060 1365.210 790.120 ;
        RECT 1366.270 790.060 1366.590 790.120 ;
        RECT 1364.890 789.920 1366.590 790.060 ;
        RECT 1364.890 789.860 1365.210 789.920 ;
        RECT 1366.270 789.860 1366.590 789.920 ;
        RECT 1365.350 738.720 1365.670 738.780 ;
        RECT 1366.270 738.720 1366.590 738.780 ;
        RECT 1365.350 738.580 1366.590 738.720 ;
        RECT 1365.350 738.520 1365.670 738.580 ;
        RECT 1366.270 738.520 1366.590 738.580 ;
        RECT 1364.890 676.160 1365.210 676.220 ;
        RECT 1365.350 676.160 1365.670 676.220 ;
        RECT 1364.890 676.020 1365.670 676.160 ;
        RECT 1364.890 675.960 1365.210 676.020 ;
        RECT 1365.350 675.960 1365.670 676.020 ;
        RECT 1365.350 579.600 1365.670 579.660 ;
        RECT 1365.155 579.460 1365.670 579.600 ;
        RECT 1365.350 579.400 1365.670 579.460 ;
        RECT 1365.350 531.660 1365.670 531.720 ;
        RECT 1365.155 531.520 1365.670 531.660 ;
        RECT 1365.350 531.460 1365.670 531.520 ;
        RECT 1365.350 255.580 1365.670 255.640 ;
        RECT 1364.980 255.440 1365.670 255.580 ;
        RECT 1364.980 255.300 1365.120 255.440 ;
        RECT 1365.350 255.380 1365.670 255.440 ;
        RECT 1364.890 255.040 1365.210 255.300 ;
        RECT 1364.890 227.700 1365.210 227.760 ;
        RECT 1365.365 227.700 1365.655 227.745 ;
        RECT 1364.890 227.560 1365.655 227.700 ;
        RECT 1364.890 227.500 1365.210 227.560 ;
        RECT 1365.365 227.515 1365.655 227.560 ;
        RECT 1364.890 185.880 1365.210 185.940 ;
        RECT 1365.365 185.880 1365.655 185.925 ;
        RECT 1364.890 185.740 1365.655 185.880 ;
        RECT 1364.890 185.680 1365.210 185.740 ;
        RECT 1365.365 185.695 1365.655 185.740 ;
        RECT 1364.890 138.620 1365.210 138.680 ;
        RECT 1364.890 138.480 1365.580 138.620 ;
        RECT 1364.890 138.420 1365.210 138.480 ;
        RECT 1365.440 138.340 1365.580 138.480 ;
        RECT 1365.350 138.080 1365.670 138.340 ;
        RECT 1363.970 90.000 1364.290 90.060 ;
        RECT 1364.430 90.000 1364.750 90.060 ;
        RECT 1363.970 89.860 1364.750 90.000 ;
        RECT 1363.970 89.800 1364.290 89.860 ;
        RECT 1364.430 89.800 1364.750 89.860 ;
        RECT 1363.970 19.960 1364.290 20.020 ;
        RECT 1389.745 19.960 1390.035 20.005 ;
        RECT 1363.970 19.820 1390.035 19.960 ;
        RECT 1363.970 19.760 1364.290 19.820 ;
        RECT 1389.745 19.775 1390.035 19.820 ;
        RECT 1391.585 15.540 1391.875 15.585 ;
        RECT 1495.530 15.540 1495.850 15.600 ;
        RECT 1391.585 15.400 1495.850 15.540 ;
        RECT 1391.585 15.355 1391.875 15.400 ;
        RECT 1495.530 15.340 1495.850 15.400 ;
      LAYER via ;
        RECT 1365.380 835.420 1365.640 835.680 ;
        RECT 1364.920 834.400 1365.180 834.660 ;
        RECT 1364.920 789.860 1365.180 790.120 ;
        RECT 1366.300 789.860 1366.560 790.120 ;
        RECT 1365.380 738.520 1365.640 738.780 ;
        RECT 1366.300 738.520 1366.560 738.780 ;
        RECT 1364.920 675.960 1365.180 676.220 ;
        RECT 1365.380 675.960 1365.640 676.220 ;
        RECT 1365.380 579.400 1365.640 579.660 ;
        RECT 1365.380 531.460 1365.640 531.720 ;
        RECT 1365.380 255.380 1365.640 255.640 ;
        RECT 1364.920 255.040 1365.180 255.300 ;
        RECT 1364.920 227.500 1365.180 227.760 ;
        RECT 1364.920 185.680 1365.180 185.940 ;
        RECT 1364.920 138.420 1365.180 138.680 ;
        RECT 1365.380 138.080 1365.640 138.340 ;
        RECT 1364.000 89.800 1364.260 90.060 ;
        RECT 1364.460 89.800 1364.720 90.060 ;
        RECT 1364.000 19.760 1364.260 20.020 ;
        RECT 1495.560 15.340 1495.820 15.600 ;
      LAYER met2 ;
        RECT 1362.990 1100.650 1363.270 1104.000 ;
        RECT 1362.990 1100.510 1365.120 1100.650 ;
        RECT 1362.990 1100.000 1363.270 1100.510 ;
        RECT 1364.980 1028.570 1365.120 1100.510 ;
        RECT 1364.520 1028.430 1365.120 1028.570 ;
        RECT 1364.520 1027.890 1364.660 1028.430 ;
        RECT 1364.520 1027.750 1365.120 1027.890 ;
        RECT 1364.980 980.290 1365.120 1027.750 ;
        RECT 1364.980 980.150 1365.580 980.290 ;
        RECT 1365.440 966.010 1365.580 980.150 ;
        RECT 1364.980 965.870 1365.580 966.010 ;
        RECT 1364.980 863.445 1365.120 965.870 ;
        RECT 1364.910 863.075 1365.190 863.445 ;
        RECT 1365.370 862.395 1365.650 862.765 ;
        RECT 1365.440 835.710 1365.580 862.395 ;
        RECT 1365.380 835.390 1365.640 835.710 ;
        RECT 1364.920 834.370 1365.180 834.690 ;
        RECT 1364.980 790.150 1365.120 834.370 ;
        RECT 1364.920 789.830 1365.180 790.150 ;
        RECT 1366.300 789.830 1366.560 790.150 ;
        RECT 1366.360 738.810 1366.500 789.830 ;
        RECT 1365.380 738.490 1365.640 738.810 ;
        RECT 1366.300 738.490 1366.560 738.810 ;
        RECT 1365.440 676.250 1365.580 738.490 ;
        RECT 1364.920 675.930 1365.180 676.250 ;
        RECT 1365.380 675.930 1365.640 676.250 ;
        RECT 1364.980 641.820 1365.120 675.930 ;
        RECT 1364.980 641.680 1365.580 641.820 ;
        RECT 1365.440 579.690 1365.580 641.680 ;
        RECT 1365.380 579.370 1365.640 579.690 ;
        RECT 1365.380 531.430 1365.640 531.750 ;
        RECT 1365.440 255.670 1365.580 531.430 ;
        RECT 1365.380 255.350 1365.640 255.670 ;
        RECT 1364.920 255.010 1365.180 255.330 ;
        RECT 1364.980 227.790 1365.120 255.010 ;
        RECT 1364.920 227.470 1365.180 227.790 ;
        RECT 1364.920 185.650 1365.180 185.970 ;
        RECT 1364.980 138.710 1365.120 185.650 ;
        RECT 1364.920 138.390 1365.180 138.710 ;
        RECT 1365.380 138.050 1365.640 138.370 ;
        RECT 1365.440 111.250 1365.580 138.050 ;
        RECT 1364.520 111.110 1365.580 111.250 ;
        RECT 1364.520 90.090 1364.660 111.110 ;
        RECT 1364.000 89.770 1364.260 90.090 ;
        RECT 1364.460 89.770 1364.720 90.090 ;
        RECT 1364.060 20.050 1364.200 89.770 ;
        RECT 1364.000 19.730 1364.260 20.050 ;
        RECT 1495.560 15.310 1495.820 15.630 ;
        RECT 1495.620 2.000 1495.760 15.310 ;
        RECT 1495.410 -4.000 1495.970 2.000 ;
      LAYER via2 ;
        RECT 1364.910 863.120 1365.190 863.400 ;
        RECT 1365.370 862.440 1365.650 862.720 ;
      LAYER met3 ;
        RECT 1364.885 863.410 1365.215 863.425 ;
        RECT 1364.670 863.095 1365.215 863.410 ;
        RECT 1364.670 862.730 1364.970 863.095 ;
        RECT 1365.345 862.730 1365.675 862.745 ;
        RECT 1364.670 862.430 1365.675 862.730 ;
        RECT 1365.345 862.415 1365.675 862.430 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1408.665 1087.065 1408.835 1089.275 ;
      LAYER mcon ;
        RECT 1408.665 1089.105 1408.835 1089.275 ;
      LAYER met1 ;
        RECT 1408.605 1089.260 1408.895 1089.305 ;
        RECT 1493.690 1089.260 1494.010 1089.320 ;
        RECT 1408.605 1089.120 1494.010 1089.260 ;
        RECT 1408.605 1089.075 1408.895 1089.120 ;
        RECT 1493.690 1089.060 1494.010 1089.120 ;
        RECT 1369.030 1087.220 1369.350 1087.280 ;
        RECT 1408.605 1087.220 1408.895 1087.265 ;
        RECT 1369.030 1087.080 1408.895 1087.220 ;
        RECT 1369.030 1087.020 1369.350 1087.080 ;
        RECT 1408.605 1087.035 1408.895 1087.080 ;
        RECT 1493.690 15.200 1494.010 15.260 ;
        RECT 1513.010 15.200 1513.330 15.260 ;
        RECT 1493.690 15.060 1513.330 15.200 ;
        RECT 1493.690 15.000 1494.010 15.060 ;
        RECT 1513.010 15.000 1513.330 15.060 ;
      LAYER via ;
        RECT 1493.720 1089.060 1493.980 1089.320 ;
        RECT 1369.060 1087.020 1369.320 1087.280 ;
        RECT 1493.720 15.000 1493.980 15.260 ;
        RECT 1513.040 15.000 1513.300 15.260 ;
      LAYER met2 ;
        RECT 1368.970 1100.580 1369.250 1104.000 ;
        RECT 1368.970 1100.000 1369.260 1100.580 ;
        RECT 1369.120 1087.310 1369.260 1100.000 ;
        RECT 1493.720 1089.030 1493.980 1089.350 ;
        RECT 1369.060 1086.990 1369.320 1087.310 ;
        RECT 1493.780 15.290 1493.920 1089.030 ;
        RECT 1493.720 14.970 1493.980 15.290 ;
        RECT 1513.040 14.970 1513.300 15.290 ;
        RECT 1513.100 2.000 1513.240 14.970 ;
        RECT 1512.890 -4.000 1513.450 2.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 710.310 44.100 710.630 44.160 ;
        RECT 1091.190 44.100 1091.510 44.160 ;
        RECT 710.310 43.960 1091.510 44.100 ;
        RECT 710.310 43.900 710.630 43.960 ;
        RECT 1091.190 43.900 1091.510 43.960 ;
      LAYER via ;
        RECT 710.340 43.900 710.600 44.160 ;
        RECT 1091.220 43.900 1091.480 44.160 ;
      LAYER met2 ;
        RECT 1093.430 1100.650 1093.710 1104.000 ;
        RECT 1092.200 1100.510 1093.710 1100.650 ;
        RECT 1092.200 1088.410 1092.340 1100.510 ;
        RECT 1093.430 1100.000 1093.710 1100.510 ;
        RECT 1091.280 1088.270 1092.340 1088.410 ;
        RECT 1091.280 44.190 1091.420 1088.270 ;
        RECT 710.340 43.870 710.600 44.190 ;
        RECT 1091.220 43.870 1091.480 44.190 ;
        RECT 710.400 2.000 710.540 43.870 ;
        RECT 710.190 -4.000 710.750 2.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1409.125 1085.705 1409.295 1087.235 ;
      LAYER mcon ;
        RECT 1409.125 1087.065 1409.295 1087.235 ;
      LAYER met1 ;
        RECT 1409.065 1087.220 1409.355 1087.265 ;
        RECT 1409.065 1087.080 1463.100 1087.220 ;
        RECT 1409.065 1087.035 1409.355 1087.080 ;
        RECT 1462.960 1086.880 1463.100 1087.080 ;
        RECT 1514.850 1086.880 1515.170 1086.940 ;
        RECT 1462.960 1086.740 1515.170 1086.880 ;
        RECT 1514.850 1086.680 1515.170 1086.740 ;
        RECT 1375.470 1085.860 1375.790 1085.920 ;
        RECT 1409.065 1085.860 1409.355 1085.905 ;
        RECT 1375.470 1085.720 1409.355 1085.860 ;
        RECT 1375.470 1085.660 1375.790 1085.720 ;
        RECT 1409.065 1085.675 1409.355 1085.720 ;
        RECT 1514.850 16.220 1515.170 16.280 ;
        RECT 1530.950 16.220 1531.270 16.280 ;
        RECT 1514.850 16.080 1531.270 16.220 ;
        RECT 1514.850 16.020 1515.170 16.080 ;
        RECT 1530.950 16.020 1531.270 16.080 ;
      LAYER via ;
        RECT 1514.880 1086.680 1515.140 1086.940 ;
        RECT 1375.500 1085.660 1375.760 1085.920 ;
        RECT 1514.880 16.020 1515.140 16.280 ;
        RECT 1530.980 16.020 1531.240 16.280 ;
      LAYER met2 ;
        RECT 1375.410 1100.580 1375.690 1104.000 ;
        RECT 1375.410 1100.000 1375.700 1100.580 ;
        RECT 1375.560 1085.950 1375.700 1100.000 ;
        RECT 1514.880 1086.650 1515.140 1086.970 ;
        RECT 1375.500 1085.630 1375.760 1085.950 ;
        RECT 1514.940 16.310 1515.080 1086.650 ;
        RECT 1514.880 15.990 1515.140 16.310 ;
        RECT 1530.980 15.990 1531.240 16.310 ;
        RECT 1531.040 2.000 1531.180 15.990 ;
        RECT 1530.830 -4.000 1531.390 2.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1381.450 1086.880 1381.770 1086.940 ;
        RECT 1386.510 1086.880 1386.830 1086.940 ;
        RECT 1381.450 1086.740 1386.830 1086.880 ;
        RECT 1381.450 1086.680 1381.770 1086.740 ;
        RECT 1386.510 1086.680 1386.830 1086.740 ;
        RECT 1548.890 16.900 1549.210 16.960 ;
        RECT 1400.860 16.760 1549.210 16.900 ;
        RECT 1386.510 16.560 1386.830 16.620 ;
        RECT 1400.860 16.560 1401.000 16.760 ;
        RECT 1548.890 16.700 1549.210 16.760 ;
        RECT 1386.510 16.420 1401.000 16.560 ;
        RECT 1386.510 16.360 1386.830 16.420 ;
      LAYER via ;
        RECT 1381.480 1086.680 1381.740 1086.940 ;
        RECT 1386.540 1086.680 1386.800 1086.940 ;
        RECT 1386.540 16.360 1386.800 16.620 ;
        RECT 1548.920 16.700 1549.180 16.960 ;
      LAYER met2 ;
        RECT 1381.390 1100.580 1381.670 1104.000 ;
        RECT 1381.390 1100.000 1381.680 1100.580 ;
        RECT 1381.540 1086.970 1381.680 1100.000 ;
        RECT 1381.480 1086.650 1381.740 1086.970 ;
        RECT 1386.540 1086.650 1386.800 1086.970 ;
        RECT 1386.600 16.650 1386.740 1086.650 ;
        RECT 1548.920 16.670 1549.180 16.990 ;
        RECT 1386.540 16.330 1386.800 16.650 ;
        RECT 1548.980 2.000 1549.120 16.670 ;
        RECT 1548.770 -4.000 1549.330 2.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1414.645 1083.665 1414.815 1086.895 ;
        RECT 1456.045 1083.665 1456.215 1086.555 ;
      LAYER mcon ;
        RECT 1414.645 1086.725 1414.815 1086.895 ;
        RECT 1456.045 1086.385 1456.215 1086.555 ;
      LAYER met1 ;
        RECT 1387.430 1086.880 1387.750 1086.940 ;
        RECT 1414.585 1086.880 1414.875 1086.925 ;
        RECT 1387.430 1086.740 1414.875 1086.880 ;
        RECT 1387.430 1086.680 1387.750 1086.740 ;
        RECT 1414.585 1086.695 1414.875 1086.740 ;
        RECT 1455.985 1086.540 1456.275 1086.585 ;
        RECT 1562.690 1086.540 1563.010 1086.600 ;
        RECT 1455.985 1086.400 1563.010 1086.540 ;
        RECT 1455.985 1086.355 1456.275 1086.400 ;
        RECT 1562.690 1086.340 1563.010 1086.400 ;
        RECT 1414.585 1083.820 1414.875 1083.865 ;
        RECT 1455.985 1083.820 1456.275 1083.865 ;
        RECT 1414.585 1083.680 1456.275 1083.820 ;
        RECT 1414.585 1083.635 1414.875 1083.680 ;
        RECT 1455.985 1083.635 1456.275 1083.680 ;
        RECT 1562.690 16.900 1563.010 16.960 ;
        RECT 1566.830 16.900 1567.150 16.960 ;
        RECT 1562.690 16.760 1567.150 16.900 ;
        RECT 1562.690 16.700 1563.010 16.760 ;
        RECT 1566.830 16.700 1567.150 16.760 ;
      LAYER via ;
        RECT 1387.460 1086.680 1387.720 1086.940 ;
        RECT 1562.720 1086.340 1562.980 1086.600 ;
        RECT 1562.720 16.700 1562.980 16.960 ;
        RECT 1566.860 16.700 1567.120 16.960 ;
      LAYER met2 ;
        RECT 1387.370 1100.580 1387.650 1104.000 ;
        RECT 1387.370 1100.000 1387.660 1100.580 ;
        RECT 1387.520 1086.970 1387.660 1100.000 ;
        RECT 1387.460 1086.650 1387.720 1086.970 ;
        RECT 1562.720 1086.310 1562.980 1086.630 ;
        RECT 1562.780 16.990 1562.920 1086.310 ;
        RECT 1562.720 16.670 1562.980 16.990 ;
        RECT 1566.860 16.670 1567.120 16.990 ;
        RECT 1566.920 2.000 1567.060 16.670 ;
        RECT 1566.710 -4.000 1567.270 2.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1438.105 20.825 1440.115 20.995 ;
        RECT 1438.105 19.975 1438.275 20.825 ;
        RECT 1439.945 20.485 1440.115 20.825 ;
        RECT 1437.645 19.805 1438.275 19.975 ;
      LAYER met1 ;
        RECT 1393.870 1086.200 1394.190 1086.260 ;
        RECT 1418.250 1086.200 1418.570 1086.260 ;
        RECT 1393.870 1086.060 1418.570 1086.200 ;
        RECT 1393.870 1086.000 1394.190 1086.060 ;
        RECT 1418.250 1086.000 1418.570 1086.060 ;
        RECT 1418.250 20.640 1418.570 20.700 ;
        RECT 1439.885 20.640 1440.175 20.685 ;
        RECT 1531.870 20.640 1532.190 20.700 ;
        RECT 1418.250 20.500 1430.900 20.640 ;
        RECT 1418.250 20.440 1418.570 20.500 ;
        RECT 1430.760 19.960 1430.900 20.500 ;
        RECT 1439.885 20.500 1532.190 20.640 ;
        RECT 1439.885 20.455 1440.175 20.500 ;
        RECT 1531.870 20.440 1532.190 20.500 ;
        RECT 1555.330 20.300 1555.650 20.360 ;
        RECT 1584.770 20.300 1585.090 20.360 ;
        RECT 1555.330 20.160 1585.090 20.300 ;
        RECT 1555.330 20.100 1555.650 20.160 ;
        RECT 1584.770 20.100 1585.090 20.160 ;
        RECT 1437.585 19.960 1437.875 20.005 ;
        RECT 1430.760 19.820 1437.875 19.960 ;
        RECT 1437.585 19.775 1437.875 19.820 ;
      LAYER via ;
        RECT 1393.900 1086.000 1394.160 1086.260 ;
        RECT 1418.280 1086.000 1418.540 1086.260 ;
        RECT 1418.280 20.440 1418.540 20.700 ;
        RECT 1531.900 20.440 1532.160 20.700 ;
        RECT 1555.360 20.100 1555.620 20.360 ;
        RECT 1584.800 20.100 1585.060 20.360 ;
      LAYER met2 ;
        RECT 1393.810 1100.580 1394.090 1104.000 ;
        RECT 1393.810 1100.000 1394.100 1100.580 ;
        RECT 1393.960 1086.290 1394.100 1100.000 ;
        RECT 1393.900 1085.970 1394.160 1086.290 ;
        RECT 1418.280 1085.970 1418.540 1086.290 ;
        RECT 1418.340 20.730 1418.480 1085.970 ;
        RECT 1418.280 20.410 1418.540 20.730 ;
        RECT 1531.890 20.555 1532.170 20.925 ;
        RECT 1555.350 20.555 1555.630 20.925 ;
        RECT 1531.900 20.410 1532.160 20.555 ;
        RECT 1555.420 20.390 1555.560 20.555 ;
        RECT 1555.360 20.070 1555.620 20.390 ;
        RECT 1584.800 20.070 1585.060 20.390 ;
        RECT 1584.860 2.000 1585.000 20.070 ;
        RECT 1584.650 -4.000 1585.210 2.000 ;
      LAYER via2 ;
        RECT 1531.890 20.600 1532.170 20.880 ;
        RECT 1555.350 20.600 1555.630 20.880 ;
      LAYER met3 ;
        RECT 1531.865 20.890 1532.195 20.905 ;
        RECT 1555.325 20.890 1555.655 20.905 ;
        RECT 1531.865 20.590 1555.655 20.890 ;
        RECT 1531.865 20.575 1532.195 20.590 ;
        RECT 1555.325 20.575 1555.655 20.590 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1399.850 20.980 1400.170 21.040 ;
        RECT 1602.250 20.980 1602.570 21.040 ;
        RECT 1399.850 20.840 1602.570 20.980 ;
        RECT 1399.850 20.780 1400.170 20.840 ;
        RECT 1602.250 20.780 1602.570 20.840 ;
      LAYER via ;
        RECT 1399.880 20.780 1400.140 21.040 ;
        RECT 1602.280 20.780 1602.540 21.040 ;
      LAYER met2 ;
        RECT 1399.790 1100.580 1400.070 1104.000 ;
        RECT 1399.790 1100.000 1400.080 1100.580 ;
        RECT 1399.940 21.070 1400.080 1100.000 ;
        RECT 1399.880 20.750 1400.140 21.070 ;
        RECT 1602.280 20.750 1602.540 21.070 ;
        RECT 1602.340 2.000 1602.480 20.750 ;
        RECT 1602.130 -4.000 1602.690 2.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1406.750 21.320 1407.070 21.380 ;
        RECT 1620.190 21.320 1620.510 21.380 ;
        RECT 1406.750 21.180 1620.510 21.320 ;
        RECT 1406.750 21.120 1407.070 21.180 ;
        RECT 1620.190 21.120 1620.510 21.180 ;
      LAYER via ;
        RECT 1406.780 21.120 1407.040 21.380 ;
        RECT 1620.220 21.120 1620.480 21.380 ;
      LAYER met2 ;
        RECT 1405.770 1100.650 1406.050 1104.000 ;
        RECT 1405.770 1100.510 1406.980 1100.650 ;
        RECT 1405.770 1100.000 1406.050 1100.510 ;
        RECT 1406.840 21.410 1406.980 1100.510 ;
        RECT 1406.780 21.090 1407.040 21.410 ;
        RECT 1620.220 21.090 1620.480 21.410 ;
        RECT 1620.280 2.000 1620.420 21.090 ;
        RECT 1620.070 -4.000 1620.630 2.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1414.185 965.685 1414.355 1007.335 ;
        RECT 1413.725 572.645 1413.895 579.955 ;
        RECT 1413.725 476.085 1413.895 524.195 ;
        RECT 1413.725 379.525 1413.895 386.835 ;
      LAYER mcon ;
        RECT 1414.185 1007.165 1414.355 1007.335 ;
        RECT 1413.725 579.785 1413.895 579.955 ;
        RECT 1413.725 524.025 1413.895 524.195 ;
        RECT 1413.725 386.665 1413.895 386.835 ;
      LAYER met1 ;
        RECT 1413.190 1027.720 1413.510 1027.780 ;
        RECT 1414.110 1027.720 1414.430 1027.780 ;
        RECT 1413.190 1027.580 1414.430 1027.720 ;
        RECT 1413.190 1027.520 1413.510 1027.580 ;
        RECT 1414.110 1027.520 1414.430 1027.580 ;
        RECT 1414.110 1007.320 1414.430 1007.380 ;
        RECT 1413.915 1007.180 1414.430 1007.320 ;
        RECT 1414.110 1007.120 1414.430 1007.180 ;
        RECT 1414.110 965.840 1414.430 965.900 ;
        RECT 1413.915 965.700 1414.430 965.840 ;
        RECT 1414.110 965.640 1414.430 965.700 ;
        RECT 1413.650 917.900 1413.970 917.960 ;
        RECT 1414.570 917.900 1414.890 917.960 ;
        RECT 1413.650 917.760 1414.890 917.900 ;
        RECT 1413.650 917.700 1413.970 917.760 ;
        RECT 1414.570 917.700 1414.890 917.760 ;
        RECT 1414.110 910.760 1414.430 910.820 ;
        RECT 1414.570 910.760 1414.890 910.820 ;
        RECT 1414.110 910.620 1414.890 910.760 ;
        RECT 1414.110 910.560 1414.430 910.620 ;
        RECT 1414.570 910.560 1414.890 910.620 ;
        RECT 1413.190 814.200 1413.510 814.260 ;
        RECT 1414.110 814.200 1414.430 814.260 ;
        RECT 1413.190 814.060 1414.430 814.200 ;
        RECT 1413.190 814.000 1413.510 814.060 ;
        RECT 1414.110 814.000 1414.430 814.060 ;
        RECT 1413.665 579.940 1413.955 579.985 ;
        RECT 1414.110 579.940 1414.430 580.000 ;
        RECT 1413.665 579.800 1414.430 579.940 ;
        RECT 1413.665 579.755 1413.955 579.800 ;
        RECT 1414.110 579.740 1414.430 579.800 ;
        RECT 1413.650 572.800 1413.970 572.860 ;
        RECT 1413.455 572.660 1413.970 572.800 ;
        RECT 1413.650 572.600 1413.970 572.660 ;
        RECT 1413.650 524.180 1413.970 524.240 ;
        RECT 1413.455 524.040 1413.970 524.180 ;
        RECT 1413.650 523.980 1413.970 524.040 ;
        RECT 1413.650 476.240 1413.970 476.300 ;
        RECT 1413.455 476.100 1413.970 476.240 ;
        RECT 1413.650 476.040 1413.970 476.100 ;
        RECT 1413.665 386.820 1413.955 386.865 ;
        RECT 1414.110 386.820 1414.430 386.880 ;
        RECT 1413.665 386.680 1414.430 386.820 ;
        RECT 1413.665 386.635 1413.955 386.680 ;
        RECT 1414.110 386.620 1414.430 386.680 ;
        RECT 1413.650 379.680 1413.970 379.740 ;
        RECT 1413.455 379.540 1413.970 379.680 ;
        RECT 1413.650 379.480 1413.970 379.540 ;
        RECT 1413.650 338.200 1413.970 338.260 ;
        RECT 1414.110 338.200 1414.430 338.260 ;
        RECT 1413.650 338.060 1414.430 338.200 ;
        RECT 1413.650 338.000 1413.970 338.060 ;
        RECT 1414.110 338.000 1414.430 338.060 ;
        RECT 1413.650 241.300 1413.970 241.360 ;
        RECT 1414.110 241.300 1414.430 241.360 ;
        RECT 1413.650 241.160 1414.430 241.300 ;
        RECT 1413.650 241.100 1413.970 241.160 ;
        RECT 1414.110 241.100 1414.430 241.160 ;
        RECT 1413.650 186.560 1413.970 186.620 ;
        RECT 1414.110 186.560 1414.430 186.620 ;
        RECT 1413.650 186.420 1414.430 186.560 ;
        RECT 1413.650 186.360 1413.970 186.420 ;
        RECT 1414.110 186.360 1414.430 186.420 ;
        RECT 1413.650 21.660 1413.970 21.720 ;
        RECT 1638.130 21.660 1638.450 21.720 ;
        RECT 1413.650 21.520 1638.450 21.660 ;
        RECT 1413.650 21.460 1413.970 21.520 ;
        RECT 1638.130 21.460 1638.450 21.520 ;
      LAYER via ;
        RECT 1413.220 1027.520 1413.480 1027.780 ;
        RECT 1414.140 1027.520 1414.400 1027.780 ;
        RECT 1414.140 1007.120 1414.400 1007.380 ;
        RECT 1414.140 965.640 1414.400 965.900 ;
        RECT 1413.680 917.700 1413.940 917.960 ;
        RECT 1414.600 917.700 1414.860 917.960 ;
        RECT 1414.140 910.560 1414.400 910.820 ;
        RECT 1414.600 910.560 1414.860 910.820 ;
        RECT 1413.220 814.000 1413.480 814.260 ;
        RECT 1414.140 814.000 1414.400 814.260 ;
        RECT 1414.140 579.740 1414.400 580.000 ;
        RECT 1413.680 572.600 1413.940 572.860 ;
        RECT 1413.680 523.980 1413.940 524.240 ;
        RECT 1413.680 476.040 1413.940 476.300 ;
        RECT 1414.140 386.620 1414.400 386.880 ;
        RECT 1413.680 379.480 1413.940 379.740 ;
        RECT 1413.680 338.000 1413.940 338.260 ;
        RECT 1414.140 338.000 1414.400 338.260 ;
        RECT 1413.680 241.100 1413.940 241.360 ;
        RECT 1414.140 241.100 1414.400 241.360 ;
        RECT 1413.680 186.360 1413.940 186.620 ;
        RECT 1414.140 186.360 1414.400 186.620 ;
        RECT 1413.680 21.460 1413.940 21.720 ;
        RECT 1638.160 21.460 1638.420 21.720 ;
      LAYER met2 ;
        RECT 1412.210 1100.580 1412.490 1104.000 ;
        RECT 1412.210 1100.000 1412.500 1100.580 ;
        RECT 1412.360 1055.885 1412.500 1100.000 ;
        RECT 1412.290 1055.515 1412.570 1055.885 ;
        RECT 1413.210 1055.515 1413.490 1055.885 ;
        RECT 1413.280 1027.810 1413.420 1055.515 ;
        RECT 1413.220 1027.490 1413.480 1027.810 ;
        RECT 1414.140 1027.490 1414.400 1027.810 ;
        RECT 1414.200 1007.410 1414.340 1027.490 ;
        RECT 1414.140 1007.090 1414.400 1007.410 ;
        RECT 1414.140 965.610 1414.400 965.930 ;
        RECT 1414.200 959.210 1414.340 965.610 ;
        RECT 1414.200 959.070 1414.800 959.210 ;
        RECT 1414.660 917.990 1414.800 959.070 ;
        RECT 1413.680 917.845 1413.940 917.990 ;
        RECT 1414.600 917.845 1414.860 917.990 ;
        RECT 1413.670 917.475 1413.950 917.845 ;
        RECT 1414.590 917.475 1414.870 917.845 ;
        RECT 1414.660 910.850 1414.800 917.475 ;
        RECT 1414.140 910.530 1414.400 910.850 ;
        RECT 1414.600 910.530 1414.860 910.850 ;
        RECT 1414.200 821.285 1414.340 910.530 ;
        RECT 1413.210 820.915 1413.490 821.285 ;
        RECT 1414.130 820.915 1414.410 821.285 ;
        RECT 1413.280 814.290 1413.420 820.915 ;
        RECT 1413.220 813.970 1413.480 814.290 ;
        RECT 1414.140 813.970 1414.400 814.290 ;
        RECT 1414.200 641.820 1414.340 813.970 ;
        RECT 1413.740 641.680 1414.340 641.820 ;
        RECT 1413.740 628.050 1413.880 641.680 ;
        RECT 1413.740 627.910 1414.340 628.050 ;
        RECT 1414.200 580.030 1414.340 627.910 ;
        RECT 1414.140 579.710 1414.400 580.030 ;
        RECT 1413.680 572.570 1413.940 572.890 ;
        RECT 1413.740 524.270 1413.880 572.570 ;
        RECT 1413.680 523.950 1413.940 524.270 ;
        RECT 1413.680 476.010 1413.940 476.330 ;
        RECT 1413.740 445.130 1413.880 476.010 ;
        RECT 1413.740 444.990 1414.340 445.130 ;
        RECT 1414.200 386.910 1414.340 444.990 ;
        RECT 1414.140 386.590 1414.400 386.910 ;
        RECT 1413.680 379.450 1413.940 379.770 ;
        RECT 1413.740 338.290 1413.880 379.450 ;
        RECT 1413.680 337.970 1413.940 338.290 ;
        RECT 1414.140 337.970 1414.400 338.290 ;
        RECT 1414.200 265.610 1414.340 337.970 ;
        RECT 1413.740 265.470 1414.340 265.610 ;
        RECT 1413.740 241.390 1413.880 265.470 ;
        RECT 1413.680 241.070 1413.940 241.390 ;
        RECT 1414.140 241.070 1414.400 241.390 ;
        RECT 1414.200 186.650 1414.340 241.070 ;
        RECT 1413.680 186.330 1413.940 186.650 ;
        RECT 1414.140 186.330 1414.400 186.650 ;
        RECT 1413.740 131.650 1413.880 186.330 ;
        RECT 1413.740 131.510 1414.340 131.650 ;
        RECT 1414.200 62.290 1414.340 131.510 ;
        RECT 1414.200 62.150 1414.800 62.290 ;
        RECT 1414.660 61.610 1414.800 62.150 ;
        RECT 1413.740 61.470 1414.800 61.610 ;
        RECT 1413.740 21.750 1413.880 61.470 ;
        RECT 1413.680 21.430 1413.940 21.750 ;
        RECT 1638.160 21.430 1638.420 21.750 ;
        RECT 1638.220 2.000 1638.360 21.430 ;
        RECT 1638.010 -4.000 1638.570 2.000 ;
      LAYER via2 ;
        RECT 1412.290 1055.560 1412.570 1055.840 ;
        RECT 1413.210 1055.560 1413.490 1055.840 ;
        RECT 1413.670 917.520 1413.950 917.800 ;
        RECT 1414.590 917.520 1414.870 917.800 ;
        RECT 1413.210 820.960 1413.490 821.240 ;
        RECT 1414.130 820.960 1414.410 821.240 ;
      LAYER met3 ;
        RECT 1412.265 1055.850 1412.595 1055.865 ;
        RECT 1413.185 1055.850 1413.515 1055.865 ;
        RECT 1412.265 1055.550 1413.515 1055.850 ;
        RECT 1412.265 1055.535 1412.595 1055.550 ;
        RECT 1413.185 1055.535 1413.515 1055.550 ;
        RECT 1413.645 917.810 1413.975 917.825 ;
        RECT 1414.565 917.810 1414.895 917.825 ;
        RECT 1413.645 917.510 1414.895 917.810 ;
        RECT 1413.645 917.495 1413.975 917.510 ;
        RECT 1414.565 917.495 1414.895 917.510 ;
        RECT 1413.185 821.250 1413.515 821.265 ;
        RECT 1414.105 821.250 1414.435 821.265 ;
        RECT 1413.185 820.950 1414.435 821.250 ;
        RECT 1413.185 820.935 1413.515 820.950 ;
        RECT 1414.105 820.935 1414.435 820.950 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1419.705 476.085 1419.875 524.195 ;
        RECT 1419.705 379.525 1419.875 427.635 ;
        RECT 1419.705 283.305 1419.875 331.075 ;
        RECT 1419.705 234.685 1419.875 282.795 ;
        RECT 1419.705 41.565 1419.875 48.875 ;
      LAYER mcon ;
        RECT 1419.705 524.025 1419.875 524.195 ;
        RECT 1419.705 427.465 1419.875 427.635 ;
        RECT 1419.705 330.905 1419.875 331.075 ;
        RECT 1419.705 282.625 1419.875 282.795 ;
        RECT 1419.705 48.705 1419.875 48.875 ;
      LAYER met1 ;
        RECT 1418.710 1062.740 1419.030 1062.800 ;
        RECT 1420.090 1062.740 1420.410 1062.800 ;
        RECT 1418.710 1062.600 1420.410 1062.740 ;
        RECT 1418.710 1062.540 1419.030 1062.600 ;
        RECT 1420.090 1062.540 1420.410 1062.600 ;
        RECT 1419.170 1055.600 1419.490 1055.660 ;
        RECT 1420.090 1055.600 1420.410 1055.660 ;
        RECT 1419.170 1055.460 1420.410 1055.600 ;
        RECT 1419.170 1055.400 1419.490 1055.460 ;
        RECT 1420.090 1055.400 1420.410 1055.460 ;
        RECT 1419.170 959.040 1419.490 959.100 ;
        RECT 1420.090 959.040 1420.410 959.100 ;
        RECT 1419.170 958.900 1420.410 959.040 ;
        RECT 1419.170 958.840 1419.490 958.900 ;
        RECT 1420.090 958.840 1420.410 958.900 ;
        RECT 1419.170 862.480 1419.490 862.540 ;
        RECT 1420.090 862.480 1420.410 862.540 ;
        RECT 1419.170 862.340 1420.410 862.480 ;
        RECT 1419.170 862.280 1419.490 862.340 ;
        RECT 1420.090 862.280 1420.410 862.340 ;
        RECT 1419.170 766.260 1419.490 766.320 ;
        RECT 1419.630 766.260 1419.950 766.320 ;
        RECT 1419.170 766.120 1419.950 766.260 ;
        RECT 1419.170 766.060 1419.490 766.120 ;
        RECT 1419.630 766.060 1419.950 766.120 ;
        RECT 1420.090 669.360 1420.410 669.420 ;
        RECT 1421.470 669.360 1421.790 669.420 ;
        RECT 1420.090 669.220 1421.790 669.360 ;
        RECT 1420.090 669.160 1420.410 669.220 ;
        RECT 1421.470 669.160 1421.790 669.220 ;
        RECT 1419.645 524.180 1419.935 524.225 ;
        RECT 1420.090 524.180 1420.410 524.240 ;
        RECT 1419.645 524.040 1420.410 524.180 ;
        RECT 1419.645 523.995 1419.935 524.040 ;
        RECT 1420.090 523.980 1420.410 524.040 ;
        RECT 1419.630 476.240 1419.950 476.300 ;
        RECT 1419.435 476.100 1419.950 476.240 ;
        RECT 1419.630 476.040 1419.950 476.100 ;
        RECT 1419.630 427.620 1419.950 427.680 ;
        RECT 1419.435 427.480 1419.950 427.620 ;
        RECT 1419.630 427.420 1419.950 427.480 ;
        RECT 1419.645 379.680 1419.935 379.725 ;
        RECT 1420.090 379.680 1420.410 379.740 ;
        RECT 1419.645 379.540 1420.410 379.680 ;
        RECT 1419.645 379.495 1419.935 379.540 ;
        RECT 1420.090 379.480 1420.410 379.540 ;
        RECT 1419.645 331.060 1419.935 331.105 ;
        RECT 1420.090 331.060 1420.410 331.120 ;
        RECT 1419.645 330.920 1420.410 331.060 ;
        RECT 1419.645 330.875 1419.935 330.920 ;
        RECT 1420.090 330.860 1420.410 330.920 ;
        RECT 1419.630 283.460 1419.950 283.520 ;
        RECT 1419.435 283.320 1419.950 283.460 ;
        RECT 1419.630 283.260 1419.950 283.320 ;
        RECT 1419.630 282.780 1419.950 282.840 ;
        RECT 1419.435 282.640 1419.950 282.780 ;
        RECT 1419.630 282.580 1419.950 282.640 ;
        RECT 1419.645 234.840 1419.935 234.885 ;
        RECT 1420.090 234.840 1420.410 234.900 ;
        RECT 1419.645 234.700 1420.410 234.840 ;
        RECT 1419.645 234.655 1419.935 234.700 ;
        RECT 1420.090 234.640 1420.410 234.700 ;
        RECT 1419.630 192.680 1419.950 192.740 ;
        RECT 1421.470 192.680 1421.790 192.740 ;
        RECT 1419.630 192.540 1421.790 192.680 ;
        RECT 1419.630 192.480 1419.950 192.540 ;
        RECT 1421.470 192.480 1421.790 192.540 ;
        RECT 1420.090 145.080 1420.410 145.140 ;
        RECT 1421.470 145.080 1421.790 145.140 ;
        RECT 1420.090 144.940 1421.790 145.080 ;
        RECT 1420.090 144.880 1420.410 144.940 ;
        RECT 1421.470 144.880 1421.790 144.940 ;
        RECT 1419.645 48.860 1419.935 48.905 ;
        RECT 1420.090 48.860 1420.410 48.920 ;
        RECT 1419.645 48.720 1420.410 48.860 ;
        RECT 1419.645 48.675 1419.935 48.720 ;
        RECT 1420.090 48.660 1420.410 48.720 ;
        RECT 1419.630 41.720 1419.950 41.780 ;
        RECT 1419.435 41.580 1419.950 41.720 ;
        RECT 1419.630 41.520 1419.950 41.580 ;
        RECT 1419.630 22.680 1419.950 22.740 ;
        RECT 1656.070 22.680 1656.390 22.740 ;
        RECT 1419.630 22.540 1656.390 22.680 ;
        RECT 1419.630 22.480 1419.950 22.540 ;
        RECT 1656.070 22.480 1656.390 22.540 ;
      LAYER via ;
        RECT 1418.740 1062.540 1419.000 1062.800 ;
        RECT 1420.120 1062.540 1420.380 1062.800 ;
        RECT 1419.200 1055.400 1419.460 1055.660 ;
        RECT 1420.120 1055.400 1420.380 1055.660 ;
        RECT 1419.200 958.840 1419.460 959.100 ;
        RECT 1420.120 958.840 1420.380 959.100 ;
        RECT 1419.200 862.280 1419.460 862.540 ;
        RECT 1420.120 862.280 1420.380 862.540 ;
        RECT 1419.200 766.060 1419.460 766.320 ;
        RECT 1419.660 766.060 1419.920 766.320 ;
        RECT 1420.120 669.160 1420.380 669.420 ;
        RECT 1421.500 669.160 1421.760 669.420 ;
        RECT 1420.120 523.980 1420.380 524.240 ;
        RECT 1419.660 476.040 1419.920 476.300 ;
        RECT 1419.660 427.420 1419.920 427.680 ;
        RECT 1420.120 379.480 1420.380 379.740 ;
        RECT 1420.120 330.860 1420.380 331.120 ;
        RECT 1419.660 283.260 1419.920 283.520 ;
        RECT 1419.660 282.580 1419.920 282.840 ;
        RECT 1420.120 234.640 1420.380 234.900 ;
        RECT 1419.660 192.480 1419.920 192.740 ;
        RECT 1421.500 192.480 1421.760 192.740 ;
        RECT 1420.120 144.880 1420.380 145.140 ;
        RECT 1421.500 144.880 1421.760 145.140 ;
        RECT 1420.120 48.660 1420.380 48.920 ;
        RECT 1419.660 41.520 1419.920 41.780 ;
        RECT 1419.660 22.480 1419.920 22.740 ;
        RECT 1656.100 22.480 1656.360 22.740 ;
      LAYER met2 ;
        RECT 1418.190 1100.650 1418.470 1104.000 ;
        RECT 1418.190 1100.510 1418.940 1100.650 ;
        RECT 1418.190 1100.000 1418.470 1100.510 ;
        RECT 1418.800 1062.830 1418.940 1100.510 ;
        RECT 1418.740 1062.510 1419.000 1062.830 ;
        RECT 1420.120 1062.510 1420.380 1062.830 ;
        RECT 1420.180 1055.690 1420.320 1062.510 ;
        RECT 1419.200 1055.370 1419.460 1055.690 ;
        RECT 1420.120 1055.370 1420.380 1055.690 ;
        RECT 1419.260 1007.605 1419.400 1055.370 ;
        RECT 1419.190 1007.235 1419.470 1007.605 ;
        RECT 1420.110 1007.235 1420.390 1007.605 ;
        RECT 1420.180 959.130 1420.320 1007.235 ;
        RECT 1419.200 958.810 1419.460 959.130 ;
        RECT 1420.120 958.810 1420.380 959.130 ;
        RECT 1419.260 911.045 1419.400 958.810 ;
        RECT 1419.190 910.675 1419.470 911.045 ;
        RECT 1420.110 910.675 1420.390 911.045 ;
        RECT 1420.180 862.570 1420.320 910.675 ;
        RECT 1419.200 862.250 1419.460 862.570 ;
        RECT 1420.120 862.250 1420.380 862.570 ;
        RECT 1419.260 814.485 1419.400 862.250 ;
        RECT 1419.190 814.115 1419.470 814.485 ;
        RECT 1420.110 814.115 1420.390 814.485 ;
        RECT 1420.180 773.570 1420.320 814.115 ;
        RECT 1419.720 773.430 1420.320 773.570 ;
        RECT 1419.720 766.350 1419.860 773.430 ;
        RECT 1419.200 766.030 1419.460 766.350 ;
        RECT 1419.660 766.030 1419.920 766.350 ;
        RECT 1419.260 738.720 1419.400 766.030 ;
        RECT 1419.260 738.580 1419.860 738.720 ;
        RECT 1419.720 693.330 1419.860 738.580 ;
        RECT 1419.260 693.190 1419.860 693.330 ;
        RECT 1419.260 689.930 1419.400 693.190 ;
        RECT 1419.260 689.790 1419.860 689.930 ;
        RECT 1419.720 669.530 1419.860 689.790 ;
        RECT 1419.720 669.450 1420.320 669.530 ;
        RECT 1419.720 669.390 1420.380 669.450 ;
        RECT 1420.120 669.130 1420.380 669.390 ;
        RECT 1421.500 669.130 1421.760 669.450 ;
        RECT 1420.180 668.975 1420.320 669.130 ;
        RECT 1421.560 621.365 1421.700 669.130 ;
        RECT 1421.490 620.995 1421.770 621.365 ;
        RECT 1420.110 531.235 1420.390 531.605 ;
        RECT 1420.180 524.270 1420.320 531.235 ;
        RECT 1420.120 523.950 1420.380 524.270 ;
        RECT 1419.660 476.010 1419.920 476.330 ;
        RECT 1419.720 427.710 1419.860 476.010 ;
        RECT 1419.660 427.390 1419.920 427.710 ;
        RECT 1420.120 379.450 1420.380 379.770 ;
        RECT 1420.180 331.150 1420.320 379.450 ;
        RECT 1420.120 330.830 1420.380 331.150 ;
        RECT 1419.660 283.230 1419.920 283.550 ;
        RECT 1419.720 282.870 1419.860 283.230 ;
        RECT 1419.660 282.550 1419.920 282.870 ;
        RECT 1420.120 234.610 1420.380 234.930 ;
        RECT 1420.180 234.330 1420.320 234.610 ;
        RECT 1419.720 234.190 1420.320 234.330 ;
        RECT 1419.720 192.770 1419.860 234.190 ;
        RECT 1419.660 192.450 1419.920 192.770 ;
        RECT 1421.500 192.450 1421.760 192.770 ;
        RECT 1421.560 145.170 1421.700 192.450 ;
        RECT 1420.120 144.850 1420.380 145.170 ;
        RECT 1421.500 144.850 1421.760 145.170 ;
        RECT 1420.180 48.950 1420.320 144.850 ;
        RECT 1420.120 48.630 1420.380 48.950 ;
        RECT 1419.660 41.490 1419.920 41.810 ;
        RECT 1419.720 22.770 1419.860 41.490 ;
        RECT 1419.660 22.450 1419.920 22.770 ;
        RECT 1656.100 22.450 1656.360 22.770 ;
        RECT 1656.160 2.000 1656.300 22.450 ;
        RECT 1655.950 -4.000 1656.510 2.000 ;
      LAYER via2 ;
        RECT 1419.190 1007.280 1419.470 1007.560 ;
        RECT 1420.110 1007.280 1420.390 1007.560 ;
        RECT 1419.190 910.720 1419.470 911.000 ;
        RECT 1420.110 910.720 1420.390 911.000 ;
        RECT 1419.190 814.160 1419.470 814.440 ;
        RECT 1420.110 814.160 1420.390 814.440 ;
        RECT 1421.490 621.040 1421.770 621.320 ;
        RECT 1420.110 531.280 1420.390 531.560 ;
      LAYER met3 ;
        RECT 1419.165 1007.570 1419.495 1007.585 ;
        RECT 1420.085 1007.570 1420.415 1007.585 ;
        RECT 1419.165 1007.270 1420.415 1007.570 ;
        RECT 1419.165 1007.255 1419.495 1007.270 ;
        RECT 1420.085 1007.255 1420.415 1007.270 ;
        RECT 1419.165 911.010 1419.495 911.025 ;
        RECT 1420.085 911.010 1420.415 911.025 ;
        RECT 1419.165 910.710 1420.415 911.010 ;
        RECT 1419.165 910.695 1419.495 910.710 ;
        RECT 1420.085 910.695 1420.415 910.710 ;
        RECT 1419.165 814.450 1419.495 814.465 ;
        RECT 1420.085 814.450 1420.415 814.465 ;
        RECT 1419.165 814.150 1420.415 814.450 ;
        RECT 1419.165 814.135 1419.495 814.150 ;
        RECT 1420.085 814.135 1420.415 814.150 ;
        RECT 1421.465 621.330 1421.795 621.345 ;
        RECT 1420.100 621.030 1421.795 621.330 ;
        RECT 1420.100 619.980 1420.400 621.030 ;
        RECT 1421.465 621.015 1421.795 621.030 ;
        RECT 1419.830 619.670 1420.400 619.980 ;
        RECT 1419.830 619.660 1420.210 619.670 ;
        RECT 1420.085 531.580 1420.415 531.585 ;
        RECT 1419.830 531.570 1420.415 531.580 ;
        RECT 1419.830 531.270 1420.640 531.570 ;
        RECT 1419.830 531.260 1420.415 531.270 ;
        RECT 1420.085 531.255 1420.415 531.260 ;
      LAYER via3 ;
        RECT 1419.860 619.660 1420.180 619.980 ;
        RECT 1419.860 531.260 1420.180 531.580 ;
      LAYER met4 ;
        RECT 1419.855 619.655 1420.185 619.985 ;
        RECT 1419.870 531.585 1420.170 619.655 ;
        RECT 1419.855 531.255 1420.185 531.585 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1426.145 834.445 1426.315 910.775 ;
        RECT 1426.605 689.605 1426.775 717.655 ;
        RECT 1426.605 282.965 1426.775 331.075 ;
      LAYER mcon ;
        RECT 1426.145 910.605 1426.315 910.775 ;
        RECT 1426.605 717.485 1426.775 717.655 ;
        RECT 1426.605 330.905 1426.775 331.075 ;
      LAYER met1 ;
        RECT 1424.230 1062.740 1424.550 1062.800 ;
        RECT 1426.530 1062.740 1426.850 1062.800 ;
        RECT 1424.230 1062.600 1426.850 1062.740 ;
        RECT 1424.230 1062.540 1424.550 1062.600 ;
        RECT 1426.530 1062.540 1426.850 1062.600 ;
        RECT 1426.070 910.760 1426.390 910.820 ;
        RECT 1425.875 910.620 1426.390 910.760 ;
        RECT 1426.070 910.560 1426.390 910.620 ;
        RECT 1426.085 834.600 1426.375 834.645 ;
        RECT 1426.530 834.600 1426.850 834.660 ;
        RECT 1426.085 834.460 1426.850 834.600 ;
        RECT 1426.085 834.415 1426.375 834.460 ;
        RECT 1426.530 834.400 1426.850 834.460 ;
        RECT 1426.530 717.640 1426.850 717.700 ;
        RECT 1426.335 717.500 1426.850 717.640 ;
        RECT 1426.530 717.440 1426.850 717.500 ;
        RECT 1426.530 689.760 1426.850 689.820 ;
        RECT 1426.335 689.620 1426.850 689.760 ;
        RECT 1426.530 689.560 1426.850 689.620 ;
        RECT 1426.530 628.220 1426.850 628.280 ;
        RECT 1426.990 628.220 1427.310 628.280 ;
        RECT 1426.530 628.080 1427.310 628.220 ;
        RECT 1426.530 628.020 1426.850 628.080 ;
        RECT 1426.990 628.020 1427.310 628.080 ;
        RECT 1426.990 545.600 1427.310 545.660 ;
        RECT 1426.620 545.460 1427.310 545.600 ;
        RECT 1426.620 544.980 1426.760 545.460 ;
        RECT 1426.990 545.400 1427.310 545.460 ;
        RECT 1426.530 544.720 1426.850 544.980 ;
        RECT 1426.070 338.200 1426.390 338.260 ;
        RECT 1426.530 338.200 1426.850 338.260 ;
        RECT 1426.070 338.060 1426.850 338.200 ;
        RECT 1426.070 338.000 1426.390 338.060 ;
        RECT 1426.530 338.000 1426.850 338.060 ;
        RECT 1426.530 331.060 1426.850 331.120 ;
        RECT 1426.335 330.920 1426.850 331.060 ;
        RECT 1426.530 330.860 1426.850 330.920 ;
        RECT 1426.545 283.120 1426.835 283.165 ;
        RECT 1426.990 283.120 1427.310 283.180 ;
        RECT 1426.545 282.980 1427.310 283.120 ;
        RECT 1426.545 282.935 1426.835 282.980 ;
        RECT 1426.990 282.920 1427.310 282.980 ;
        RECT 1426.530 241.640 1426.850 241.700 ;
        RECT 1426.990 241.640 1427.310 241.700 ;
        RECT 1426.530 241.500 1427.310 241.640 ;
        RECT 1426.530 241.440 1426.850 241.500 ;
        RECT 1426.990 241.440 1427.310 241.500 ;
        RECT 1426.990 159.020 1427.310 159.080 ;
        RECT 1426.620 158.880 1427.310 159.020 ;
        RECT 1426.620 158.740 1426.760 158.880 ;
        RECT 1426.990 158.820 1427.310 158.880 ;
        RECT 1426.530 158.480 1426.850 158.740 ;
        RECT 1426.990 62.460 1427.310 62.520 ;
        RECT 1426.620 62.320 1427.310 62.460 ;
        RECT 1426.620 62.180 1426.760 62.320 ;
        RECT 1426.990 62.260 1427.310 62.320 ;
        RECT 1426.530 61.920 1426.850 62.180 ;
        RECT 1426.530 23.020 1426.850 23.080 ;
        RECT 1673.550 23.020 1673.870 23.080 ;
        RECT 1426.530 22.880 1673.870 23.020 ;
        RECT 1426.530 22.820 1426.850 22.880 ;
        RECT 1673.550 22.820 1673.870 22.880 ;
      LAYER via ;
        RECT 1424.260 1062.540 1424.520 1062.800 ;
        RECT 1426.560 1062.540 1426.820 1062.800 ;
        RECT 1426.100 910.560 1426.360 910.820 ;
        RECT 1426.560 834.400 1426.820 834.660 ;
        RECT 1426.560 717.440 1426.820 717.700 ;
        RECT 1426.560 689.560 1426.820 689.820 ;
        RECT 1426.560 628.020 1426.820 628.280 ;
        RECT 1427.020 628.020 1427.280 628.280 ;
        RECT 1427.020 545.400 1427.280 545.660 ;
        RECT 1426.560 544.720 1426.820 544.980 ;
        RECT 1426.100 338.000 1426.360 338.260 ;
        RECT 1426.560 338.000 1426.820 338.260 ;
        RECT 1426.560 330.860 1426.820 331.120 ;
        RECT 1427.020 282.920 1427.280 283.180 ;
        RECT 1426.560 241.440 1426.820 241.700 ;
        RECT 1427.020 241.440 1427.280 241.700 ;
        RECT 1427.020 158.820 1427.280 159.080 ;
        RECT 1426.560 158.480 1426.820 158.740 ;
        RECT 1427.020 62.260 1427.280 62.520 ;
        RECT 1426.560 61.920 1426.820 62.180 ;
        RECT 1426.560 22.820 1426.820 23.080 ;
        RECT 1673.580 22.820 1673.840 23.080 ;
      LAYER met2 ;
        RECT 1424.170 1100.580 1424.450 1104.000 ;
        RECT 1424.170 1100.000 1424.460 1100.580 ;
        RECT 1424.320 1062.830 1424.460 1100.000 ;
        RECT 1424.260 1062.510 1424.520 1062.830 ;
        RECT 1426.560 1062.570 1426.820 1062.830 ;
        RECT 1426.160 1062.510 1426.820 1062.570 ;
        RECT 1426.160 1062.430 1426.760 1062.510 ;
        RECT 1426.160 960.005 1426.300 1062.430 ;
        RECT 1426.090 959.635 1426.370 960.005 ;
        RECT 1426.550 958.955 1426.830 959.325 ;
        RECT 1426.620 917.730 1426.760 958.955 ;
        RECT 1426.160 917.590 1426.760 917.730 ;
        RECT 1426.160 910.850 1426.300 917.590 ;
        RECT 1426.100 910.530 1426.360 910.850 ;
        RECT 1426.560 834.370 1426.820 834.690 ;
        RECT 1426.620 796.690 1426.760 834.370 ;
        RECT 1426.620 796.550 1427.220 796.690 ;
        RECT 1427.080 724.610 1427.220 796.550 ;
        RECT 1426.620 724.470 1427.220 724.610 ;
        RECT 1426.620 717.730 1426.760 724.470 ;
        RECT 1426.560 717.410 1426.820 717.730 ;
        RECT 1426.560 689.530 1426.820 689.850 ;
        RECT 1426.620 669.530 1426.760 689.530 ;
        RECT 1426.620 669.390 1427.220 669.530 ;
        RECT 1427.080 628.310 1427.220 669.390 ;
        RECT 1426.560 627.990 1426.820 628.310 ;
        RECT 1427.020 627.990 1427.280 628.310 ;
        RECT 1426.620 603.570 1426.760 627.990 ;
        RECT 1426.620 603.430 1427.220 603.570 ;
        RECT 1427.080 545.690 1427.220 603.430 ;
        RECT 1427.020 545.370 1427.280 545.690 ;
        RECT 1426.560 544.690 1426.820 545.010 ;
        RECT 1426.620 507.010 1426.760 544.690 ;
        RECT 1426.620 506.870 1427.220 507.010 ;
        RECT 1427.080 449.040 1427.220 506.870 ;
        RECT 1426.620 448.900 1427.220 449.040 ;
        RECT 1426.620 403.650 1426.760 448.900 ;
        RECT 1426.160 403.510 1426.760 403.650 ;
        RECT 1426.160 338.290 1426.300 403.510 ;
        RECT 1426.100 337.970 1426.360 338.290 ;
        RECT 1426.560 337.970 1426.820 338.290 ;
        RECT 1426.620 331.150 1426.760 337.970 ;
        RECT 1426.560 330.830 1426.820 331.150 ;
        RECT 1427.020 282.890 1427.280 283.210 ;
        RECT 1427.080 241.730 1427.220 282.890 ;
        RECT 1426.560 241.410 1426.820 241.730 ;
        RECT 1427.020 241.410 1427.280 241.730 ;
        RECT 1426.620 217.330 1426.760 241.410 ;
        RECT 1426.620 217.190 1427.220 217.330 ;
        RECT 1427.080 159.110 1427.220 217.190 ;
        RECT 1427.020 158.790 1427.280 159.110 ;
        RECT 1426.560 158.450 1426.820 158.770 ;
        RECT 1426.620 131.650 1426.760 158.450 ;
        RECT 1426.620 131.510 1427.220 131.650 ;
        RECT 1427.080 62.550 1427.220 131.510 ;
        RECT 1427.020 62.230 1427.280 62.550 ;
        RECT 1426.560 61.890 1426.820 62.210 ;
        RECT 1426.620 23.110 1426.760 61.890 ;
        RECT 1426.560 22.790 1426.820 23.110 ;
        RECT 1673.580 22.790 1673.840 23.110 ;
        RECT 1673.640 2.000 1673.780 22.790 ;
        RECT 1673.430 -4.000 1673.990 2.000 ;
      LAYER via2 ;
        RECT 1426.090 959.680 1426.370 959.960 ;
        RECT 1426.550 959.000 1426.830 959.280 ;
      LAYER met3 ;
        RECT 1426.065 959.970 1426.395 959.985 ;
        RECT 1426.065 959.655 1426.610 959.970 ;
        RECT 1426.310 959.305 1426.610 959.655 ;
        RECT 1426.310 958.990 1426.855 959.305 ;
        RECT 1426.525 958.975 1426.855 958.990 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1433.505 766.105 1433.675 814.215 ;
        RECT 1433.045 689.605 1433.215 717.655 ;
        RECT 1433.045 282.965 1433.215 331.075 ;
      LAYER mcon ;
        RECT 1433.505 814.045 1433.675 814.215 ;
        RECT 1433.045 717.485 1433.215 717.655 ;
        RECT 1433.045 330.905 1433.215 331.075 ;
      LAYER met1 ;
        RECT 1430.670 1062.740 1430.990 1062.800 ;
        RECT 1432.970 1062.740 1433.290 1062.800 ;
        RECT 1430.670 1062.600 1433.290 1062.740 ;
        RECT 1430.670 1062.540 1430.990 1062.600 ;
        RECT 1432.970 1062.540 1433.290 1062.600 ;
        RECT 1432.970 1028.200 1433.290 1028.460 ;
        RECT 1433.060 1027.720 1433.200 1028.200 ;
        RECT 1433.430 1027.720 1433.750 1027.780 ;
        RECT 1433.060 1027.580 1433.750 1027.720 ;
        RECT 1433.430 1027.520 1433.750 1027.580 ;
        RECT 1432.510 966.180 1432.830 966.240 ;
        RECT 1433.430 966.180 1433.750 966.240 ;
        RECT 1432.510 966.040 1433.750 966.180 ;
        RECT 1432.510 965.980 1432.830 966.040 ;
        RECT 1433.430 965.980 1433.750 966.040 ;
        RECT 1433.430 918.240 1433.750 918.300 ;
        RECT 1433.060 918.100 1433.750 918.240 ;
        RECT 1433.060 917.960 1433.200 918.100 ;
        RECT 1433.430 918.040 1433.750 918.100 ;
        RECT 1432.970 917.700 1433.290 917.960 ;
        RECT 1432.510 869.420 1432.830 869.680 ;
        RECT 1432.600 868.940 1432.740 869.420 ;
        RECT 1432.970 868.940 1433.290 869.000 ;
        RECT 1432.600 868.800 1433.290 868.940 ;
        RECT 1432.970 868.740 1433.290 868.800 ;
        RECT 1432.970 821.000 1433.290 821.060 ;
        RECT 1433.430 821.000 1433.750 821.060 ;
        RECT 1432.970 820.860 1433.750 821.000 ;
        RECT 1432.970 820.800 1433.290 820.860 ;
        RECT 1433.430 820.800 1433.750 820.860 ;
        RECT 1433.430 814.200 1433.750 814.260 ;
        RECT 1433.235 814.060 1433.750 814.200 ;
        RECT 1433.430 814.000 1433.750 814.060 ;
        RECT 1433.430 766.260 1433.750 766.320 ;
        RECT 1433.235 766.120 1433.750 766.260 ;
        RECT 1433.430 766.060 1433.750 766.120 ;
        RECT 1432.970 717.640 1433.290 717.700 ;
        RECT 1432.775 717.500 1433.290 717.640 ;
        RECT 1432.970 717.440 1433.290 717.500 ;
        RECT 1432.970 689.760 1433.290 689.820 ;
        RECT 1432.775 689.620 1433.290 689.760 ;
        RECT 1432.970 689.560 1433.290 689.620 ;
        RECT 1432.970 628.220 1433.290 628.280 ;
        RECT 1433.430 628.220 1433.750 628.280 ;
        RECT 1432.970 628.080 1433.750 628.220 ;
        RECT 1432.970 628.020 1433.290 628.080 ;
        RECT 1433.430 628.020 1433.750 628.080 ;
        RECT 1432.050 579.600 1432.370 579.660 ;
        RECT 1433.430 579.600 1433.750 579.660 ;
        RECT 1432.050 579.460 1433.750 579.600 ;
        RECT 1432.050 579.400 1432.370 579.460 ;
        RECT 1433.430 579.400 1433.750 579.460 ;
        RECT 1432.510 338.200 1432.830 338.260 ;
        RECT 1432.970 338.200 1433.290 338.260 ;
        RECT 1432.510 338.060 1433.290 338.200 ;
        RECT 1432.510 338.000 1432.830 338.060 ;
        RECT 1432.970 338.000 1433.290 338.060 ;
        RECT 1432.970 331.060 1433.290 331.120 ;
        RECT 1432.775 330.920 1433.290 331.060 ;
        RECT 1432.970 330.860 1433.290 330.920 ;
        RECT 1432.985 283.120 1433.275 283.165 ;
        RECT 1433.430 283.120 1433.750 283.180 ;
        RECT 1432.985 282.980 1433.750 283.120 ;
        RECT 1432.985 282.935 1433.275 282.980 ;
        RECT 1433.430 282.920 1433.750 282.980 ;
        RECT 1432.970 241.640 1433.290 241.700 ;
        RECT 1433.430 241.640 1433.750 241.700 ;
        RECT 1432.970 241.500 1433.750 241.640 ;
        RECT 1432.970 241.440 1433.290 241.500 ;
        RECT 1433.430 241.440 1433.750 241.500 ;
        RECT 1433.430 159.020 1433.750 159.080 ;
        RECT 1433.060 158.880 1433.750 159.020 ;
        RECT 1433.060 158.740 1433.200 158.880 ;
        RECT 1433.430 158.820 1433.750 158.880 ;
        RECT 1432.970 158.480 1433.290 158.740 ;
        RECT 1433.430 62.460 1433.750 62.520 ;
        RECT 1433.060 62.320 1433.750 62.460 ;
        RECT 1433.060 62.180 1433.200 62.320 ;
        RECT 1433.430 62.260 1433.750 62.320 ;
        RECT 1432.970 61.920 1433.290 62.180 ;
        RECT 1432.970 23.700 1433.290 23.760 ;
        RECT 1691.490 23.700 1691.810 23.760 ;
        RECT 1432.970 23.560 1691.810 23.700 ;
        RECT 1432.970 23.500 1433.290 23.560 ;
        RECT 1691.490 23.500 1691.810 23.560 ;
      LAYER via ;
        RECT 1430.700 1062.540 1430.960 1062.800 ;
        RECT 1433.000 1062.540 1433.260 1062.800 ;
        RECT 1433.000 1028.200 1433.260 1028.460 ;
        RECT 1433.460 1027.520 1433.720 1027.780 ;
        RECT 1432.540 965.980 1432.800 966.240 ;
        RECT 1433.460 965.980 1433.720 966.240 ;
        RECT 1433.460 918.040 1433.720 918.300 ;
        RECT 1433.000 917.700 1433.260 917.960 ;
        RECT 1432.540 869.420 1432.800 869.680 ;
        RECT 1433.000 868.740 1433.260 869.000 ;
        RECT 1433.000 820.800 1433.260 821.060 ;
        RECT 1433.460 820.800 1433.720 821.060 ;
        RECT 1433.460 814.000 1433.720 814.260 ;
        RECT 1433.460 766.060 1433.720 766.320 ;
        RECT 1433.000 717.440 1433.260 717.700 ;
        RECT 1433.000 689.560 1433.260 689.820 ;
        RECT 1433.000 628.020 1433.260 628.280 ;
        RECT 1433.460 628.020 1433.720 628.280 ;
        RECT 1432.080 579.400 1432.340 579.660 ;
        RECT 1433.460 579.400 1433.720 579.660 ;
        RECT 1432.540 338.000 1432.800 338.260 ;
        RECT 1433.000 338.000 1433.260 338.260 ;
        RECT 1433.000 330.860 1433.260 331.120 ;
        RECT 1433.460 282.920 1433.720 283.180 ;
        RECT 1433.000 241.440 1433.260 241.700 ;
        RECT 1433.460 241.440 1433.720 241.700 ;
        RECT 1433.460 158.820 1433.720 159.080 ;
        RECT 1433.000 158.480 1433.260 158.740 ;
        RECT 1433.460 62.260 1433.720 62.520 ;
        RECT 1433.000 61.920 1433.260 62.180 ;
        RECT 1433.000 23.500 1433.260 23.760 ;
        RECT 1691.520 23.500 1691.780 23.760 ;
      LAYER met2 ;
        RECT 1430.610 1100.580 1430.890 1104.000 ;
        RECT 1430.610 1100.000 1430.900 1100.580 ;
        RECT 1430.760 1062.830 1430.900 1100.000 ;
        RECT 1430.700 1062.510 1430.960 1062.830 ;
        RECT 1433.000 1062.510 1433.260 1062.830 ;
        RECT 1433.060 1028.490 1433.200 1062.510 ;
        RECT 1433.000 1028.170 1433.260 1028.490 ;
        RECT 1433.460 1027.490 1433.720 1027.810 ;
        RECT 1433.520 1014.405 1433.660 1027.490 ;
        RECT 1432.530 1014.035 1432.810 1014.405 ;
        RECT 1433.450 1014.035 1433.730 1014.405 ;
        RECT 1432.600 966.270 1432.740 1014.035 ;
        RECT 1432.540 965.950 1432.800 966.270 ;
        RECT 1433.460 965.950 1433.720 966.270 ;
        RECT 1433.520 918.330 1433.660 965.950 ;
        RECT 1433.460 918.010 1433.720 918.330 ;
        RECT 1433.000 917.845 1433.260 917.990 ;
        RECT 1432.990 917.475 1433.270 917.845 ;
        RECT 1432.530 916.795 1432.810 917.165 ;
        RECT 1432.600 869.710 1432.740 916.795 ;
        RECT 1432.540 869.390 1432.800 869.710 ;
        RECT 1433.000 868.710 1433.260 869.030 ;
        RECT 1433.060 821.090 1433.200 868.710 ;
        RECT 1433.000 820.770 1433.260 821.090 ;
        RECT 1433.460 820.770 1433.720 821.090 ;
        RECT 1433.520 814.290 1433.660 820.770 ;
        RECT 1433.460 813.970 1433.720 814.290 ;
        RECT 1433.460 766.030 1433.720 766.350 ;
        RECT 1433.520 724.610 1433.660 766.030 ;
        RECT 1433.060 724.470 1433.660 724.610 ;
        RECT 1433.060 717.730 1433.200 724.470 ;
        RECT 1433.000 717.410 1433.260 717.730 ;
        RECT 1433.000 689.530 1433.260 689.850 ;
        RECT 1433.060 669.530 1433.200 689.530 ;
        RECT 1433.060 669.390 1433.660 669.530 ;
        RECT 1433.520 628.310 1433.660 669.390 ;
        RECT 1433.000 627.990 1433.260 628.310 ;
        RECT 1433.460 627.990 1433.720 628.310 ;
        RECT 1433.060 603.570 1433.200 627.990 ;
        RECT 1433.060 603.430 1433.660 603.570 ;
        RECT 1433.520 579.690 1433.660 603.430 ;
        RECT 1432.080 579.370 1432.340 579.690 ;
        RECT 1433.460 579.370 1433.720 579.690 ;
        RECT 1432.140 531.605 1432.280 579.370 ;
        RECT 1432.070 531.235 1432.350 531.605 ;
        RECT 1432.990 531.235 1433.270 531.605 ;
        RECT 1433.060 507.010 1433.200 531.235 ;
        RECT 1433.060 506.870 1433.660 507.010 ;
        RECT 1433.520 449.040 1433.660 506.870 ;
        RECT 1433.060 448.900 1433.660 449.040 ;
        RECT 1433.060 403.650 1433.200 448.900 ;
        RECT 1432.600 403.510 1433.200 403.650 ;
        RECT 1432.600 338.290 1432.740 403.510 ;
        RECT 1432.540 337.970 1432.800 338.290 ;
        RECT 1433.000 337.970 1433.260 338.290 ;
        RECT 1433.060 331.150 1433.200 337.970 ;
        RECT 1433.000 330.830 1433.260 331.150 ;
        RECT 1433.460 282.890 1433.720 283.210 ;
        RECT 1433.520 241.730 1433.660 282.890 ;
        RECT 1433.000 241.410 1433.260 241.730 ;
        RECT 1433.460 241.410 1433.720 241.730 ;
        RECT 1433.060 217.330 1433.200 241.410 ;
        RECT 1433.060 217.190 1433.660 217.330 ;
        RECT 1433.520 159.110 1433.660 217.190 ;
        RECT 1433.460 158.790 1433.720 159.110 ;
        RECT 1433.000 158.450 1433.260 158.770 ;
        RECT 1433.060 131.650 1433.200 158.450 ;
        RECT 1433.060 131.510 1433.660 131.650 ;
        RECT 1433.520 62.550 1433.660 131.510 ;
        RECT 1433.460 62.230 1433.720 62.550 ;
        RECT 1433.000 61.890 1433.260 62.210 ;
        RECT 1433.060 23.790 1433.200 61.890 ;
        RECT 1433.000 23.470 1433.260 23.790 ;
        RECT 1691.520 23.470 1691.780 23.790 ;
        RECT 1691.580 2.000 1691.720 23.470 ;
        RECT 1691.370 -4.000 1691.930 2.000 ;
      LAYER via2 ;
        RECT 1432.530 1014.080 1432.810 1014.360 ;
        RECT 1433.450 1014.080 1433.730 1014.360 ;
        RECT 1432.990 917.520 1433.270 917.800 ;
        RECT 1432.530 916.840 1432.810 917.120 ;
        RECT 1432.070 531.280 1432.350 531.560 ;
        RECT 1432.990 531.280 1433.270 531.560 ;
      LAYER met3 ;
        RECT 1432.505 1014.370 1432.835 1014.385 ;
        RECT 1433.425 1014.370 1433.755 1014.385 ;
        RECT 1432.505 1014.070 1433.755 1014.370 ;
        RECT 1432.505 1014.055 1432.835 1014.070 ;
        RECT 1433.425 1014.055 1433.755 1014.070 ;
        RECT 1432.965 917.810 1433.295 917.825 ;
        RECT 1432.750 917.495 1433.295 917.810 ;
        RECT 1432.750 917.145 1433.050 917.495 ;
        RECT 1432.505 916.830 1433.050 917.145 ;
        RECT 1432.505 916.815 1432.835 916.830 ;
        RECT 1432.045 531.570 1432.375 531.585 ;
        RECT 1432.965 531.570 1433.295 531.585 ;
        RECT 1432.045 531.270 1433.295 531.570 ;
        RECT 1432.045 531.255 1432.375 531.270 ;
        RECT 1432.965 531.255 1433.295 531.270 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 728.250 43.760 728.570 43.820 ;
        RECT 1098.090 43.760 1098.410 43.820 ;
        RECT 728.250 43.620 1098.410 43.760 ;
        RECT 728.250 43.560 728.570 43.620 ;
        RECT 1098.090 43.560 1098.410 43.620 ;
      LAYER via ;
        RECT 728.280 43.560 728.540 43.820 ;
        RECT 1098.120 43.560 1098.380 43.820 ;
      LAYER met2 ;
        RECT 1099.870 1100.650 1100.150 1104.000 ;
        RECT 1098.180 1100.510 1100.150 1100.650 ;
        RECT 1098.180 43.850 1098.320 1100.510 ;
        RECT 1099.870 1100.000 1100.150 1100.510 ;
        RECT 728.280 43.530 728.540 43.850 ;
        RECT 1098.120 43.530 1098.380 43.850 ;
        RECT 728.340 2.000 728.480 43.530 ;
        RECT 728.130 -4.000 728.690 2.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1436.650 1085.180 1436.970 1085.240 ;
        RECT 1441.250 1085.180 1441.570 1085.240 ;
        RECT 1436.650 1085.040 1441.570 1085.180 ;
        RECT 1436.650 1084.980 1436.970 1085.040 ;
        RECT 1441.250 1084.980 1441.570 1085.040 ;
        RECT 1441.250 27.440 1441.570 27.500 ;
        RECT 1709.430 27.440 1709.750 27.500 ;
        RECT 1441.250 27.300 1709.750 27.440 ;
        RECT 1441.250 27.240 1441.570 27.300 ;
        RECT 1709.430 27.240 1709.750 27.300 ;
      LAYER via ;
        RECT 1436.680 1084.980 1436.940 1085.240 ;
        RECT 1441.280 1084.980 1441.540 1085.240 ;
        RECT 1441.280 27.240 1441.540 27.500 ;
        RECT 1709.460 27.240 1709.720 27.500 ;
      LAYER met2 ;
        RECT 1436.590 1100.580 1436.870 1104.000 ;
        RECT 1436.590 1100.000 1436.880 1100.580 ;
        RECT 1436.740 1085.270 1436.880 1100.000 ;
        RECT 1436.680 1084.950 1436.940 1085.270 ;
        RECT 1441.280 1084.950 1441.540 1085.270 ;
        RECT 1441.340 27.530 1441.480 1084.950 ;
        RECT 1441.280 27.210 1441.540 27.530 ;
        RECT 1709.460 27.210 1709.720 27.530 ;
        RECT 1709.520 2.000 1709.660 27.210 ;
        RECT 1709.310 -4.000 1709.870 2.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1442.630 1086.540 1442.950 1086.600 ;
        RECT 1448.150 1086.540 1448.470 1086.600 ;
        RECT 1442.630 1086.400 1448.470 1086.540 ;
        RECT 1442.630 1086.340 1442.950 1086.400 ;
        RECT 1448.150 1086.340 1448.470 1086.400 ;
        RECT 1448.150 26.760 1448.470 26.820 ;
        RECT 1727.370 26.760 1727.690 26.820 ;
        RECT 1448.150 26.620 1727.690 26.760 ;
        RECT 1448.150 26.560 1448.470 26.620 ;
        RECT 1727.370 26.560 1727.690 26.620 ;
      LAYER via ;
        RECT 1442.660 1086.340 1442.920 1086.600 ;
        RECT 1448.180 1086.340 1448.440 1086.600 ;
        RECT 1448.180 26.560 1448.440 26.820 ;
        RECT 1727.400 26.560 1727.660 26.820 ;
      LAYER met2 ;
        RECT 1442.570 1100.580 1442.850 1104.000 ;
        RECT 1442.570 1100.000 1442.860 1100.580 ;
        RECT 1442.720 1086.630 1442.860 1100.000 ;
        RECT 1442.660 1086.310 1442.920 1086.630 ;
        RECT 1448.180 1086.310 1448.440 1086.630 ;
        RECT 1448.240 26.850 1448.380 1086.310 ;
        RECT 1448.180 26.530 1448.440 26.850 ;
        RECT 1727.400 26.530 1727.660 26.850 ;
        RECT 1727.460 2.000 1727.600 26.530 ;
        RECT 1727.250 -4.000 1727.810 2.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1447.690 40.020 1448.010 40.080 ;
        RECT 1745.310 40.020 1745.630 40.080 ;
        RECT 1447.690 39.880 1745.630 40.020 ;
        RECT 1447.690 39.820 1448.010 39.880 ;
        RECT 1745.310 39.820 1745.630 39.880 ;
      LAYER via ;
        RECT 1447.720 39.820 1447.980 40.080 ;
        RECT 1745.340 39.820 1745.600 40.080 ;
      LAYER met2 ;
        RECT 1448.550 1100.650 1448.830 1104.000 ;
        RECT 1447.780 1100.510 1448.830 1100.650 ;
        RECT 1447.780 40.110 1447.920 1100.510 ;
        RECT 1448.550 1100.000 1448.830 1100.510 ;
        RECT 1447.720 39.790 1447.980 40.110 ;
        RECT 1745.340 39.790 1745.600 40.110 ;
        RECT 1745.400 2.000 1745.540 39.790 ;
        RECT 1745.190 -4.000 1745.750 2.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1454.590 39.680 1454.910 39.740 ;
        RECT 1762.790 39.680 1763.110 39.740 ;
        RECT 1454.590 39.540 1763.110 39.680 ;
        RECT 1454.590 39.480 1454.910 39.540 ;
        RECT 1762.790 39.480 1763.110 39.540 ;
      LAYER via ;
        RECT 1454.620 39.480 1454.880 39.740 ;
        RECT 1762.820 39.480 1763.080 39.740 ;
      LAYER met2 ;
        RECT 1454.990 1100.650 1455.270 1104.000 ;
        RECT 1454.680 1100.510 1455.270 1100.650 ;
        RECT 1454.680 39.770 1454.820 1100.510 ;
        RECT 1454.990 1100.000 1455.270 1100.510 ;
        RECT 1454.620 39.450 1454.880 39.770 ;
        RECT 1762.820 39.450 1763.080 39.770 ;
        RECT 1762.880 2.000 1763.020 39.450 ;
        RECT 1762.670 -4.000 1763.230 2.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1461.490 39.340 1461.810 39.400 ;
        RECT 1780.730 39.340 1781.050 39.400 ;
        RECT 1461.490 39.200 1781.050 39.340 ;
        RECT 1461.490 39.140 1461.810 39.200 ;
        RECT 1780.730 39.140 1781.050 39.200 ;
      LAYER via ;
        RECT 1461.520 39.140 1461.780 39.400 ;
        RECT 1780.760 39.140 1781.020 39.400 ;
      LAYER met2 ;
        RECT 1460.970 1100.650 1461.250 1104.000 ;
        RECT 1460.970 1100.510 1461.720 1100.650 ;
        RECT 1460.970 1100.000 1461.250 1100.510 ;
        RECT 1461.580 39.430 1461.720 1100.510 ;
        RECT 1461.520 39.110 1461.780 39.430 ;
        RECT 1780.760 39.110 1781.020 39.430 ;
        RECT 1780.820 2.000 1780.960 39.110 ;
        RECT 1780.610 -4.000 1781.170 2.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1468.390 39.000 1468.710 39.060 ;
        RECT 1798.670 39.000 1798.990 39.060 ;
        RECT 1468.390 38.860 1798.990 39.000 ;
        RECT 1468.390 38.800 1468.710 38.860 ;
        RECT 1798.670 38.800 1798.990 38.860 ;
      LAYER via ;
        RECT 1468.420 38.800 1468.680 39.060 ;
        RECT 1798.700 38.800 1798.960 39.060 ;
      LAYER met2 ;
        RECT 1466.950 1100.650 1467.230 1104.000 ;
        RECT 1466.950 1100.510 1468.620 1100.650 ;
        RECT 1466.950 1100.000 1467.230 1100.510 ;
        RECT 1468.480 39.090 1468.620 1100.510 ;
        RECT 1468.420 38.770 1468.680 39.090 ;
        RECT 1798.700 38.770 1798.960 39.090 ;
        RECT 1798.760 2.000 1798.900 38.770 ;
        RECT 1798.550 -4.000 1799.110 2.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1473.450 1062.740 1473.770 1062.800 ;
        RECT 1475.290 1062.740 1475.610 1062.800 ;
        RECT 1473.450 1062.600 1475.610 1062.740 ;
        RECT 1473.450 1062.540 1473.770 1062.600 ;
        RECT 1475.290 1062.540 1475.610 1062.600 ;
        RECT 1474.830 38.660 1475.150 38.720 ;
        RECT 1816.610 38.660 1816.930 38.720 ;
        RECT 1474.830 38.520 1816.930 38.660 ;
        RECT 1474.830 38.460 1475.150 38.520 ;
        RECT 1816.610 38.460 1816.930 38.520 ;
      LAYER via ;
        RECT 1473.480 1062.540 1473.740 1062.800 ;
        RECT 1475.320 1062.540 1475.580 1062.800 ;
        RECT 1474.860 38.460 1475.120 38.720 ;
        RECT 1816.640 38.460 1816.900 38.720 ;
      LAYER met2 ;
        RECT 1473.390 1100.580 1473.670 1104.000 ;
        RECT 1473.390 1100.000 1473.680 1100.580 ;
        RECT 1473.540 1062.830 1473.680 1100.000 ;
        RECT 1473.480 1062.510 1473.740 1062.830 ;
        RECT 1475.320 1062.510 1475.580 1062.830 ;
        RECT 1475.380 980.290 1475.520 1062.510 ;
        RECT 1474.920 980.150 1475.520 980.290 ;
        RECT 1474.920 979.610 1475.060 980.150 ;
        RECT 1474.920 979.470 1475.520 979.610 ;
        RECT 1475.380 835.450 1475.520 979.470 ;
        RECT 1474.920 835.310 1475.520 835.450 ;
        RECT 1474.920 834.770 1475.060 835.310 ;
        RECT 1474.920 834.630 1475.520 834.770 ;
        RECT 1475.380 738.890 1475.520 834.630 ;
        RECT 1474.920 738.750 1475.520 738.890 ;
        RECT 1474.920 738.210 1475.060 738.750 ;
        RECT 1474.920 738.070 1475.520 738.210 ;
        RECT 1475.380 642.330 1475.520 738.070 ;
        RECT 1474.920 642.190 1475.520 642.330 ;
        RECT 1474.920 641.650 1475.060 642.190 ;
        RECT 1474.920 641.510 1475.520 641.650 ;
        RECT 1475.380 545.770 1475.520 641.510 ;
        RECT 1474.920 545.630 1475.520 545.770 ;
        RECT 1474.920 545.090 1475.060 545.630 ;
        RECT 1474.920 544.950 1475.520 545.090 ;
        RECT 1475.380 449.210 1475.520 544.950 ;
        RECT 1474.920 449.070 1475.520 449.210 ;
        RECT 1474.920 448.530 1475.060 449.070 ;
        RECT 1474.920 448.390 1475.520 448.530 ;
        RECT 1475.380 351.970 1475.520 448.390 ;
        RECT 1474.920 351.830 1475.520 351.970 ;
        RECT 1474.920 351.290 1475.060 351.830 ;
        RECT 1474.920 351.150 1475.520 351.290 ;
        RECT 1475.380 255.410 1475.520 351.150 ;
        RECT 1474.920 255.270 1475.520 255.410 ;
        RECT 1474.920 254.730 1475.060 255.270 ;
        RECT 1474.920 254.590 1475.520 254.730 ;
        RECT 1475.380 158.850 1475.520 254.590 ;
        RECT 1474.920 158.710 1475.520 158.850 ;
        RECT 1474.920 158.170 1475.060 158.710 ;
        RECT 1474.920 158.030 1475.520 158.170 ;
        RECT 1475.380 62.290 1475.520 158.030 ;
        RECT 1474.920 62.150 1475.520 62.290 ;
        RECT 1474.920 38.750 1475.060 62.150 ;
        RECT 1474.860 38.430 1475.120 38.750 ;
        RECT 1816.640 38.430 1816.900 38.750 ;
        RECT 1816.700 2.000 1816.840 38.430 ;
        RECT 1816.490 -4.000 1817.050 2.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1479.430 1088.580 1479.750 1088.640 ;
        RECT 1482.650 1088.580 1482.970 1088.640 ;
        RECT 1479.430 1088.440 1482.970 1088.580 ;
        RECT 1479.430 1088.380 1479.750 1088.440 ;
        RECT 1482.650 1088.380 1482.970 1088.440 ;
        RECT 1482.650 38.320 1482.970 38.380 ;
        RECT 1834.550 38.320 1834.870 38.380 ;
        RECT 1482.650 38.180 1834.870 38.320 ;
        RECT 1482.650 38.120 1482.970 38.180 ;
        RECT 1834.550 38.120 1834.870 38.180 ;
      LAYER via ;
        RECT 1479.460 1088.380 1479.720 1088.640 ;
        RECT 1482.680 1088.380 1482.940 1088.640 ;
        RECT 1482.680 38.120 1482.940 38.380 ;
        RECT 1834.580 38.120 1834.840 38.380 ;
      LAYER met2 ;
        RECT 1479.370 1100.580 1479.650 1104.000 ;
        RECT 1479.370 1100.000 1479.660 1100.580 ;
        RECT 1479.520 1088.670 1479.660 1100.000 ;
        RECT 1479.460 1088.350 1479.720 1088.670 ;
        RECT 1482.680 1088.350 1482.940 1088.670 ;
        RECT 1482.740 38.410 1482.880 1088.350 ;
        RECT 1482.680 38.090 1482.940 38.410 ;
        RECT 1834.580 38.090 1834.840 38.410 ;
        RECT 1834.640 2.000 1834.780 38.090 ;
        RECT 1834.430 -4.000 1834.990 2.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1485.410 1085.860 1485.730 1085.920 ;
        RECT 1489.090 1085.860 1489.410 1085.920 ;
        RECT 1485.410 1085.720 1489.410 1085.860 ;
        RECT 1485.410 1085.660 1485.730 1085.720 ;
        RECT 1489.090 1085.660 1489.410 1085.720 ;
        RECT 1489.090 56.340 1489.410 56.400 ;
        RECT 1849.270 56.340 1849.590 56.400 ;
        RECT 1489.090 56.200 1849.590 56.340 ;
        RECT 1489.090 56.140 1489.410 56.200 ;
        RECT 1849.270 56.140 1849.590 56.200 ;
      LAYER via ;
        RECT 1485.440 1085.660 1485.700 1085.920 ;
        RECT 1489.120 1085.660 1489.380 1085.920 ;
        RECT 1489.120 56.140 1489.380 56.400 ;
        RECT 1849.300 56.140 1849.560 56.400 ;
      LAYER met2 ;
        RECT 1485.350 1100.580 1485.630 1104.000 ;
        RECT 1485.350 1100.000 1485.640 1100.580 ;
        RECT 1485.500 1085.950 1485.640 1100.000 ;
        RECT 1485.440 1085.630 1485.700 1085.950 ;
        RECT 1489.120 1085.630 1489.380 1085.950 ;
        RECT 1489.180 56.430 1489.320 1085.630 ;
        RECT 1489.120 56.110 1489.380 56.430 ;
        RECT 1849.300 56.110 1849.560 56.430 ;
        RECT 1849.360 2.450 1849.500 56.110 ;
        RECT 1849.360 2.310 1852.260 2.450 ;
        RECT 1852.120 2.000 1852.260 2.310 ;
        RECT 1851.910 -4.000 1852.470 2.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1491.850 1085.520 1492.170 1085.580 ;
        RECT 1496.450 1085.520 1496.770 1085.580 ;
        RECT 1491.850 1085.380 1496.770 1085.520 ;
        RECT 1491.850 1085.320 1492.170 1085.380 ;
        RECT 1496.450 1085.320 1496.770 1085.380 ;
        RECT 1496.450 56.680 1496.770 56.740 ;
        RECT 1870.430 56.680 1870.750 56.740 ;
        RECT 1496.450 56.540 1870.750 56.680 ;
        RECT 1496.450 56.480 1496.770 56.540 ;
        RECT 1870.430 56.480 1870.750 56.540 ;
      LAYER via ;
        RECT 1491.880 1085.320 1492.140 1085.580 ;
        RECT 1496.480 1085.320 1496.740 1085.580 ;
        RECT 1496.480 56.480 1496.740 56.740 ;
        RECT 1870.460 56.480 1870.720 56.740 ;
      LAYER met2 ;
        RECT 1491.790 1100.580 1492.070 1104.000 ;
        RECT 1491.790 1100.000 1492.080 1100.580 ;
        RECT 1491.940 1085.610 1492.080 1100.000 ;
        RECT 1491.880 1085.290 1492.140 1085.610 ;
        RECT 1496.480 1085.290 1496.740 1085.610 ;
        RECT 1496.540 56.770 1496.680 1085.290 ;
        RECT 1496.480 56.450 1496.740 56.770 ;
        RECT 1870.460 56.450 1870.720 56.770 ;
        RECT 1870.520 7.890 1870.660 56.450 ;
        RECT 1870.060 7.750 1870.660 7.890 ;
        RECT 1870.060 2.000 1870.200 7.750 ;
        RECT 1869.850 -4.000 1870.410 2.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 751.710 50.220 752.030 50.280 ;
        RECT 1105.450 50.220 1105.770 50.280 ;
        RECT 751.710 50.080 1105.770 50.220 ;
        RECT 751.710 50.020 752.030 50.080 ;
        RECT 1105.450 50.020 1105.770 50.080 ;
      LAYER via ;
        RECT 751.740 50.020 752.000 50.280 ;
        RECT 1105.480 50.020 1105.740 50.280 ;
      LAYER met2 ;
        RECT 1105.850 1100.650 1106.130 1104.000 ;
        RECT 1105.540 1100.510 1106.130 1100.650 ;
        RECT 1105.540 50.310 1105.680 1100.510 ;
        RECT 1105.850 1100.000 1106.130 1100.510 ;
        RECT 751.740 49.990 752.000 50.310 ;
        RECT 1105.480 49.990 1105.740 50.310 ;
        RECT 751.800 16.730 751.940 49.990 ;
        RECT 746.280 16.590 751.940 16.730 ;
        RECT 746.280 2.000 746.420 16.590 ;
        RECT 746.070 -4.000 746.630 2.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1497.830 1088.240 1498.150 1088.300 ;
        RECT 1502.890 1088.240 1503.210 1088.300 ;
        RECT 1497.830 1088.100 1503.210 1088.240 ;
        RECT 1497.830 1088.040 1498.150 1088.100 ;
        RECT 1502.890 1088.040 1503.210 1088.100 ;
        RECT 1502.890 57.020 1503.210 57.080 ;
        RECT 1883.770 57.020 1884.090 57.080 ;
        RECT 1502.890 56.880 1884.090 57.020 ;
        RECT 1502.890 56.820 1503.210 56.880 ;
        RECT 1883.770 56.820 1884.090 56.880 ;
        RECT 1883.770 2.620 1884.090 2.680 ;
        RECT 1887.910 2.620 1888.230 2.680 ;
        RECT 1883.770 2.480 1888.230 2.620 ;
        RECT 1883.770 2.420 1884.090 2.480 ;
        RECT 1887.910 2.420 1888.230 2.480 ;
      LAYER via ;
        RECT 1497.860 1088.040 1498.120 1088.300 ;
        RECT 1502.920 1088.040 1503.180 1088.300 ;
        RECT 1502.920 56.820 1503.180 57.080 ;
        RECT 1883.800 56.820 1884.060 57.080 ;
        RECT 1883.800 2.420 1884.060 2.680 ;
        RECT 1887.940 2.420 1888.200 2.680 ;
      LAYER met2 ;
        RECT 1497.770 1100.580 1498.050 1104.000 ;
        RECT 1497.770 1100.000 1498.060 1100.580 ;
        RECT 1497.920 1088.330 1498.060 1100.000 ;
        RECT 1497.860 1088.010 1498.120 1088.330 ;
        RECT 1502.920 1088.010 1503.180 1088.330 ;
        RECT 1502.980 57.110 1503.120 1088.010 ;
        RECT 1502.920 56.790 1503.180 57.110 ;
        RECT 1883.800 56.790 1884.060 57.110 ;
        RECT 1883.860 2.710 1884.000 56.790 ;
        RECT 1883.800 2.390 1884.060 2.710 ;
        RECT 1887.940 2.390 1888.200 2.710 ;
        RECT 1888.000 2.000 1888.140 2.390 ;
        RECT 1887.790 -4.000 1888.350 2.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1503.350 57.360 1503.670 57.420 ;
        RECT 1904.470 57.360 1904.790 57.420 ;
        RECT 1503.350 57.220 1904.790 57.360 ;
        RECT 1503.350 57.160 1503.670 57.220 ;
        RECT 1904.470 57.160 1904.790 57.220 ;
      LAYER via ;
        RECT 1503.380 57.160 1503.640 57.420 ;
        RECT 1904.500 57.160 1904.760 57.420 ;
      LAYER met2 ;
        RECT 1503.750 1100.650 1504.030 1104.000 ;
        RECT 1503.440 1100.510 1504.030 1100.650 ;
        RECT 1503.440 57.450 1503.580 1100.510 ;
        RECT 1503.750 1100.000 1504.030 1100.510 ;
        RECT 1503.380 57.130 1503.640 57.450 ;
        RECT 1904.500 57.130 1904.760 57.450 ;
        RECT 1904.560 2.450 1904.700 57.130 ;
        RECT 1904.560 2.310 1906.080 2.450 ;
        RECT 1905.940 2.000 1906.080 2.310 ;
        RECT 1905.730 -4.000 1906.290 2.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1510.250 57.700 1510.570 57.760 ;
        RECT 1918.270 57.700 1918.590 57.760 ;
        RECT 1510.250 57.560 1918.590 57.700 ;
        RECT 1510.250 57.500 1510.570 57.560 ;
        RECT 1918.270 57.500 1918.590 57.560 ;
        RECT 1918.270 2.620 1918.590 2.680 ;
        RECT 1923.330 2.620 1923.650 2.680 ;
        RECT 1918.270 2.480 1923.650 2.620 ;
        RECT 1918.270 2.420 1918.590 2.480 ;
        RECT 1923.330 2.420 1923.650 2.480 ;
      LAYER via ;
        RECT 1510.280 57.500 1510.540 57.760 ;
        RECT 1918.300 57.500 1918.560 57.760 ;
        RECT 1918.300 2.420 1918.560 2.680 ;
        RECT 1923.360 2.420 1923.620 2.680 ;
      LAYER met2 ;
        RECT 1510.190 1100.580 1510.470 1104.000 ;
        RECT 1510.190 1100.000 1510.480 1100.580 ;
        RECT 1510.340 57.790 1510.480 1100.000 ;
        RECT 1510.280 57.470 1510.540 57.790 ;
        RECT 1918.300 57.470 1918.560 57.790 ;
        RECT 1918.360 2.710 1918.500 57.470 ;
        RECT 1918.300 2.390 1918.560 2.710 ;
        RECT 1923.360 2.390 1923.620 2.710 ;
        RECT 1923.420 2.000 1923.560 2.390 ;
        RECT 1923.210 -4.000 1923.770 2.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1517.150 58.040 1517.470 58.100 ;
        RECT 1938.970 58.040 1939.290 58.100 ;
        RECT 1517.150 57.900 1939.290 58.040 ;
        RECT 1517.150 57.840 1517.470 57.900 ;
        RECT 1938.970 57.840 1939.290 57.900 ;
      LAYER via ;
        RECT 1517.180 57.840 1517.440 58.100 ;
        RECT 1939.000 57.840 1939.260 58.100 ;
      LAYER met2 ;
        RECT 1516.170 1100.650 1516.450 1104.000 ;
        RECT 1516.170 1100.510 1517.380 1100.650 ;
        RECT 1516.170 1100.000 1516.450 1100.510 ;
        RECT 1517.240 58.130 1517.380 1100.510 ;
        RECT 1517.180 57.810 1517.440 58.130 ;
        RECT 1939.000 57.810 1939.260 58.130 ;
        RECT 1939.060 2.450 1939.200 57.810 ;
        RECT 1939.060 2.310 1941.500 2.450 ;
        RECT 1941.360 2.000 1941.500 2.310 ;
        RECT 1941.150 -4.000 1941.710 2.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1524.050 58.380 1524.370 58.440 ;
        RECT 1952.770 58.380 1953.090 58.440 ;
        RECT 1524.050 58.240 1953.090 58.380 ;
        RECT 1524.050 58.180 1524.370 58.240 ;
        RECT 1952.770 58.180 1953.090 58.240 ;
        RECT 1952.770 14.520 1953.090 14.580 ;
        RECT 1959.210 14.520 1959.530 14.580 ;
        RECT 1952.770 14.380 1959.530 14.520 ;
        RECT 1952.770 14.320 1953.090 14.380 ;
        RECT 1959.210 14.320 1959.530 14.380 ;
      LAYER via ;
        RECT 1524.080 58.180 1524.340 58.440 ;
        RECT 1952.800 58.180 1953.060 58.440 ;
        RECT 1952.800 14.320 1953.060 14.580 ;
        RECT 1959.240 14.320 1959.500 14.580 ;
      LAYER met2 ;
        RECT 1522.150 1100.650 1522.430 1104.000 ;
        RECT 1522.150 1100.510 1524.280 1100.650 ;
        RECT 1522.150 1100.000 1522.430 1100.510 ;
        RECT 1524.140 58.470 1524.280 1100.510 ;
        RECT 1524.080 58.150 1524.340 58.470 ;
        RECT 1952.800 58.150 1953.060 58.470 ;
        RECT 1952.860 14.610 1953.000 58.150 ;
        RECT 1952.800 14.290 1953.060 14.610 ;
        RECT 1959.240 14.290 1959.500 14.610 ;
        RECT 1959.300 2.000 1959.440 14.290 ;
        RECT 1959.090 -4.000 1959.650 2.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1531.410 41.720 1531.730 41.780 ;
        RECT 1977.150 41.720 1977.470 41.780 ;
        RECT 1531.410 41.580 1977.470 41.720 ;
        RECT 1531.410 41.520 1531.730 41.580 ;
        RECT 1977.150 41.520 1977.470 41.580 ;
      LAYER via ;
        RECT 1531.440 41.520 1531.700 41.780 ;
        RECT 1977.180 41.520 1977.440 41.780 ;
      LAYER met2 ;
        RECT 1528.130 1100.650 1528.410 1104.000 ;
        RECT 1528.130 1100.510 1530.260 1100.650 ;
        RECT 1528.130 1100.000 1528.410 1100.510 ;
        RECT 1530.120 1084.330 1530.260 1100.510 ;
        RECT 1530.120 1084.190 1531.640 1084.330 ;
        RECT 1531.500 41.810 1531.640 1084.190 ;
        RECT 1531.440 41.490 1531.700 41.810 ;
        RECT 1977.180 41.490 1977.440 41.810 ;
        RECT 1977.240 2.000 1977.380 41.490 ;
        RECT 1977.030 -4.000 1977.590 2.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1534.630 1083.480 1534.950 1083.540 ;
        RECT 1538.310 1083.480 1538.630 1083.540 ;
        RECT 1534.630 1083.340 1538.630 1083.480 ;
        RECT 1534.630 1083.280 1534.950 1083.340 ;
        RECT 1538.310 1083.280 1538.630 1083.340 ;
        RECT 1538.310 42.060 1538.630 42.120 ;
        RECT 1995.090 42.060 1995.410 42.120 ;
        RECT 1538.310 41.920 1995.410 42.060 ;
        RECT 1538.310 41.860 1538.630 41.920 ;
        RECT 1995.090 41.860 1995.410 41.920 ;
      LAYER via ;
        RECT 1534.660 1083.280 1534.920 1083.540 ;
        RECT 1538.340 1083.280 1538.600 1083.540 ;
        RECT 1538.340 41.860 1538.600 42.120 ;
        RECT 1995.120 41.860 1995.380 42.120 ;
      LAYER met2 ;
        RECT 1534.570 1100.580 1534.850 1104.000 ;
        RECT 1534.570 1100.000 1534.860 1100.580 ;
        RECT 1534.720 1083.570 1534.860 1100.000 ;
        RECT 1534.660 1083.250 1534.920 1083.570 ;
        RECT 1538.340 1083.250 1538.600 1083.570 ;
        RECT 1538.400 42.150 1538.540 1083.250 ;
        RECT 1538.340 41.830 1538.600 42.150 ;
        RECT 1995.120 41.830 1995.380 42.150 ;
        RECT 1995.180 2.000 1995.320 41.830 ;
        RECT 1994.970 -4.000 1995.530 2.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1540.610 1083.480 1540.930 1083.540 ;
        RECT 1544.750 1083.480 1545.070 1083.540 ;
        RECT 1540.610 1083.340 1545.070 1083.480 ;
        RECT 1540.610 1083.280 1540.930 1083.340 ;
        RECT 1544.750 1083.280 1545.070 1083.340 ;
        RECT 1544.750 42.400 1545.070 42.460 ;
        RECT 2012.570 42.400 2012.890 42.460 ;
        RECT 1544.750 42.260 2012.890 42.400 ;
        RECT 1544.750 42.200 1545.070 42.260 ;
        RECT 2012.570 42.200 2012.890 42.260 ;
      LAYER via ;
        RECT 1540.640 1083.280 1540.900 1083.540 ;
        RECT 1544.780 1083.280 1545.040 1083.540 ;
        RECT 1544.780 42.200 1545.040 42.460 ;
        RECT 2012.600 42.200 2012.860 42.460 ;
      LAYER met2 ;
        RECT 1540.550 1100.580 1540.830 1104.000 ;
        RECT 1540.550 1100.000 1540.840 1100.580 ;
        RECT 1540.700 1083.570 1540.840 1100.000 ;
        RECT 1540.640 1083.250 1540.900 1083.570 ;
        RECT 1544.780 1083.250 1545.040 1083.570 ;
        RECT 1544.840 42.490 1544.980 1083.250 ;
        RECT 1544.780 42.170 1545.040 42.490 ;
        RECT 2012.600 42.170 2012.860 42.490 ;
        RECT 2012.660 2.000 2012.800 42.170 ;
        RECT 2012.450 -4.000 2013.010 2.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1546.590 1083.480 1546.910 1083.540 ;
        RECT 1551.650 1083.480 1551.970 1083.540 ;
        RECT 1546.590 1083.340 1551.970 1083.480 ;
        RECT 1546.590 1083.280 1546.910 1083.340 ;
        RECT 1551.650 1083.280 1551.970 1083.340 ;
        RECT 1551.650 42.740 1551.970 42.800 ;
        RECT 2030.510 42.740 2030.830 42.800 ;
        RECT 1551.650 42.600 2030.830 42.740 ;
        RECT 1551.650 42.540 1551.970 42.600 ;
        RECT 2030.510 42.540 2030.830 42.600 ;
      LAYER via ;
        RECT 1546.620 1083.280 1546.880 1083.540 ;
        RECT 1551.680 1083.280 1551.940 1083.540 ;
        RECT 1551.680 42.540 1551.940 42.800 ;
        RECT 2030.540 42.540 2030.800 42.800 ;
      LAYER met2 ;
        RECT 1546.530 1100.580 1546.810 1104.000 ;
        RECT 1546.530 1100.000 1546.820 1100.580 ;
        RECT 1546.680 1083.570 1546.820 1100.000 ;
        RECT 1546.620 1083.250 1546.880 1083.570 ;
        RECT 1551.680 1083.250 1551.940 1083.570 ;
        RECT 1551.740 42.830 1551.880 1083.250 ;
        RECT 1551.680 42.510 1551.940 42.830 ;
        RECT 2030.540 42.510 2030.800 42.830 ;
        RECT 2030.600 2.000 2030.740 42.510 ;
        RECT 2030.390 -4.000 2030.950 2.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1553.030 1083.480 1553.350 1083.540 ;
        RECT 1558.090 1083.480 1558.410 1083.540 ;
        RECT 1553.030 1083.340 1558.410 1083.480 ;
        RECT 1553.030 1083.280 1553.350 1083.340 ;
        RECT 1558.090 1083.280 1558.410 1083.340 ;
        RECT 1558.090 43.080 1558.410 43.140 ;
        RECT 2048.450 43.080 2048.770 43.140 ;
        RECT 1558.090 42.940 2048.770 43.080 ;
        RECT 1558.090 42.880 1558.410 42.940 ;
        RECT 2048.450 42.880 2048.770 42.940 ;
      LAYER via ;
        RECT 1553.060 1083.280 1553.320 1083.540 ;
        RECT 1558.120 1083.280 1558.380 1083.540 ;
        RECT 1558.120 42.880 1558.380 43.140 ;
        RECT 2048.480 42.880 2048.740 43.140 ;
      LAYER met2 ;
        RECT 1552.970 1100.580 1553.250 1104.000 ;
        RECT 1552.970 1100.000 1553.260 1100.580 ;
        RECT 1553.120 1083.570 1553.260 1100.000 ;
        RECT 1553.060 1083.250 1553.320 1083.570 ;
        RECT 1558.120 1083.250 1558.380 1083.570 ;
        RECT 1558.180 43.170 1558.320 1083.250 ;
        RECT 1558.120 42.850 1558.380 43.170 ;
        RECT 2048.480 42.850 2048.740 43.170 ;
        RECT 2048.540 2.000 2048.680 42.850 ;
        RECT 2048.330 -4.000 2048.890 2.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 765.510 49.880 765.830 49.940 ;
        RECT 1111.890 49.880 1112.210 49.940 ;
        RECT 765.510 49.740 1112.210 49.880 ;
        RECT 765.510 49.680 765.830 49.740 ;
        RECT 1111.890 49.680 1112.210 49.740 ;
      LAYER via ;
        RECT 765.540 49.680 765.800 49.940 ;
        RECT 1111.920 49.680 1112.180 49.940 ;
      LAYER met2 ;
        RECT 1111.830 1100.580 1112.110 1104.000 ;
        RECT 1111.830 1100.000 1112.120 1100.580 ;
        RECT 1111.980 49.970 1112.120 1100.000 ;
        RECT 765.540 49.650 765.800 49.970 ;
        RECT 1111.920 49.650 1112.180 49.970 ;
        RECT 765.600 17.410 765.740 49.650 ;
        RECT 763.760 17.270 765.740 17.410 ;
        RECT 763.760 2.000 763.900 17.270 ;
        RECT 763.550 -4.000 764.110 2.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1558.550 43.420 1558.870 43.480 ;
        RECT 2066.390 43.420 2066.710 43.480 ;
        RECT 1558.550 43.280 2066.710 43.420 ;
        RECT 1558.550 43.220 1558.870 43.280 ;
        RECT 2066.390 43.220 2066.710 43.280 ;
      LAYER via ;
        RECT 1558.580 43.220 1558.840 43.480 ;
        RECT 2066.420 43.220 2066.680 43.480 ;
      LAYER met2 ;
        RECT 1558.950 1100.650 1559.230 1104.000 ;
        RECT 1558.640 1100.510 1559.230 1100.650 ;
        RECT 1558.640 43.510 1558.780 1100.510 ;
        RECT 1558.950 1100.000 1559.230 1100.510 ;
        RECT 1558.580 43.190 1558.840 43.510 ;
        RECT 2066.420 43.190 2066.680 43.510 ;
        RECT 2066.480 2.000 2066.620 43.190 ;
        RECT 2066.270 -4.000 2066.830 2.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1565.450 43.760 1565.770 43.820 ;
        RECT 2084.330 43.760 2084.650 43.820 ;
        RECT 1565.450 43.620 2084.650 43.760 ;
        RECT 1565.450 43.560 1565.770 43.620 ;
        RECT 2084.330 43.560 2084.650 43.620 ;
      LAYER via ;
        RECT 1565.480 43.560 1565.740 43.820 ;
        RECT 2084.360 43.560 2084.620 43.820 ;
      LAYER met2 ;
        RECT 1564.930 1100.650 1565.210 1104.000 ;
        RECT 1564.930 1100.510 1565.680 1100.650 ;
        RECT 1564.930 1100.000 1565.210 1100.510 ;
        RECT 1565.540 43.850 1565.680 1100.510 ;
        RECT 1565.480 43.530 1565.740 43.850 ;
        RECT 2084.360 43.530 2084.620 43.850 ;
        RECT 2084.420 2.000 2084.560 43.530 ;
        RECT 2084.210 -4.000 2084.770 2.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1572.350 44.100 1572.670 44.160 ;
        RECT 2101.810 44.100 2102.130 44.160 ;
        RECT 1572.350 43.960 2102.130 44.100 ;
        RECT 1572.350 43.900 1572.670 43.960 ;
        RECT 2101.810 43.900 2102.130 43.960 ;
      LAYER via ;
        RECT 1572.380 43.900 1572.640 44.160 ;
        RECT 2101.840 43.900 2102.100 44.160 ;
      LAYER met2 ;
        RECT 1571.370 1100.650 1571.650 1104.000 ;
        RECT 1571.370 1100.510 1572.580 1100.650 ;
        RECT 1571.370 1100.000 1571.650 1100.510 ;
        RECT 1572.440 44.190 1572.580 1100.510 ;
        RECT 1572.380 43.870 1572.640 44.190 ;
        RECT 2101.840 43.870 2102.100 44.190 ;
        RECT 2101.900 2.000 2102.040 43.870 ;
        RECT 2101.690 -4.000 2102.250 2.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1579.325 1014.305 1579.495 1028.415 ;
        RECT 1578.865 959.225 1579.035 980.475 ;
        RECT 1578.405 910.945 1578.575 958.715 ;
        RECT 1579.325 662.405 1579.495 710.515 ;
        RECT 1579.325 572.645 1579.495 593.895 ;
        RECT 1579.325 524.365 1579.495 545.615 ;
        RECT 1578.865 434.945 1579.035 484.755 ;
      LAYER mcon ;
        RECT 1579.325 1028.245 1579.495 1028.415 ;
        RECT 1578.865 980.305 1579.035 980.475 ;
        RECT 1578.405 958.545 1578.575 958.715 ;
        RECT 1579.325 710.345 1579.495 710.515 ;
        RECT 1579.325 593.725 1579.495 593.895 ;
        RECT 1579.325 545.445 1579.495 545.615 ;
        RECT 1578.865 484.585 1579.035 484.755 ;
      LAYER met1 ;
        RECT 1578.790 1097.080 1579.110 1097.140 ;
        RECT 1579.710 1097.080 1580.030 1097.140 ;
        RECT 1578.790 1096.940 1580.030 1097.080 ;
        RECT 1578.790 1096.880 1579.110 1096.940 ;
        RECT 1579.710 1096.880 1580.030 1096.940 ;
        RECT 1579.250 1028.400 1579.570 1028.460 ;
        RECT 1579.055 1028.260 1579.570 1028.400 ;
        RECT 1579.250 1028.200 1579.570 1028.260 ;
        RECT 1579.250 1014.460 1579.570 1014.520 ;
        RECT 1579.055 1014.320 1579.570 1014.460 ;
        RECT 1579.250 1014.260 1579.570 1014.320 ;
        RECT 1578.805 980.460 1579.095 980.505 ;
        RECT 1579.250 980.460 1579.570 980.520 ;
        RECT 1578.805 980.320 1579.570 980.460 ;
        RECT 1578.805 980.275 1579.095 980.320 ;
        RECT 1579.250 980.260 1579.570 980.320 ;
        RECT 1578.790 959.380 1579.110 959.440 ;
        RECT 1578.595 959.240 1579.110 959.380 ;
        RECT 1578.790 959.180 1579.110 959.240 ;
        RECT 1578.345 958.700 1578.635 958.745 ;
        RECT 1578.790 958.700 1579.110 958.760 ;
        RECT 1578.345 958.560 1579.110 958.700 ;
        RECT 1578.345 958.515 1578.635 958.560 ;
        RECT 1578.790 958.500 1579.110 958.560 ;
        RECT 1578.330 911.100 1578.650 911.160 ;
        RECT 1578.135 910.960 1578.650 911.100 ;
        RECT 1578.330 910.900 1578.650 910.960 ;
        RECT 1578.330 821.340 1578.650 821.400 ;
        RECT 1578.790 821.340 1579.110 821.400 ;
        RECT 1578.330 821.200 1579.110 821.340 ;
        RECT 1578.330 821.140 1578.650 821.200 ;
        RECT 1578.790 821.140 1579.110 821.200 ;
        RECT 1578.790 766.600 1579.110 766.660 ;
        RECT 1579.250 766.600 1579.570 766.660 ;
        RECT 1578.790 766.460 1579.570 766.600 ;
        RECT 1578.790 766.400 1579.110 766.460 ;
        RECT 1579.250 766.400 1579.570 766.460 ;
        RECT 1578.790 738.520 1579.110 738.780 ;
        RECT 1578.880 738.100 1579.020 738.520 ;
        RECT 1578.790 737.840 1579.110 738.100 ;
        RECT 1579.250 710.500 1579.570 710.560 ;
        RECT 1579.055 710.360 1579.570 710.500 ;
        RECT 1579.250 710.300 1579.570 710.360 ;
        RECT 1579.250 662.560 1579.570 662.620 ;
        RECT 1579.055 662.420 1579.570 662.560 ;
        RECT 1579.250 662.360 1579.570 662.420 ;
        RECT 1579.250 593.880 1579.570 593.940 ;
        RECT 1579.055 593.740 1579.570 593.880 ;
        RECT 1579.250 593.680 1579.570 593.740 ;
        RECT 1579.250 572.800 1579.570 572.860 ;
        RECT 1579.055 572.660 1579.570 572.800 ;
        RECT 1579.250 572.600 1579.570 572.660 ;
        RECT 1579.250 545.600 1579.570 545.660 ;
        RECT 1579.055 545.460 1579.570 545.600 ;
        RECT 1579.250 545.400 1579.570 545.460 ;
        RECT 1579.250 524.520 1579.570 524.580 ;
        RECT 1579.055 524.380 1579.570 524.520 ;
        RECT 1579.250 524.320 1579.570 524.380 ;
        RECT 1578.790 484.740 1579.110 484.800 ;
        RECT 1578.595 484.600 1579.110 484.740 ;
        RECT 1578.790 484.540 1579.110 484.600 ;
        RECT 1578.790 435.100 1579.110 435.160 ;
        RECT 1578.595 434.960 1579.110 435.100 ;
        RECT 1578.790 434.900 1579.110 434.960 ;
        RECT 1578.790 289.920 1579.110 289.980 ;
        RECT 1579.250 289.920 1579.570 289.980 ;
        RECT 1578.790 289.780 1579.570 289.920 ;
        RECT 1578.790 289.720 1579.110 289.780 ;
        RECT 1579.250 289.720 1579.570 289.780 ;
        RECT 1579.250 44.440 1579.570 44.500 ;
        RECT 2119.750 44.440 2120.070 44.500 ;
        RECT 1579.250 44.300 2120.070 44.440 ;
        RECT 1579.250 44.240 1579.570 44.300 ;
        RECT 2119.750 44.240 2120.070 44.300 ;
      LAYER via ;
        RECT 1578.820 1096.880 1579.080 1097.140 ;
        RECT 1579.740 1096.880 1580.000 1097.140 ;
        RECT 1579.280 1028.200 1579.540 1028.460 ;
        RECT 1579.280 1014.260 1579.540 1014.520 ;
        RECT 1579.280 980.260 1579.540 980.520 ;
        RECT 1578.820 959.180 1579.080 959.440 ;
        RECT 1578.820 958.500 1579.080 958.760 ;
        RECT 1578.360 910.900 1578.620 911.160 ;
        RECT 1578.360 821.140 1578.620 821.400 ;
        RECT 1578.820 821.140 1579.080 821.400 ;
        RECT 1578.820 766.400 1579.080 766.660 ;
        RECT 1579.280 766.400 1579.540 766.660 ;
        RECT 1578.820 738.520 1579.080 738.780 ;
        RECT 1578.820 737.840 1579.080 738.100 ;
        RECT 1579.280 710.300 1579.540 710.560 ;
        RECT 1579.280 662.360 1579.540 662.620 ;
        RECT 1579.280 593.680 1579.540 593.940 ;
        RECT 1579.280 572.600 1579.540 572.860 ;
        RECT 1579.280 545.400 1579.540 545.660 ;
        RECT 1579.280 524.320 1579.540 524.580 ;
        RECT 1578.820 484.540 1579.080 484.800 ;
        RECT 1578.820 434.900 1579.080 435.160 ;
        RECT 1578.820 289.720 1579.080 289.980 ;
        RECT 1579.280 289.720 1579.540 289.980 ;
        RECT 1579.280 44.240 1579.540 44.500 ;
        RECT 2119.780 44.240 2120.040 44.500 ;
      LAYER met2 ;
        RECT 1577.350 1100.650 1577.630 1104.000 ;
        RECT 1577.350 1100.510 1579.020 1100.650 ;
        RECT 1577.350 1100.000 1577.630 1100.510 ;
        RECT 1578.880 1097.170 1579.020 1100.510 ;
        RECT 1578.820 1096.850 1579.080 1097.170 ;
        RECT 1579.740 1096.850 1580.000 1097.170 ;
        RECT 1579.800 1089.090 1579.940 1096.850 ;
        RECT 1579.340 1088.950 1579.940 1089.090 ;
        RECT 1579.340 1028.490 1579.480 1088.950 ;
        RECT 1579.280 1028.170 1579.540 1028.490 ;
        RECT 1579.280 1014.230 1579.540 1014.550 ;
        RECT 1579.340 980.550 1579.480 1014.230 ;
        RECT 1579.280 980.230 1579.540 980.550 ;
        RECT 1578.820 959.150 1579.080 959.470 ;
        RECT 1578.880 958.790 1579.020 959.150 ;
        RECT 1578.820 958.470 1579.080 958.790 ;
        RECT 1578.360 910.870 1578.620 911.190 ;
        RECT 1578.420 870.130 1578.560 910.870 ;
        RECT 1577.960 869.990 1578.560 870.130 ;
        RECT 1577.960 868.770 1578.100 869.990 ;
        RECT 1577.960 868.630 1578.560 868.770 ;
        RECT 1578.420 821.430 1578.560 868.630 ;
        RECT 1578.360 821.110 1578.620 821.430 ;
        RECT 1578.820 821.110 1579.080 821.430 ;
        RECT 1578.880 787.850 1579.020 821.110 ;
        RECT 1578.880 787.710 1579.480 787.850 ;
        RECT 1579.340 766.690 1579.480 787.710 ;
        RECT 1578.820 766.370 1579.080 766.690 ;
        RECT 1579.280 766.370 1579.540 766.690 ;
        RECT 1578.880 738.810 1579.020 766.370 ;
        RECT 1578.820 738.490 1579.080 738.810 ;
        RECT 1578.820 737.810 1579.080 738.130 ;
        RECT 1578.880 717.810 1579.020 737.810 ;
        RECT 1578.880 717.670 1579.480 717.810 ;
        RECT 1579.340 710.590 1579.480 717.670 ;
        RECT 1579.280 710.270 1579.540 710.590 ;
        RECT 1579.280 662.330 1579.540 662.650 ;
        RECT 1579.340 593.970 1579.480 662.330 ;
        RECT 1579.280 593.650 1579.540 593.970 ;
        RECT 1579.280 572.570 1579.540 572.890 ;
        RECT 1579.340 545.690 1579.480 572.570 ;
        RECT 1579.280 545.370 1579.540 545.690 ;
        RECT 1579.280 524.290 1579.540 524.610 ;
        RECT 1579.340 524.010 1579.480 524.290 ;
        RECT 1578.880 523.870 1579.480 524.010 ;
        RECT 1578.880 484.830 1579.020 523.870 ;
        RECT 1578.820 484.510 1579.080 484.830 ;
        RECT 1578.820 434.870 1579.080 435.190 ;
        RECT 1578.880 290.010 1579.020 434.870 ;
        RECT 1578.820 289.690 1579.080 290.010 ;
        RECT 1579.280 289.690 1579.540 290.010 ;
        RECT 1579.340 110.570 1579.480 289.690 ;
        RECT 1578.880 110.430 1579.480 110.570 ;
        RECT 1578.880 109.890 1579.020 110.430 ;
        RECT 1578.880 109.750 1579.480 109.890 ;
        RECT 1579.340 44.530 1579.480 109.750 ;
        RECT 1579.280 44.210 1579.540 44.530 ;
        RECT 2119.780 44.210 2120.040 44.530 ;
        RECT 2119.840 2.000 2119.980 44.210 ;
        RECT 2119.630 -4.000 2120.190 2.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1585.765 786.505 1585.935 814.215 ;
        RECT 1586.225 717.825 1586.395 738.395 ;
        RECT 1586.225 483.225 1586.395 548.675 ;
        RECT 1585.765 186.405 1585.935 234.515 ;
        RECT 1585.765 96.645 1585.935 144.415 ;
      LAYER mcon ;
        RECT 1585.765 814.045 1585.935 814.215 ;
        RECT 1586.225 738.225 1586.395 738.395 ;
        RECT 1586.225 548.505 1586.395 548.675 ;
        RECT 1585.765 234.345 1585.935 234.515 ;
        RECT 1585.765 144.245 1585.935 144.415 ;
      LAYER met1 ;
        RECT 1585.230 835.280 1585.550 835.340 ;
        RECT 1585.230 835.140 1585.920 835.280 ;
        RECT 1585.230 835.080 1585.550 835.140 ;
        RECT 1585.780 835.000 1585.920 835.140 ;
        RECT 1585.690 834.740 1586.010 835.000 ;
        RECT 1585.690 814.200 1586.010 814.260 ;
        RECT 1585.495 814.060 1586.010 814.200 ;
        RECT 1585.690 814.000 1586.010 814.060 ;
        RECT 1585.690 786.660 1586.010 786.720 ;
        RECT 1585.495 786.520 1586.010 786.660 ;
        RECT 1585.690 786.460 1586.010 786.520 ;
        RECT 1586.150 738.380 1586.470 738.440 ;
        RECT 1585.955 738.240 1586.470 738.380 ;
        RECT 1586.150 738.180 1586.470 738.240 ;
        RECT 1586.150 717.980 1586.470 718.040 ;
        RECT 1585.955 717.840 1586.470 717.980 ;
        RECT 1586.150 717.780 1586.470 717.840 ;
        RECT 1585.690 676.160 1586.010 676.220 ;
        RECT 1586.150 676.160 1586.470 676.220 ;
        RECT 1585.690 676.020 1586.470 676.160 ;
        RECT 1585.690 675.960 1586.010 676.020 ;
        RECT 1586.150 675.960 1586.470 676.020 ;
        RECT 1586.150 548.660 1586.470 548.720 ;
        RECT 1585.955 548.520 1586.470 548.660 ;
        RECT 1586.150 548.460 1586.470 548.520 ;
        RECT 1586.150 483.380 1586.470 483.440 ;
        RECT 1585.955 483.240 1586.470 483.380 ;
        RECT 1586.150 483.180 1586.470 483.240 ;
        RECT 1585.230 338.200 1585.550 338.260 ;
        RECT 1586.150 338.200 1586.470 338.260 ;
        RECT 1585.230 338.060 1586.470 338.200 ;
        RECT 1585.230 338.000 1585.550 338.060 ;
        RECT 1586.150 338.000 1586.470 338.060 ;
        RECT 1585.690 234.500 1586.010 234.560 ;
        RECT 1585.495 234.360 1586.010 234.500 ;
        RECT 1585.690 234.300 1586.010 234.360 ;
        RECT 1585.705 186.560 1585.995 186.605 ;
        RECT 1586.150 186.560 1586.470 186.620 ;
        RECT 1585.705 186.420 1586.470 186.560 ;
        RECT 1585.705 186.375 1585.995 186.420 ;
        RECT 1586.150 186.360 1586.470 186.420 ;
        RECT 1585.690 145.080 1586.010 145.140 ;
        RECT 1586.150 145.080 1586.470 145.140 ;
        RECT 1585.690 144.940 1586.470 145.080 ;
        RECT 1585.690 144.880 1586.010 144.940 ;
        RECT 1586.150 144.880 1586.470 144.940 ;
        RECT 1585.690 144.400 1586.010 144.460 ;
        RECT 1585.495 144.260 1586.010 144.400 ;
        RECT 1585.690 144.200 1586.010 144.260 ;
        RECT 1585.705 96.800 1585.995 96.845 ;
        RECT 1586.150 96.800 1586.470 96.860 ;
        RECT 1585.705 96.660 1586.470 96.800 ;
        RECT 1585.705 96.615 1585.995 96.660 ;
        RECT 1586.150 96.600 1586.470 96.660 ;
        RECT 1585.230 48.180 1585.550 48.240 ;
        RECT 2137.690 48.180 2138.010 48.240 ;
        RECT 1585.230 48.040 2138.010 48.180 ;
        RECT 1585.230 47.980 1585.550 48.040 ;
        RECT 2137.690 47.980 2138.010 48.040 ;
      LAYER via ;
        RECT 1585.260 835.080 1585.520 835.340 ;
        RECT 1585.720 834.740 1585.980 835.000 ;
        RECT 1585.720 814.000 1585.980 814.260 ;
        RECT 1585.720 786.460 1585.980 786.720 ;
        RECT 1586.180 738.180 1586.440 738.440 ;
        RECT 1586.180 717.780 1586.440 718.040 ;
        RECT 1585.720 675.960 1585.980 676.220 ;
        RECT 1586.180 675.960 1586.440 676.220 ;
        RECT 1586.180 548.460 1586.440 548.720 ;
        RECT 1586.180 483.180 1586.440 483.440 ;
        RECT 1585.260 338.000 1585.520 338.260 ;
        RECT 1586.180 338.000 1586.440 338.260 ;
        RECT 1585.720 234.300 1585.980 234.560 ;
        RECT 1586.180 186.360 1586.440 186.620 ;
        RECT 1585.720 144.880 1585.980 145.140 ;
        RECT 1586.180 144.880 1586.440 145.140 ;
        RECT 1585.720 144.200 1585.980 144.460 ;
        RECT 1586.180 96.600 1586.440 96.860 ;
        RECT 1585.260 47.980 1585.520 48.240 ;
        RECT 2137.720 47.980 2137.980 48.240 ;
      LAYER met2 ;
        RECT 1583.330 1100.650 1583.610 1104.000 ;
        RECT 1583.330 1100.510 1585.460 1100.650 ;
        RECT 1583.330 1100.000 1583.610 1100.510 ;
        RECT 1585.320 1085.010 1585.460 1100.510 ;
        RECT 1585.320 1084.870 1586.380 1085.010 ;
        RECT 1586.240 1028.570 1586.380 1084.870 ;
        RECT 1585.320 1028.430 1586.380 1028.570 ;
        RECT 1585.320 1027.890 1585.460 1028.430 ;
        RECT 1585.320 1027.750 1585.920 1027.890 ;
        RECT 1585.780 932.010 1585.920 1027.750 ;
        RECT 1585.320 931.870 1585.920 932.010 ;
        RECT 1585.320 931.330 1585.460 931.870 ;
        RECT 1585.320 931.190 1586.380 931.330 ;
        RECT 1586.240 869.565 1586.380 931.190 ;
        RECT 1585.250 869.195 1585.530 869.565 ;
        RECT 1586.170 869.195 1586.450 869.565 ;
        RECT 1585.320 835.370 1585.460 869.195 ;
        RECT 1585.260 835.050 1585.520 835.370 ;
        RECT 1585.720 834.710 1585.980 835.030 ;
        RECT 1585.780 814.290 1585.920 834.710 ;
        RECT 1585.720 813.970 1585.980 814.290 ;
        RECT 1585.720 786.430 1585.980 786.750 ;
        RECT 1585.780 766.090 1585.920 786.430 ;
        RECT 1585.780 765.950 1586.380 766.090 ;
        RECT 1586.240 738.470 1586.380 765.950 ;
        RECT 1586.180 738.150 1586.440 738.470 ;
        RECT 1586.180 717.750 1586.440 718.070 ;
        RECT 1586.240 676.250 1586.380 717.750 ;
        RECT 1585.720 675.930 1585.980 676.250 ;
        RECT 1586.180 675.930 1586.440 676.250 ;
        RECT 1585.780 641.820 1585.920 675.930 ;
        RECT 1585.780 641.680 1586.380 641.820 ;
        RECT 1586.240 548.750 1586.380 641.680 ;
        RECT 1586.180 548.430 1586.440 548.750 ;
        RECT 1586.180 483.150 1586.440 483.470 ;
        RECT 1586.240 338.290 1586.380 483.150 ;
        RECT 1585.260 337.970 1585.520 338.290 ;
        RECT 1586.180 337.970 1586.440 338.290 ;
        RECT 1585.320 337.805 1585.460 337.970 ;
        RECT 1584.330 337.435 1584.610 337.805 ;
        RECT 1585.250 337.435 1585.530 337.805 ;
        RECT 1584.400 290.205 1584.540 337.435 ;
        RECT 1584.330 289.835 1584.610 290.205 ;
        RECT 1585.250 289.155 1585.530 289.525 ;
        RECT 1585.320 254.730 1585.460 289.155 ;
        RECT 1585.320 254.590 1585.920 254.730 ;
        RECT 1585.780 234.590 1585.920 254.590 ;
        RECT 1585.720 234.270 1585.980 234.590 ;
        RECT 1586.180 186.330 1586.440 186.650 ;
        RECT 1586.240 145.170 1586.380 186.330 ;
        RECT 1585.720 144.850 1585.980 145.170 ;
        RECT 1586.180 144.850 1586.440 145.170 ;
        RECT 1585.780 144.490 1585.920 144.850 ;
        RECT 1585.720 144.170 1585.980 144.490 ;
        RECT 1586.180 96.570 1586.440 96.890 ;
        RECT 1586.240 62.970 1586.380 96.570 ;
        RECT 1585.780 62.830 1586.380 62.970 ;
        RECT 1585.780 62.290 1585.920 62.830 ;
        RECT 1585.320 62.150 1585.920 62.290 ;
        RECT 1585.320 48.270 1585.460 62.150 ;
        RECT 1585.260 47.950 1585.520 48.270 ;
        RECT 2137.720 47.950 2137.980 48.270 ;
        RECT 2137.780 2.000 2137.920 47.950 ;
        RECT 2137.570 -4.000 2138.130 2.000 ;
      LAYER via2 ;
        RECT 1585.250 869.240 1585.530 869.520 ;
        RECT 1586.170 869.240 1586.450 869.520 ;
        RECT 1584.330 337.480 1584.610 337.760 ;
        RECT 1585.250 337.480 1585.530 337.760 ;
        RECT 1584.330 289.880 1584.610 290.160 ;
        RECT 1585.250 289.200 1585.530 289.480 ;
      LAYER met3 ;
        RECT 1585.225 869.530 1585.555 869.545 ;
        RECT 1586.145 869.530 1586.475 869.545 ;
        RECT 1585.225 869.230 1586.475 869.530 ;
        RECT 1585.225 869.215 1585.555 869.230 ;
        RECT 1586.145 869.215 1586.475 869.230 ;
        RECT 1584.305 337.770 1584.635 337.785 ;
        RECT 1585.225 337.770 1585.555 337.785 ;
        RECT 1584.305 337.470 1585.555 337.770 ;
        RECT 1584.305 337.455 1584.635 337.470 ;
        RECT 1585.225 337.455 1585.555 337.470 ;
        RECT 1584.305 290.170 1584.635 290.185 ;
        RECT 1584.305 289.870 1586.690 290.170 ;
        RECT 1584.305 289.855 1584.635 289.870 ;
        RECT 1585.225 289.490 1585.555 289.505 ;
        RECT 1586.390 289.490 1586.690 289.870 ;
        RECT 1585.225 289.190 1586.690 289.490 ;
        RECT 1585.225 289.175 1585.555 289.190 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1592.205 821.185 1592.375 845.835 ;
        RECT 1592.205 786.505 1592.375 814.215 ;
        RECT 1592.205 669.885 1592.375 717.655 ;
        RECT 1592.205 627.725 1592.375 669.375 ;
        RECT 1592.665 572.645 1592.835 620.755 ;
        RECT 1591.745 524.365 1591.915 546.975 ;
        RECT 1591.285 379.525 1591.455 387.855 ;
        RECT 1591.745 234.685 1591.915 282.795 ;
      LAYER mcon ;
        RECT 1592.205 845.665 1592.375 845.835 ;
        RECT 1592.205 814.045 1592.375 814.215 ;
        RECT 1592.205 717.485 1592.375 717.655 ;
        RECT 1592.205 669.205 1592.375 669.375 ;
        RECT 1592.665 620.585 1592.835 620.755 ;
        RECT 1591.745 546.805 1591.915 546.975 ;
        RECT 1591.285 387.685 1591.455 387.855 ;
        RECT 1591.745 282.625 1591.915 282.795 ;
      LAYER met1 ;
        RECT 1590.750 1085.180 1591.070 1085.240 ;
        RECT 1592.590 1085.180 1592.910 1085.240 ;
        RECT 1590.750 1085.040 1592.910 1085.180 ;
        RECT 1590.750 1084.980 1591.070 1085.040 ;
        RECT 1592.590 1084.980 1592.910 1085.040 ;
        RECT 1592.145 845.820 1592.435 845.865 ;
        RECT 1592.590 845.820 1592.910 845.880 ;
        RECT 1592.145 845.680 1592.910 845.820 ;
        RECT 1592.145 845.635 1592.435 845.680 ;
        RECT 1592.590 845.620 1592.910 845.680 ;
        RECT 1592.130 821.340 1592.450 821.400 ;
        RECT 1591.935 821.200 1592.450 821.340 ;
        RECT 1592.130 821.140 1592.450 821.200 ;
        RECT 1592.130 814.200 1592.450 814.260 ;
        RECT 1591.935 814.060 1592.450 814.200 ;
        RECT 1592.130 814.000 1592.450 814.060 ;
        RECT 1592.130 786.660 1592.450 786.720 ;
        RECT 1591.935 786.520 1592.450 786.660 ;
        RECT 1592.130 786.460 1592.450 786.520 ;
        RECT 1592.145 717.640 1592.435 717.685 ;
        RECT 1592.590 717.640 1592.910 717.700 ;
        RECT 1592.145 717.500 1592.910 717.640 ;
        RECT 1592.145 717.455 1592.435 717.500 ;
        RECT 1592.590 717.440 1592.910 717.500 ;
        RECT 1592.130 670.040 1592.450 670.100 ;
        RECT 1591.935 669.900 1592.450 670.040 ;
        RECT 1592.130 669.840 1592.450 669.900 ;
        RECT 1592.130 669.360 1592.450 669.420 ;
        RECT 1591.935 669.220 1592.450 669.360 ;
        RECT 1592.130 669.160 1592.450 669.220 ;
        RECT 1592.130 627.880 1592.450 627.940 ;
        RECT 1591.935 627.740 1592.450 627.880 ;
        RECT 1592.130 627.680 1592.450 627.740 ;
        RECT 1592.590 620.740 1592.910 620.800 ;
        RECT 1592.395 620.600 1592.910 620.740 ;
        RECT 1592.590 620.540 1592.910 620.600 ;
        RECT 1592.590 572.800 1592.910 572.860 ;
        RECT 1592.395 572.660 1592.910 572.800 ;
        RECT 1592.590 572.600 1592.910 572.660 ;
        RECT 1591.685 546.960 1591.975 547.005 ;
        RECT 1592.590 546.960 1592.910 547.020 ;
        RECT 1591.685 546.820 1592.910 546.960 ;
        RECT 1591.685 546.775 1591.975 546.820 ;
        RECT 1592.590 546.760 1592.910 546.820 ;
        RECT 1591.670 524.520 1591.990 524.580 ;
        RECT 1591.475 524.380 1591.990 524.520 ;
        RECT 1591.670 524.320 1591.990 524.380 ;
        RECT 1591.225 387.840 1591.515 387.885 ;
        RECT 1592.590 387.840 1592.910 387.900 ;
        RECT 1591.225 387.700 1592.910 387.840 ;
        RECT 1591.225 387.655 1591.515 387.700 ;
        RECT 1592.590 387.640 1592.910 387.700 ;
        RECT 1591.210 379.680 1591.530 379.740 ;
        RECT 1591.015 379.540 1591.530 379.680 ;
        RECT 1591.210 379.480 1591.530 379.540 ;
        RECT 1591.670 289.580 1591.990 289.640 ;
        RECT 1592.590 289.580 1592.910 289.640 ;
        RECT 1591.670 289.440 1592.910 289.580 ;
        RECT 1591.670 289.380 1591.990 289.440 ;
        RECT 1592.590 289.380 1592.910 289.440 ;
        RECT 1591.670 282.780 1591.990 282.840 ;
        RECT 1591.475 282.640 1591.990 282.780 ;
        RECT 1591.670 282.580 1591.990 282.640 ;
        RECT 1591.685 234.840 1591.975 234.885 ;
        RECT 1592.130 234.840 1592.450 234.900 ;
        RECT 1591.685 234.700 1592.450 234.840 ;
        RECT 1591.685 234.655 1591.975 234.700 ;
        RECT 1592.130 234.640 1592.450 234.700 ;
        RECT 1592.130 169.020 1592.450 169.280 ;
        RECT 1592.220 168.880 1592.360 169.020 ;
        RECT 1592.590 168.880 1592.910 168.940 ;
        RECT 1592.220 168.740 1592.910 168.880 ;
        RECT 1592.590 168.680 1592.910 168.740 ;
        RECT 1591.670 47.840 1591.990 47.900 ;
        RECT 2155.630 47.840 2155.950 47.900 ;
        RECT 1591.670 47.700 2155.950 47.840 ;
        RECT 1591.670 47.640 1591.990 47.700 ;
        RECT 2155.630 47.640 2155.950 47.700 ;
      LAYER via ;
        RECT 1590.780 1084.980 1591.040 1085.240 ;
        RECT 1592.620 1084.980 1592.880 1085.240 ;
        RECT 1592.620 845.620 1592.880 845.880 ;
        RECT 1592.160 821.140 1592.420 821.400 ;
        RECT 1592.160 814.000 1592.420 814.260 ;
        RECT 1592.160 786.460 1592.420 786.720 ;
        RECT 1592.620 717.440 1592.880 717.700 ;
        RECT 1592.160 669.840 1592.420 670.100 ;
        RECT 1592.160 669.160 1592.420 669.420 ;
        RECT 1592.160 627.680 1592.420 627.940 ;
        RECT 1592.620 620.540 1592.880 620.800 ;
        RECT 1592.620 572.600 1592.880 572.860 ;
        RECT 1592.620 546.760 1592.880 547.020 ;
        RECT 1591.700 524.320 1591.960 524.580 ;
        RECT 1592.620 387.640 1592.880 387.900 ;
        RECT 1591.240 379.480 1591.500 379.740 ;
        RECT 1591.700 289.380 1591.960 289.640 ;
        RECT 1592.620 289.380 1592.880 289.640 ;
        RECT 1591.700 282.580 1591.960 282.840 ;
        RECT 1592.160 234.640 1592.420 234.900 ;
        RECT 1592.160 169.020 1592.420 169.280 ;
        RECT 1592.620 168.680 1592.880 168.940 ;
        RECT 1591.700 47.640 1591.960 47.900 ;
        RECT 2155.660 47.640 2155.920 47.900 ;
      LAYER met2 ;
        RECT 1589.770 1100.650 1590.050 1104.000 ;
        RECT 1589.770 1100.510 1590.980 1100.650 ;
        RECT 1589.770 1100.000 1590.050 1100.510 ;
        RECT 1590.840 1085.270 1590.980 1100.510 ;
        RECT 1590.780 1084.950 1591.040 1085.270 ;
        RECT 1592.620 1084.950 1592.880 1085.270 ;
        RECT 1592.680 1028.570 1592.820 1084.950 ;
        RECT 1591.760 1028.430 1592.820 1028.570 ;
        RECT 1591.760 1027.890 1591.900 1028.430 ;
        RECT 1591.760 1027.750 1592.360 1027.890 ;
        RECT 1592.220 932.010 1592.360 1027.750 ;
        RECT 1591.760 931.870 1592.360 932.010 ;
        RECT 1591.760 931.330 1591.900 931.870 ;
        RECT 1591.760 931.190 1592.820 931.330 ;
        RECT 1592.680 845.910 1592.820 931.190 ;
        RECT 1592.620 845.590 1592.880 845.910 ;
        RECT 1592.160 821.110 1592.420 821.430 ;
        RECT 1592.220 814.290 1592.360 821.110 ;
        RECT 1592.160 813.970 1592.420 814.290 ;
        RECT 1592.160 786.430 1592.420 786.750 ;
        RECT 1592.220 766.090 1592.360 786.430 ;
        RECT 1592.220 765.950 1592.820 766.090 ;
        RECT 1592.680 739.005 1592.820 765.950 ;
        RECT 1592.610 738.635 1592.890 739.005 ;
        RECT 1592.610 717.555 1592.890 717.925 ;
        RECT 1592.620 717.410 1592.880 717.555 ;
        RECT 1592.160 669.810 1592.420 670.130 ;
        RECT 1592.220 669.450 1592.360 669.810 ;
        RECT 1592.160 669.130 1592.420 669.450 ;
        RECT 1592.160 627.650 1592.420 627.970 ;
        RECT 1592.220 621.250 1592.360 627.650 ;
        RECT 1592.220 621.110 1592.820 621.250 ;
        RECT 1592.680 620.830 1592.820 621.110 ;
        RECT 1592.620 620.510 1592.880 620.830 ;
        RECT 1592.620 572.570 1592.880 572.890 ;
        RECT 1592.680 547.050 1592.820 572.570 ;
        RECT 1592.620 546.730 1592.880 547.050 ;
        RECT 1591.700 524.290 1591.960 524.610 ;
        RECT 1591.760 483.325 1591.900 524.290 ;
        RECT 1591.690 482.955 1591.970 483.325 ;
        RECT 1592.610 482.955 1592.890 483.325 ;
        RECT 1592.680 387.930 1592.820 482.955 ;
        RECT 1592.620 387.610 1592.880 387.930 ;
        RECT 1591.240 379.450 1591.500 379.770 ;
        RECT 1591.300 351.290 1591.440 379.450 ;
        RECT 1591.300 351.150 1591.900 351.290 ;
        RECT 1591.760 337.805 1591.900 351.150 ;
        RECT 1591.690 337.435 1591.970 337.805 ;
        RECT 1592.610 336.755 1592.890 337.125 ;
        RECT 1592.680 289.670 1592.820 336.755 ;
        RECT 1591.700 289.350 1591.960 289.670 ;
        RECT 1592.620 289.350 1592.880 289.670 ;
        RECT 1591.760 282.870 1591.900 289.350 ;
        RECT 1591.700 282.550 1591.960 282.870 ;
        RECT 1592.160 234.610 1592.420 234.930 ;
        RECT 1592.220 234.445 1592.360 234.610 ;
        RECT 1592.150 234.075 1592.430 234.445 ;
        RECT 1591.690 233.395 1591.970 233.765 ;
        RECT 1591.760 206.450 1591.900 233.395 ;
        RECT 1591.760 206.310 1592.360 206.450 ;
        RECT 1592.220 169.310 1592.360 206.310 ;
        RECT 1592.160 168.990 1592.420 169.310 ;
        RECT 1592.620 168.650 1592.880 168.970 ;
        RECT 1592.680 62.970 1592.820 168.650 ;
        RECT 1592.220 62.830 1592.820 62.970 ;
        RECT 1592.220 62.290 1592.360 62.830 ;
        RECT 1591.760 62.150 1592.360 62.290 ;
        RECT 1591.760 47.930 1591.900 62.150 ;
        RECT 1591.700 47.610 1591.960 47.930 ;
        RECT 2155.660 47.610 2155.920 47.930 ;
        RECT 2155.720 2.000 2155.860 47.610 ;
        RECT 2155.510 -4.000 2156.070 2.000 ;
      LAYER via2 ;
        RECT 1592.610 738.680 1592.890 738.960 ;
        RECT 1592.610 717.600 1592.890 717.880 ;
        RECT 1591.690 483.000 1591.970 483.280 ;
        RECT 1592.610 483.000 1592.890 483.280 ;
        RECT 1591.690 337.480 1591.970 337.760 ;
        RECT 1592.610 336.800 1592.890 337.080 ;
        RECT 1592.150 234.120 1592.430 234.400 ;
        RECT 1591.690 233.440 1591.970 233.720 ;
      LAYER met3 ;
        RECT 1592.585 738.980 1592.915 738.985 ;
        RECT 1592.585 738.970 1593.170 738.980 ;
        RECT 1592.585 738.670 1593.370 738.970 ;
        RECT 1592.585 738.660 1593.170 738.670 ;
        RECT 1592.585 738.655 1592.915 738.660 ;
        RECT 1592.585 717.900 1592.915 717.905 ;
        RECT 1592.585 717.890 1593.170 717.900 ;
        RECT 1592.585 717.590 1593.370 717.890 ;
        RECT 1592.585 717.580 1593.170 717.590 ;
        RECT 1592.585 717.575 1592.915 717.580 ;
        RECT 1591.665 483.290 1591.995 483.305 ;
        RECT 1592.585 483.290 1592.915 483.305 ;
        RECT 1591.665 482.990 1592.915 483.290 ;
        RECT 1591.665 482.975 1591.995 482.990 ;
        RECT 1592.585 482.975 1592.915 482.990 ;
        RECT 1591.665 337.770 1591.995 337.785 ;
        RECT 1590.990 337.470 1591.995 337.770 ;
        RECT 1590.990 337.090 1591.290 337.470 ;
        RECT 1591.665 337.455 1591.995 337.470 ;
        RECT 1592.585 337.090 1592.915 337.105 ;
        RECT 1590.990 336.790 1592.915 337.090 ;
        RECT 1592.585 336.775 1592.915 336.790 ;
        RECT 1592.125 234.410 1592.455 234.425 ;
        RECT 1592.125 234.110 1593.130 234.410 ;
        RECT 1592.125 234.095 1592.455 234.110 ;
        RECT 1591.665 233.730 1591.995 233.745 ;
        RECT 1592.830 233.730 1593.130 234.110 ;
        RECT 1591.665 233.430 1593.130 233.730 ;
        RECT 1591.665 233.415 1591.995 233.430 ;
      LAYER via3 ;
        RECT 1592.820 738.660 1593.140 738.980 ;
        RECT 1592.820 717.580 1593.140 717.900 ;
      LAYER met4 ;
        RECT 1592.815 738.655 1593.145 738.985 ;
        RECT 1592.830 717.905 1593.130 738.655 ;
        RECT 1592.815 717.575 1593.145 717.905 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1595.810 1083.480 1596.130 1083.540 ;
        RECT 1599.950 1083.480 1600.270 1083.540 ;
        RECT 1595.810 1083.340 1600.270 1083.480 ;
        RECT 1595.810 1083.280 1596.130 1083.340 ;
        RECT 1599.950 1083.280 1600.270 1083.340 ;
        RECT 1599.950 47.500 1600.270 47.560 ;
        RECT 2173.110 47.500 2173.430 47.560 ;
        RECT 1599.950 47.360 2173.430 47.500 ;
        RECT 1599.950 47.300 1600.270 47.360 ;
        RECT 2173.110 47.300 2173.430 47.360 ;
      LAYER via ;
        RECT 1595.840 1083.280 1596.100 1083.540 ;
        RECT 1599.980 1083.280 1600.240 1083.540 ;
        RECT 1599.980 47.300 1600.240 47.560 ;
        RECT 2173.140 47.300 2173.400 47.560 ;
      LAYER met2 ;
        RECT 1595.750 1100.580 1596.030 1104.000 ;
        RECT 1595.750 1100.000 1596.040 1100.580 ;
        RECT 1595.900 1083.570 1596.040 1100.000 ;
        RECT 1595.840 1083.250 1596.100 1083.570 ;
        RECT 1599.980 1083.250 1600.240 1083.570 ;
        RECT 1600.040 47.590 1600.180 1083.250 ;
        RECT 1599.980 47.270 1600.240 47.590 ;
        RECT 2173.140 47.270 2173.400 47.590 ;
        RECT 2173.200 2.000 2173.340 47.270 ;
        RECT 2172.990 -4.000 2173.550 2.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1601.790 1083.480 1602.110 1083.540 ;
        RECT 1606.850 1083.480 1607.170 1083.540 ;
        RECT 1601.790 1083.340 1607.170 1083.480 ;
        RECT 1601.790 1083.280 1602.110 1083.340 ;
        RECT 1606.850 1083.280 1607.170 1083.340 ;
        RECT 1606.850 47.160 1607.170 47.220 ;
        RECT 2191.050 47.160 2191.370 47.220 ;
        RECT 1606.850 47.020 2191.370 47.160 ;
        RECT 1606.850 46.960 1607.170 47.020 ;
        RECT 2191.050 46.960 2191.370 47.020 ;
      LAYER via ;
        RECT 1601.820 1083.280 1602.080 1083.540 ;
        RECT 1606.880 1083.280 1607.140 1083.540 ;
        RECT 1606.880 46.960 1607.140 47.220 ;
        RECT 2191.080 46.960 2191.340 47.220 ;
      LAYER met2 ;
        RECT 1601.730 1100.580 1602.010 1104.000 ;
        RECT 1601.730 1100.000 1602.020 1100.580 ;
        RECT 1601.880 1083.570 1602.020 1100.000 ;
        RECT 1601.820 1083.250 1602.080 1083.570 ;
        RECT 1606.880 1083.250 1607.140 1083.570 ;
        RECT 1606.940 47.250 1607.080 1083.250 ;
        RECT 1606.880 46.930 1607.140 47.250 ;
        RECT 2191.080 46.930 2191.340 47.250 ;
        RECT 2191.140 2.000 2191.280 46.930 ;
        RECT 2190.930 -4.000 2191.490 2.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1608.230 1089.600 1608.550 1089.660 ;
        RECT 1613.290 1089.600 1613.610 1089.660 ;
        RECT 1608.230 1089.460 1613.610 1089.600 ;
        RECT 1608.230 1089.400 1608.550 1089.460 ;
        RECT 1613.290 1089.400 1613.610 1089.460 ;
        RECT 1613.290 46.820 1613.610 46.880 ;
        RECT 2208.990 46.820 2209.310 46.880 ;
        RECT 1613.290 46.680 2209.310 46.820 ;
        RECT 1613.290 46.620 1613.610 46.680 ;
        RECT 2208.990 46.620 2209.310 46.680 ;
      LAYER via ;
        RECT 1608.260 1089.400 1608.520 1089.660 ;
        RECT 1613.320 1089.400 1613.580 1089.660 ;
        RECT 1613.320 46.620 1613.580 46.880 ;
        RECT 2209.020 46.620 2209.280 46.880 ;
      LAYER met2 ;
        RECT 1608.170 1100.580 1608.450 1104.000 ;
        RECT 1608.170 1100.000 1608.460 1100.580 ;
        RECT 1608.320 1089.690 1608.460 1100.000 ;
        RECT 1608.260 1089.370 1608.520 1089.690 ;
        RECT 1613.320 1089.370 1613.580 1089.690 ;
        RECT 1613.380 46.910 1613.520 1089.370 ;
        RECT 1613.320 46.590 1613.580 46.910 ;
        RECT 2209.020 46.590 2209.280 46.910 ;
        RECT 2209.080 2.000 2209.220 46.590 ;
        RECT 2208.870 -4.000 2209.430 2.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1613.750 46.480 1614.070 46.540 ;
        RECT 2226.930 46.480 2227.250 46.540 ;
        RECT 1613.750 46.340 2227.250 46.480 ;
        RECT 1613.750 46.280 1614.070 46.340 ;
        RECT 2226.930 46.280 2227.250 46.340 ;
      LAYER via ;
        RECT 1613.780 46.280 1614.040 46.540 ;
        RECT 2226.960 46.280 2227.220 46.540 ;
      LAYER met2 ;
        RECT 1614.150 1100.650 1614.430 1104.000 ;
        RECT 1613.840 1100.510 1614.430 1100.650 ;
        RECT 1613.840 46.570 1613.980 1100.510 ;
        RECT 1614.150 1100.000 1614.430 1100.510 ;
        RECT 1613.780 46.250 1614.040 46.570 ;
        RECT 2226.960 46.250 2227.220 46.570 ;
        RECT 2227.020 2.000 2227.160 46.250 ;
        RECT 2226.810 -4.000 2227.370 2.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 786.210 49.540 786.530 49.600 ;
        RECT 1119.250 49.540 1119.570 49.600 ;
        RECT 786.210 49.400 1119.570 49.540 ;
        RECT 786.210 49.340 786.530 49.400 ;
        RECT 1119.250 49.340 1119.570 49.400 ;
      LAYER via ;
        RECT 786.240 49.340 786.500 49.600 ;
        RECT 1119.280 49.340 1119.540 49.600 ;
      LAYER met2 ;
        RECT 1118.270 1101.330 1118.550 1104.000 ;
        RECT 1118.270 1101.190 1119.480 1101.330 ;
        RECT 1118.270 1100.000 1118.550 1101.190 ;
        RECT 1119.340 49.630 1119.480 1101.190 ;
        RECT 786.240 49.310 786.500 49.630 ;
        RECT 1119.280 49.310 1119.540 49.630 ;
        RECT 786.300 17.410 786.440 49.310 ;
        RECT 781.700 17.270 786.440 17.410 ;
        RECT 781.700 2.000 781.840 17.270 ;
        RECT 781.490 -4.000 782.050 2.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1620.650 46.140 1620.970 46.200 ;
        RECT 2244.870 46.140 2245.190 46.200 ;
        RECT 1620.650 46.000 2245.190 46.140 ;
        RECT 1620.650 45.940 1620.970 46.000 ;
        RECT 2244.870 45.940 2245.190 46.000 ;
      LAYER via ;
        RECT 1620.680 45.940 1620.940 46.200 ;
        RECT 2244.900 45.940 2245.160 46.200 ;
      LAYER met2 ;
        RECT 1620.130 1100.650 1620.410 1104.000 ;
        RECT 1620.130 1100.510 1620.880 1100.650 ;
        RECT 1620.130 1100.000 1620.410 1100.510 ;
        RECT 1620.740 46.230 1620.880 1100.510 ;
        RECT 1620.680 45.910 1620.940 46.230 ;
        RECT 2244.900 45.910 2245.160 46.230 ;
        RECT 2244.960 2.000 2245.100 45.910 ;
        RECT 2244.750 -4.000 2245.310 2.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1627.550 45.800 1627.870 45.860 ;
        RECT 2262.350 45.800 2262.670 45.860 ;
        RECT 1627.550 45.660 2262.670 45.800 ;
        RECT 1627.550 45.600 1627.870 45.660 ;
        RECT 2262.350 45.600 2262.670 45.660 ;
      LAYER via ;
        RECT 1627.580 45.600 1627.840 45.860 ;
        RECT 2262.380 45.600 2262.640 45.860 ;
      LAYER met2 ;
        RECT 1626.110 1100.650 1626.390 1104.000 ;
        RECT 1626.110 1100.510 1627.780 1100.650 ;
        RECT 1626.110 1100.000 1626.390 1100.510 ;
        RECT 1627.640 45.890 1627.780 1100.510 ;
        RECT 1627.580 45.570 1627.840 45.890 ;
        RECT 2262.380 45.570 2262.640 45.890 ;
        RECT 2262.440 2.000 2262.580 45.570 ;
        RECT 2262.230 -4.000 2262.790 2.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1633.990 45.460 1634.310 45.520 ;
        RECT 2280.290 45.460 2280.610 45.520 ;
        RECT 1633.990 45.320 2280.610 45.460 ;
        RECT 1633.990 45.260 1634.310 45.320 ;
        RECT 2280.290 45.260 2280.610 45.320 ;
      LAYER via ;
        RECT 1634.020 45.260 1634.280 45.520 ;
        RECT 2280.320 45.260 2280.580 45.520 ;
      LAYER met2 ;
        RECT 1632.550 1100.650 1632.830 1104.000 ;
        RECT 1632.550 1100.510 1633.300 1100.650 ;
        RECT 1632.550 1100.000 1632.830 1100.510 ;
        RECT 1633.160 1085.690 1633.300 1100.510 ;
        RECT 1633.160 1085.550 1634.680 1085.690 ;
        RECT 1634.540 980.290 1634.680 1085.550 ;
        RECT 1634.080 980.150 1634.680 980.290 ;
        RECT 1634.080 979.610 1634.220 980.150 ;
        RECT 1634.080 979.470 1634.680 979.610 ;
        RECT 1634.540 835.450 1634.680 979.470 ;
        RECT 1634.080 835.310 1634.680 835.450 ;
        RECT 1634.080 834.770 1634.220 835.310 ;
        RECT 1634.080 834.630 1634.680 834.770 ;
        RECT 1634.540 738.890 1634.680 834.630 ;
        RECT 1634.080 738.750 1634.680 738.890 ;
        RECT 1634.080 738.210 1634.220 738.750 ;
        RECT 1634.080 738.070 1634.680 738.210 ;
        RECT 1634.540 642.330 1634.680 738.070 ;
        RECT 1634.080 642.190 1634.680 642.330 ;
        RECT 1634.080 641.650 1634.220 642.190 ;
        RECT 1634.080 641.510 1634.680 641.650 ;
        RECT 1634.540 545.770 1634.680 641.510 ;
        RECT 1634.080 545.630 1634.680 545.770 ;
        RECT 1634.080 545.090 1634.220 545.630 ;
        RECT 1634.080 544.950 1634.680 545.090 ;
        RECT 1634.540 449.210 1634.680 544.950 ;
        RECT 1634.080 449.070 1634.680 449.210 ;
        RECT 1634.080 448.530 1634.220 449.070 ;
        RECT 1634.080 448.390 1634.680 448.530 ;
        RECT 1634.540 351.970 1634.680 448.390 ;
        RECT 1634.080 351.830 1634.680 351.970 ;
        RECT 1634.080 351.290 1634.220 351.830 ;
        RECT 1634.080 351.150 1634.680 351.290 ;
        RECT 1634.540 255.410 1634.680 351.150 ;
        RECT 1634.080 255.270 1634.680 255.410 ;
        RECT 1634.080 254.730 1634.220 255.270 ;
        RECT 1634.080 254.590 1634.680 254.730 ;
        RECT 1634.540 158.850 1634.680 254.590 ;
        RECT 1634.080 158.710 1634.680 158.850 ;
        RECT 1634.080 158.170 1634.220 158.710 ;
        RECT 1634.080 158.030 1634.680 158.170 ;
        RECT 1634.540 62.290 1634.680 158.030 ;
        RECT 1634.080 62.150 1634.680 62.290 ;
        RECT 1634.080 45.550 1634.220 62.150 ;
        RECT 1634.020 45.230 1634.280 45.550 ;
        RECT 2280.320 45.230 2280.580 45.550 ;
        RECT 2280.380 2.000 2280.520 45.230 ;
        RECT 2280.170 -4.000 2280.730 2.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1640.505 1027.905 1640.675 1055.615 ;
        RECT 1640.965 931.345 1641.135 965.515 ;
        RECT 1641.425 724.625 1641.595 738.395 ;
        RECT 1641.425 620.925 1641.595 641.835 ;
        RECT 1640.505 138.125 1640.675 159.035 ;
        RECT 1640.965 48.365 1641.135 96.475 ;
      LAYER mcon ;
        RECT 1640.505 1055.445 1640.675 1055.615 ;
        RECT 1640.965 965.345 1641.135 965.515 ;
        RECT 1641.425 738.225 1641.595 738.395 ;
        RECT 1641.425 641.665 1641.595 641.835 ;
        RECT 1640.505 158.865 1640.675 159.035 ;
        RECT 1640.965 96.305 1641.135 96.475 ;
      LAYER met1 ;
        RECT 1640.430 1055.600 1640.750 1055.660 ;
        RECT 1640.235 1055.460 1640.750 1055.600 ;
        RECT 1640.430 1055.400 1640.750 1055.460 ;
        RECT 1640.445 1028.060 1640.735 1028.105 ;
        RECT 1640.890 1028.060 1641.210 1028.120 ;
        RECT 1640.445 1027.920 1641.210 1028.060 ;
        RECT 1640.445 1027.875 1640.735 1027.920 ;
        RECT 1640.890 1027.860 1641.210 1027.920 ;
        RECT 1640.905 965.500 1641.195 965.545 ;
        RECT 1641.350 965.500 1641.670 965.560 ;
        RECT 1640.905 965.360 1641.670 965.500 ;
        RECT 1640.905 965.315 1641.195 965.360 ;
        RECT 1641.350 965.300 1641.670 965.360 ;
        RECT 1640.890 931.500 1641.210 931.560 ;
        RECT 1640.695 931.360 1641.210 931.500 ;
        RECT 1640.890 931.300 1641.210 931.360 ;
        RECT 1639.970 845.480 1640.290 845.540 ;
        RECT 1640.890 845.480 1641.210 845.540 ;
        RECT 1639.970 845.340 1641.210 845.480 ;
        RECT 1639.970 845.280 1640.290 845.340 ;
        RECT 1640.890 845.280 1641.210 845.340 ;
        RECT 1640.890 786.800 1641.210 787.060 ;
        RECT 1640.980 786.320 1641.120 786.800 ;
        RECT 1641.350 786.320 1641.670 786.380 ;
        RECT 1640.980 786.180 1641.670 786.320 ;
        RECT 1641.350 786.120 1641.670 786.180 ;
        RECT 1641.350 738.380 1641.670 738.440 ;
        RECT 1641.155 738.240 1641.670 738.380 ;
        RECT 1641.350 738.180 1641.670 738.240 ;
        RECT 1641.350 724.780 1641.670 724.840 ;
        RECT 1641.155 724.640 1641.670 724.780 ;
        RECT 1641.350 724.580 1641.670 724.640 ;
        RECT 1641.350 641.820 1641.670 641.880 ;
        RECT 1641.155 641.680 1641.670 641.820 ;
        RECT 1641.350 641.620 1641.670 641.680 ;
        RECT 1641.350 621.080 1641.670 621.140 ;
        RECT 1641.155 620.940 1641.670 621.080 ;
        RECT 1641.350 620.880 1641.670 620.940 ;
        RECT 1640.890 572.800 1641.210 572.860 ;
        RECT 1641.350 572.800 1641.670 572.860 ;
        RECT 1640.890 572.660 1641.670 572.800 ;
        RECT 1640.890 572.600 1641.210 572.660 ;
        RECT 1641.350 572.600 1641.670 572.660 ;
        RECT 1641.350 545.060 1641.670 545.320 ;
        RECT 1641.440 544.640 1641.580 545.060 ;
        RECT 1641.350 544.380 1641.670 544.640 ;
        RECT 1640.890 289.920 1641.210 289.980 ;
        RECT 1641.350 289.920 1641.670 289.980 ;
        RECT 1640.890 289.780 1641.670 289.920 ;
        RECT 1640.890 289.720 1641.210 289.780 ;
        RECT 1641.350 289.720 1641.670 289.780 ;
        RECT 1639.510 265.780 1639.830 265.840 ;
        RECT 1641.350 265.780 1641.670 265.840 ;
        RECT 1639.510 265.640 1641.670 265.780 ;
        RECT 1639.510 265.580 1639.830 265.640 ;
        RECT 1641.350 265.580 1641.670 265.640 ;
        RECT 1641.350 187.040 1641.670 187.300 ;
        RECT 1641.440 186.620 1641.580 187.040 ;
        RECT 1641.350 186.360 1641.670 186.620 ;
        RECT 1640.445 159.020 1640.735 159.065 ;
        RECT 1640.890 159.020 1641.210 159.080 ;
        RECT 1640.445 158.880 1641.210 159.020 ;
        RECT 1640.445 158.835 1640.735 158.880 ;
        RECT 1640.890 158.820 1641.210 158.880 ;
        RECT 1640.430 138.280 1640.750 138.340 ;
        RECT 1640.235 138.140 1640.750 138.280 ;
        RECT 1640.430 138.080 1640.750 138.140 ;
        RECT 1640.905 96.460 1641.195 96.505 ;
        RECT 1641.350 96.460 1641.670 96.520 ;
        RECT 1640.905 96.320 1641.670 96.460 ;
        RECT 1640.905 96.275 1641.195 96.320 ;
        RECT 1641.350 96.260 1641.670 96.320 ;
        RECT 1640.890 48.520 1641.210 48.580 ;
        RECT 1640.695 48.380 1641.210 48.520 ;
        RECT 1640.890 48.320 1641.210 48.380 ;
        RECT 1640.890 45.120 1641.210 45.180 ;
        RECT 2298.230 45.120 2298.550 45.180 ;
        RECT 1640.890 44.980 2298.550 45.120 ;
        RECT 1640.890 44.920 1641.210 44.980 ;
        RECT 2298.230 44.920 2298.550 44.980 ;
      LAYER via ;
        RECT 1640.460 1055.400 1640.720 1055.660 ;
        RECT 1640.920 1027.860 1641.180 1028.120 ;
        RECT 1641.380 965.300 1641.640 965.560 ;
        RECT 1640.920 931.300 1641.180 931.560 ;
        RECT 1640.000 845.280 1640.260 845.540 ;
        RECT 1640.920 845.280 1641.180 845.540 ;
        RECT 1640.920 786.800 1641.180 787.060 ;
        RECT 1641.380 786.120 1641.640 786.380 ;
        RECT 1641.380 738.180 1641.640 738.440 ;
        RECT 1641.380 724.580 1641.640 724.840 ;
        RECT 1641.380 641.620 1641.640 641.880 ;
        RECT 1641.380 620.880 1641.640 621.140 ;
        RECT 1640.920 572.600 1641.180 572.860 ;
        RECT 1641.380 572.600 1641.640 572.860 ;
        RECT 1641.380 545.060 1641.640 545.320 ;
        RECT 1641.380 544.380 1641.640 544.640 ;
        RECT 1640.920 289.720 1641.180 289.980 ;
        RECT 1641.380 289.720 1641.640 289.980 ;
        RECT 1639.540 265.580 1639.800 265.840 ;
        RECT 1641.380 265.580 1641.640 265.840 ;
        RECT 1641.380 187.040 1641.640 187.300 ;
        RECT 1641.380 186.360 1641.640 186.620 ;
        RECT 1640.920 158.820 1641.180 159.080 ;
        RECT 1640.460 138.080 1640.720 138.340 ;
        RECT 1641.380 96.260 1641.640 96.520 ;
        RECT 1640.920 48.320 1641.180 48.580 ;
        RECT 1640.920 44.920 1641.180 45.180 ;
        RECT 2298.260 44.920 2298.520 45.180 ;
      LAYER met2 ;
        RECT 1638.530 1100.650 1638.810 1104.000 ;
        RECT 1638.530 1100.510 1640.660 1100.650 ;
        RECT 1638.530 1100.000 1638.810 1100.510 ;
        RECT 1640.520 1055.690 1640.660 1100.510 ;
        RECT 1640.460 1055.370 1640.720 1055.690 ;
        RECT 1640.920 1027.830 1641.180 1028.150 ;
        RECT 1640.980 1007.490 1641.120 1027.830 ;
        RECT 1640.980 1007.350 1641.580 1007.490 ;
        RECT 1641.440 965.590 1641.580 1007.350 ;
        RECT 1641.380 965.270 1641.640 965.590 ;
        RECT 1640.920 931.270 1641.180 931.590 ;
        RECT 1640.980 893.930 1641.120 931.270 ;
        RECT 1640.520 893.790 1641.120 893.930 ;
        RECT 1640.520 870.245 1640.660 893.790 ;
        RECT 1640.450 869.875 1640.730 870.245 ;
        RECT 1641.370 869.875 1641.650 870.245 ;
        RECT 1641.440 869.450 1641.580 869.875 ;
        RECT 1640.980 869.310 1641.580 869.450 ;
        RECT 1640.980 845.570 1641.120 869.310 ;
        RECT 1640.000 845.250 1640.260 845.570 ;
        RECT 1640.920 845.250 1641.180 845.570 ;
        RECT 1640.060 821.285 1640.200 845.250 ;
        RECT 1639.990 820.915 1640.270 821.285 ;
        RECT 1640.910 820.915 1641.190 821.285 ;
        RECT 1640.980 787.090 1641.120 820.915 ;
        RECT 1640.920 786.770 1641.180 787.090 ;
        RECT 1641.380 786.090 1641.640 786.410 ;
        RECT 1641.440 738.470 1641.580 786.090 ;
        RECT 1641.380 738.150 1641.640 738.470 ;
        RECT 1641.380 724.550 1641.640 724.870 ;
        RECT 1641.440 641.910 1641.580 724.550 ;
        RECT 1641.380 641.590 1641.640 641.910 ;
        RECT 1641.380 620.850 1641.640 621.170 ;
        RECT 1641.440 620.570 1641.580 620.850 ;
        RECT 1640.980 620.430 1641.580 620.570 ;
        RECT 1640.980 572.890 1641.120 620.430 ;
        RECT 1640.920 572.570 1641.180 572.890 ;
        RECT 1641.380 572.570 1641.640 572.890 ;
        RECT 1641.440 545.350 1641.580 572.570 ;
        RECT 1641.380 545.030 1641.640 545.350 ;
        RECT 1641.380 544.350 1641.640 544.670 ;
        RECT 1641.440 290.770 1641.580 544.350 ;
        RECT 1640.980 290.630 1641.580 290.770 ;
        RECT 1640.980 290.010 1641.120 290.630 ;
        RECT 1640.920 289.690 1641.180 290.010 ;
        RECT 1641.380 289.690 1641.640 290.010 ;
        RECT 1641.440 265.870 1641.580 289.690 ;
        RECT 1639.540 265.550 1639.800 265.870 ;
        RECT 1641.380 265.550 1641.640 265.870 ;
        RECT 1639.600 241.925 1639.740 265.550 ;
        RECT 1639.530 241.555 1639.810 241.925 ;
        RECT 1640.450 241.810 1640.730 241.925 ;
        RECT 1640.450 241.670 1641.120 241.810 ;
        RECT 1640.450 241.555 1640.730 241.670 ;
        RECT 1640.980 210.530 1641.120 241.670 ;
        RECT 1640.980 210.390 1641.580 210.530 ;
        RECT 1641.440 187.330 1641.580 210.390 ;
        RECT 1641.380 187.010 1641.640 187.330 ;
        RECT 1641.380 186.330 1641.640 186.650 ;
        RECT 1641.440 186.050 1641.580 186.330 ;
        RECT 1640.980 185.910 1641.580 186.050 ;
        RECT 1640.980 159.110 1641.120 185.910 ;
        RECT 1640.920 158.790 1641.180 159.110 ;
        RECT 1640.460 138.050 1640.720 138.370 ;
        RECT 1640.520 109.890 1640.660 138.050 ;
        RECT 1640.520 109.750 1641.580 109.890 ;
        RECT 1641.440 96.550 1641.580 109.750 ;
        RECT 1641.380 96.230 1641.640 96.550 ;
        RECT 1640.920 48.290 1641.180 48.610 ;
        RECT 1640.980 45.210 1641.120 48.290 ;
        RECT 1640.920 44.890 1641.180 45.210 ;
        RECT 2298.260 44.890 2298.520 45.210 ;
        RECT 2298.320 2.000 2298.460 44.890 ;
        RECT 2298.110 -4.000 2298.670 2.000 ;
      LAYER via2 ;
        RECT 1640.450 869.920 1640.730 870.200 ;
        RECT 1641.370 869.920 1641.650 870.200 ;
        RECT 1639.990 820.960 1640.270 821.240 ;
        RECT 1640.910 820.960 1641.190 821.240 ;
        RECT 1639.530 241.600 1639.810 241.880 ;
        RECT 1640.450 241.600 1640.730 241.880 ;
      LAYER met3 ;
        RECT 1640.425 870.210 1640.755 870.225 ;
        RECT 1641.345 870.210 1641.675 870.225 ;
        RECT 1640.425 869.910 1641.675 870.210 ;
        RECT 1640.425 869.895 1640.755 869.910 ;
        RECT 1641.345 869.895 1641.675 869.910 ;
        RECT 1639.965 821.250 1640.295 821.265 ;
        RECT 1640.885 821.250 1641.215 821.265 ;
        RECT 1639.965 820.950 1641.215 821.250 ;
        RECT 1639.965 820.935 1640.295 820.950 ;
        RECT 1640.885 820.935 1641.215 820.950 ;
        RECT 1639.505 241.890 1639.835 241.905 ;
        RECT 1640.425 241.890 1640.755 241.905 ;
        RECT 1639.505 241.590 1640.755 241.890 ;
        RECT 1639.505 241.575 1639.835 241.590 ;
        RECT 1640.425 241.575 1640.755 241.590 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1646.945 1007.165 1647.115 1048.815 ;
        RECT 1647.865 907.885 1648.035 959.055 ;
        RECT 1647.865 676.345 1648.035 724.455 ;
        RECT 1647.865 579.785 1648.035 627.895 ;
        RECT 1647.865 483.225 1648.035 531.335 ;
        RECT 1647.865 282.965 1648.035 331.075 ;
        RECT 1646.945 186.405 1647.115 210.715 ;
        RECT 1647.405 96.645 1647.575 144.755 ;
        RECT 1647.405 48.365 1647.575 62.475 ;
      LAYER mcon ;
        RECT 1646.945 1048.645 1647.115 1048.815 ;
        RECT 1647.865 958.885 1648.035 959.055 ;
        RECT 1647.865 724.285 1648.035 724.455 ;
        RECT 1647.865 627.725 1648.035 627.895 ;
        RECT 1647.865 531.165 1648.035 531.335 ;
        RECT 1647.865 330.905 1648.035 331.075 ;
        RECT 1646.945 210.545 1647.115 210.715 ;
        RECT 1647.405 144.585 1647.575 144.755 ;
        RECT 1647.405 62.305 1647.575 62.475 ;
      LAYER met1 ;
        RECT 1646.870 1048.800 1647.190 1048.860 ;
        RECT 1646.675 1048.660 1647.190 1048.800 ;
        RECT 1646.870 1048.600 1647.190 1048.660 ;
        RECT 1646.885 1007.320 1647.175 1007.365 ;
        RECT 1647.330 1007.320 1647.650 1007.380 ;
        RECT 1646.885 1007.180 1647.650 1007.320 ;
        RECT 1646.885 1007.135 1647.175 1007.180 ;
        RECT 1647.330 1007.120 1647.650 1007.180 ;
        RECT 1647.790 959.040 1648.110 959.100 ;
        RECT 1647.595 958.900 1648.110 959.040 ;
        RECT 1647.790 958.840 1648.110 958.900 ;
        RECT 1646.870 908.040 1647.190 908.100 ;
        RECT 1647.805 908.040 1648.095 908.085 ;
        RECT 1646.870 907.900 1648.095 908.040 ;
        RECT 1646.870 907.840 1647.190 907.900 ;
        RECT 1647.805 907.855 1648.095 907.900 ;
        RECT 1646.870 869.620 1647.190 869.680 ;
        RECT 1647.790 869.620 1648.110 869.680 ;
        RECT 1646.870 869.480 1648.110 869.620 ;
        RECT 1646.870 869.420 1647.190 869.480 ;
        RECT 1647.790 869.420 1648.110 869.480 ;
        RECT 1646.410 845.480 1646.730 845.540 ;
        RECT 1647.330 845.480 1647.650 845.540 ;
        RECT 1646.410 845.340 1647.650 845.480 ;
        RECT 1646.410 845.280 1646.730 845.340 ;
        RECT 1647.330 845.280 1647.650 845.340 ;
        RECT 1647.330 786.800 1647.650 787.060 ;
        RECT 1647.420 786.320 1647.560 786.800 ;
        RECT 1647.790 786.320 1648.110 786.380 ;
        RECT 1647.420 786.180 1648.110 786.320 ;
        RECT 1647.790 786.120 1648.110 786.180 ;
        RECT 1647.790 724.440 1648.110 724.500 ;
        RECT 1647.595 724.300 1648.110 724.440 ;
        RECT 1647.790 724.240 1648.110 724.300 ;
        RECT 1647.790 676.500 1648.110 676.560 ;
        RECT 1647.595 676.360 1648.110 676.500 ;
        RECT 1647.790 676.300 1648.110 676.360 ;
        RECT 1647.790 627.880 1648.110 627.940 ;
        RECT 1647.595 627.740 1648.110 627.880 ;
        RECT 1647.790 627.680 1648.110 627.740 ;
        RECT 1647.790 579.940 1648.110 580.000 ;
        RECT 1647.595 579.800 1648.110 579.940 ;
        RECT 1647.790 579.740 1648.110 579.800 ;
        RECT 1647.790 531.320 1648.110 531.380 ;
        RECT 1647.595 531.180 1648.110 531.320 ;
        RECT 1647.790 531.120 1648.110 531.180 ;
        RECT 1647.790 483.380 1648.110 483.440 ;
        RECT 1647.595 483.240 1648.110 483.380 ;
        RECT 1647.790 483.180 1648.110 483.240 ;
        RECT 1647.790 338.680 1648.110 338.940 ;
        RECT 1647.880 338.260 1648.020 338.680 ;
        RECT 1647.790 338.000 1648.110 338.260 ;
        RECT 1647.790 331.060 1648.110 331.120 ;
        RECT 1647.595 330.920 1648.110 331.060 ;
        RECT 1647.790 330.860 1648.110 330.920 ;
        RECT 1647.790 283.120 1648.110 283.180 ;
        RECT 1647.595 282.980 1648.110 283.120 ;
        RECT 1647.790 282.920 1648.110 282.980 ;
        RECT 1646.885 210.700 1647.175 210.745 ;
        RECT 1647.330 210.700 1647.650 210.760 ;
        RECT 1646.885 210.560 1647.650 210.700 ;
        RECT 1646.885 210.515 1647.175 210.560 ;
        RECT 1647.330 210.500 1647.650 210.560 ;
        RECT 1646.870 186.560 1647.190 186.620 ;
        RECT 1646.675 186.420 1647.190 186.560 ;
        RECT 1646.870 186.360 1647.190 186.420 ;
        RECT 1647.330 144.740 1647.650 144.800 ;
        RECT 1647.135 144.600 1647.650 144.740 ;
        RECT 1647.330 144.540 1647.650 144.600 ;
        RECT 1647.345 96.800 1647.635 96.845 ;
        RECT 1647.790 96.800 1648.110 96.860 ;
        RECT 1647.345 96.660 1648.110 96.800 ;
        RECT 1647.345 96.615 1647.635 96.660 ;
        RECT 1647.790 96.600 1648.110 96.660 ;
        RECT 1647.330 62.460 1647.650 62.520 ;
        RECT 1647.135 62.320 1647.650 62.460 ;
        RECT 1647.330 62.260 1647.650 62.320 ;
        RECT 1647.330 48.520 1647.650 48.580 ;
        RECT 1647.135 48.380 1647.650 48.520 ;
        RECT 1647.330 48.320 1647.650 48.380 ;
        RECT 1647.330 44.780 1647.650 44.840 ;
        RECT 2316.170 44.780 2316.490 44.840 ;
        RECT 1647.330 44.640 2316.490 44.780 ;
        RECT 1647.330 44.580 1647.650 44.640 ;
        RECT 2316.170 44.580 2316.490 44.640 ;
      LAYER via ;
        RECT 1646.900 1048.600 1647.160 1048.860 ;
        RECT 1647.360 1007.120 1647.620 1007.380 ;
        RECT 1647.820 958.840 1648.080 959.100 ;
        RECT 1646.900 907.840 1647.160 908.100 ;
        RECT 1646.900 869.420 1647.160 869.680 ;
        RECT 1647.820 869.420 1648.080 869.680 ;
        RECT 1646.440 845.280 1646.700 845.540 ;
        RECT 1647.360 845.280 1647.620 845.540 ;
        RECT 1647.360 786.800 1647.620 787.060 ;
        RECT 1647.820 786.120 1648.080 786.380 ;
        RECT 1647.820 724.240 1648.080 724.500 ;
        RECT 1647.820 676.300 1648.080 676.560 ;
        RECT 1647.820 627.680 1648.080 627.940 ;
        RECT 1647.820 579.740 1648.080 580.000 ;
        RECT 1647.820 531.120 1648.080 531.380 ;
        RECT 1647.820 483.180 1648.080 483.440 ;
        RECT 1647.820 338.680 1648.080 338.940 ;
        RECT 1647.820 338.000 1648.080 338.260 ;
        RECT 1647.820 330.860 1648.080 331.120 ;
        RECT 1647.820 282.920 1648.080 283.180 ;
        RECT 1647.360 210.500 1647.620 210.760 ;
        RECT 1646.900 186.360 1647.160 186.620 ;
        RECT 1647.360 144.540 1647.620 144.800 ;
        RECT 1647.820 96.600 1648.080 96.860 ;
        RECT 1647.360 62.260 1647.620 62.520 ;
        RECT 1647.360 48.320 1647.620 48.580 ;
        RECT 1647.360 44.580 1647.620 44.840 ;
        RECT 2316.200 44.580 2316.460 44.840 ;
      LAYER met2 ;
        RECT 1644.510 1100.650 1644.790 1104.000 ;
        RECT 1644.510 1100.510 1646.180 1100.650 ;
        RECT 1644.510 1100.000 1644.790 1100.510 ;
        RECT 1646.040 1088.410 1646.180 1100.510 ;
        RECT 1646.040 1088.270 1647.100 1088.410 ;
        RECT 1646.960 1048.890 1647.100 1088.270 ;
        RECT 1646.900 1048.570 1647.160 1048.890 ;
        RECT 1647.360 1007.090 1647.620 1007.410 ;
        RECT 1647.420 1000.690 1647.560 1007.090 ;
        RECT 1647.420 1000.550 1648.020 1000.690 ;
        RECT 1647.880 959.130 1648.020 1000.550 ;
        RECT 1647.820 958.810 1648.080 959.130 ;
        RECT 1646.900 907.810 1647.160 908.130 ;
        RECT 1646.960 869.710 1647.100 907.810 ;
        RECT 1646.900 869.390 1647.160 869.710 ;
        RECT 1647.820 869.450 1648.080 869.710 ;
        RECT 1647.420 869.390 1648.080 869.450 ;
        RECT 1647.420 869.310 1648.020 869.390 ;
        RECT 1647.420 845.570 1647.560 869.310 ;
        RECT 1646.440 845.250 1646.700 845.570 ;
        RECT 1647.360 845.250 1647.620 845.570 ;
        RECT 1646.500 821.285 1646.640 845.250 ;
        RECT 1646.430 820.915 1646.710 821.285 ;
        RECT 1647.350 820.915 1647.630 821.285 ;
        RECT 1647.420 787.090 1647.560 820.915 ;
        RECT 1647.360 786.770 1647.620 787.090 ;
        RECT 1647.820 786.090 1648.080 786.410 ;
        RECT 1647.880 739.005 1648.020 786.090 ;
        RECT 1647.810 738.635 1648.090 739.005 ;
        RECT 1647.810 724.355 1648.090 724.725 ;
        RECT 1647.820 724.210 1648.080 724.355 ;
        RECT 1647.820 676.270 1648.080 676.590 ;
        RECT 1647.880 642.445 1648.020 676.270 ;
        RECT 1647.810 642.075 1648.090 642.445 ;
        RECT 1647.810 627.795 1648.090 628.165 ;
        RECT 1647.820 627.650 1648.080 627.795 ;
        RECT 1647.820 579.710 1648.080 580.030 ;
        RECT 1647.880 545.885 1648.020 579.710 ;
        RECT 1647.810 545.515 1648.090 545.885 ;
        RECT 1647.810 531.235 1648.090 531.605 ;
        RECT 1647.820 531.090 1648.080 531.235 ;
        RECT 1647.820 483.150 1648.080 483.470 ;
        RECT 1647.880 338.970 1648.020 483.150 ;
        RECT 1647.820 338.650 1648.080 338.970 ;
        RECT 1647.820 337.970 1648.080 338.290 ;
        RECT 1647.880 331.150 1648.020 337.970 ;
        RECT 1647.820 330.830 1648.080 331.150 ;
        RECT 1647.820 282.890 1648.080 283.210 ;
        RECT 1647.880 256.205 1648.020 282.890 ;
        RECT 1647.810 255.835 1648.090 256.205 ;
        RECT 1647.350 241.555 1647.630 241.925 ;
        RECT 1647.420 210.790 1647.560 241.555 ;
        RECT 1647.360 210.470 1647.620 210.790 ;
        RECT 1646.900 186.330 1647.160 186.650 ;
        RECT 1646.960 145.250 1647.100 186.330 ;
        RECT 1646.960 145.110 1647.560 145.250 ;
        RECT 1647.420 144.830 1647.560 145.110 ;
        RECT 1647.360 144.510 1647.620 144.830 ;
        RECT 1647.820 96.570 1648.080 96.890 ;
        RECT 1647.880 96.290 1648.020 96.570 ;
        RECT 1647.420 96.150 1648.020 96.290 ;
        RECT 1647.420 62.550 1647.560 96.150 ;
        RECT 1647.360 62.230 1647.620 62.550 ;
        RECT 1647.360 48.290 1647.620 48.610 ;
        RECT 1647.420 44.870 1647.560 48.290 ;
        RECT 1647.360 44.550 1647.620 44.870 ;
        RECT 2316.200 44.550 2316.460 44.870 ;
        RECT 2316.260 2.000 2316.400 44.550 ;
        RECT 2316.050 -4.000 2316.610 2.000 ;
      LAYER via2 ;
        RECT 1646.430 820.960 1646.710 821.240 ;
        RECT 1647.350 820.960 1647.630 821.240 ;
        RECT 1647.810 738.680 1648.090 738.960 ;
        RECT 1647.810 724.400 1648.090 724.680 ;
        RECT 1647.810 642.120 1648.090 642.400 ;
        RECT 1647.810 627.840 1648.090 628.120 ;
        RECT 1647.810 545.560 1648.090 545.840 ;
        RECT 1647.810 531.280 1648.090 531.560 ;
        RECT 1647.810 255.880 1648.090 256.160 ;
        RECT 1647.350 241.600 1647.630 241.880 ;
      LAYER met3 ;
        RECT 1646.405 821.250 1646.735 821.265 ;
        RECT 1647.325 821.250 1647.655 821.265 ;
        RECT 1646.405 820.950 1647.655 821.250 ;
        RECT 1646.405 820.935 1646.735 820.950 ;
        RECT 1647.325 820.935 1647.655 820.950 ;
        RECT 1647.785 738.980 1648.115 738.985 ;
        RECT 1647.785 738.970 1648.370 738.980 ;
        RECT 1647.785 738.670 1648.570 738.970 ;
        RECT 1647.785 738.660 1648.370 738.670 ;
        RECT 1647.785 738.655 1648.115 738.660 ;
        RECT 1647.785 724.700 1648.115 724.705 ;
        RECT 1647.785 724.690 1648.370 724.700 ;
        RECT 1647.785 724.390 1648.570 724.690 ;
        RECT 1647.785 724.380 1648.370 724.390 ;
        RECT 1647.785 724.375 1648.115 724.380 ;
        RECT 1647.785 642.420 1648.115 642.425 ;
        RECT 1647.785 642.410 1648.370 642.420 ;
        RECT 1647.785 642.110 1648.570 642.410 ;
        RECT 1647.785 642.100 1648.370 642.110 ;
        RECT 1647.785 642.095 1648.115 642.100 ;
        RECT 1647.785 628.140 1648.115 628.145 ;
        RECT 1647.785 628.130 1648.370 628.140 ;
        RECT 1647.785 627.830 1648.570 628.130 ;
        RECT 1647.785 627.820 1648.370 627.830 ;
        RECT 1647.785 627.815 1648.115 627.820 ;
        RECT 1647.785 545.860 1648.115 545.865 ;
        RECT 1647.785 545.850 1648.370 545.860 ;
        RECT 1647.785 545.550 1648.570 545.850 ;
        RECT 1647.785 545.540 1648.370 545.550 ;
        RECT 1647.785 545.535 1648.115 545.540 ;
        RECT 1647.785 531.580 1648.115 531.585 ;
        RECT 1647.785 531.570 1648.370 531.580 ;
        RECT 1647.785 531.270 1648.570 531.570 ;
        RECT 1647.785 531.260 1648.370 531.270 ;
        RECT 1647.785 531.255 1648.115 531.260 ;
        RECT 1647.070 256.170 1647.450 256.180 ;
        RECT 1647.785 256.170 1648.115 256.185 ;
        RECT 1647.070 255.870 1648.115 256.170 ;
        RECT 1647.070 255.860 1647.450 255.870 ;
        RECT 1647.785 255.855 1648.115 255.870 ;
        RECT 1647.325 241.900 1647.655 241.905 ;
        RECT 1647.070 241.890 1647.655 241.900 ;
        RECT 1647.070 241.590 1647.880 241.890 ;
        RECT 1647.070 241.580 1647.655 241.590 ;
        RECT 1647.325 241.575 1647.655 241.580 ;
      LAYER via3 ;
        RECT 1648.020 738.660 1648.340 738.980 ;
        RECT 1648.020 724.380 1648.340 724.700 ;
        RECT 1648.020 642.100 1648.340 642.420 ;
        RECT 1648.020 627.820 1648.340 628.140 ;
        RECT 1648.020 545.540 1648.340 545.860 ;
        RECT 1648.020 531.260 1648.340 531.580 ;
        RECT 1647.100 255.860 1647.420 256.180 ;
        RECT 1647.100 241.580 1647.420 241.900 ;
      LAYER met4 ;
        RECT 1648.015 738.655 1648.345 738.985 ;
        RECT 1648.030 724.705 1648.330 738.655 ;
        RECT 1648.015 724.375 1648.345 724.705 ;
        RECT 1648.015 642.095 1648.345 642.425 ;
        RECT 1648.030 628.145 1648.330 642.095 ;
        RECT 1648.015 627.815 1648.345 628.145 ;
        RECT 1648.015 545.535 1648.345 545.865 ;
        RECT 1648.030 531.585 1648.330 545.535 ;
        RECT 1648.015 531.255 1648.345 531.585 ;
        RECT 1647.095 255.855 1647.425 256.185 ;
        RECT 1647.110 241.905 1647.410 255.855 ;
        RECT 1647.095 241.575 1647.425 241.905 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1651.010 1087.900 1651.330 1087.960 ;
        RECT 1655.150 1087.900 1655.470 1087.960 ;
        RECT 1651.010 1087.760 1655.470 1087.900 ;
        RECT 1651.010 1087.700 1651.330 1087.760 ;
        RECT 1655.150 1087.700 1655.470 1087.760 ;
      LAYER via ;
        RECT 1651.040 1087.700 1651.300 1087.960 ;
        RECT 1655.180 1087.700 1655.440 1087.960 ;
      LAYER met2 ;
        RECT 1650.950 1100.580 1651.230 1104.000 ;
        RECT 1650.950 1100.000 1651.240 1100.580 ;
        RECT 1651.100 1087.990 1651.240 1100.000 ;
        RECT 1651.040 1087.670 1651.300 1087.990 ;
        RECT 1655.180 1087.670 1655.440 1087.990 ;
        RECT 1655.240 44.725 1655.380 1087.670 ;
        RECT 1655.170 44.355 1655.450 44.725 ;
        RECT 2334.130 44.355 2334.410 44.725 ;
        RECT 2334.200 2.000 2334.340 44.355 ;
        RECT 2333.990 -4.000 2334.550 2.000 ;
      LAYER via2 ;
        RECT 1655.170 44.400 1655.450 44.680 ;
        RECT 2334.130 44.400 2334.410 44.680 ;
      LAYER met3 ;
        RECT 1655.145 44.690 1655.475 44.705 ;
        RECT 2334.105 44.690 2334.435 44.705 ;
        RECT 1655.145 44.390 2334.435 44.690 ;
        RECT 1655.145 44.375 1655.475 44.390 ;
        RECT 2334.105 44.375 2334.435 44.390 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1656.990 1088.580 1657.310 1088.640 ;
        RECT 1662.050 1088.580 1662.370 1088.640 ;
        RECT 1656.990 1088.440 1662.370 1088.580 ;
        RECT 1656.990 1088.380 1657.310 1088.440 ;
        RECT 1662.050 1088.380 1662.370 1088.440 ;
        RECT 1662.050 62.120 1662.370 62.180 ;
        RECT 2346.070 62.120 2346.390 62.180 ;
        RECT 1662.050 61.980 2346.390 62.120 ;
        RECT 1662.050 61.920 1662.370 61.980 ;
        RECT 2346.070 61.920 2346.390 61.980 ;
      LAYER via ;
        RECT 1657.020 1088.380 1657.280 1088.640 ;
        RECT 1662.080 1088.380 1662.340 1088.640 ;
        RECT 1662.080 61.920 1662.340 62.180 ;
        RECT 2346.100 61.920 2346.360 62.180 ;
      LAYER met2 ;
        RECT 1656.930 1100.580 1657.210 1104.000 ;
        RECT 1656.930 1100.000 1657.220 1100.580 ;
        RECT 1657.080 1088.670 1657.220 1100.000 ;
        RECT 1657.020 1088.350 1657.280 1088.670 ;
        RECT 1662.080 1088.350 1662.340 1088.670 ;
        RECT 1662.140 62.210 1662.280 1088.350 ;
        RECT 1662.080 61.890 1662.340 62.210 ;
        RECT 2346.100 61.890 2346.360 62.210 ;
        RECT 2346.160 16.730 2346.300 61.890 ;
        RECT 2346.160 16.590 2351.820 16.730 ;
        RECT 2351.680 2.000 2351.820 16.590 ;
        RECT 2351.470 -4.000 2352.030 2.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1662.970 1087.220 1663.290 1087.280 ;
        RECT 1668.490 1087.220 1668.810 1087.280 ;
        RECT 1662.970 1087.080 1668.810 1087.220 ;
        RECT 1662.970 1087.020 1663.290 1087.080 ;
        RECT 1668.490 1087.020 1668.810 1087.080 ;
        RECT 1668.490 61.780 1668.810 61.840 ;
        RECT 2366.770 61.780 2367.090 61.840 ;
        RECT 1668.490 61.640 2367.090 61.780 ;
        RECT 1668.490 61.580 1668.810 61.640 ;
        RECT 2366.770 61.580 2367.090 61.640 ;
      LAYER via ;
        RECT 1663.000 1087.020 1663.260 1087.280 ;
        RECT 1668.520 1087.020 1668.780 1087.280 ;
        RECT 1668.520 61.580 1668.780 61.840 ;
        RECT 2366.800 61.580 2367.060 61.840 ;
      LAYER met2 ;
        RECT 1662.910 1100.580 1663.190 1104.000 ;
        RECT 1662.910 1100.000 1663.200 1100.580 ;
        RECT 1663.060 1087.310 1663.200 1100.000 ;
        RECT 1663.000 1086.990 1663.260 1087.310 ;
        RECT 1668.520 1086.990 1668.780 1087.310 ;
        RECT 1668.580 61.870 1668.720 1086.990 ;
        RECT 1668.520 61.550 1668.780 61.870 ;
        RECT 2366.800 61.550 2367.060 61.870 ;
        RECT 2366.860 2.450 2367.000 61.550 ;
        RECT 2366.860 2.310 2369.760 2.450 ;
        RECT 2369.620 2.000 2369.760 2.310 ;
        RECT 2369.410 -4.000 2369.970 2.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1668.030 63.480 1668.350 63.540 ;
        RECT 2387.930 63.480 2388.250 63.540 ;
        RECT 1668.030 63.340 2388.250 63.480 ;
        RECT 1668.030 63.280 1668.350 63.340 ;
        RECT 2387.930 63.280 2388.250 63.340 ;
      LAYER via ;
        RECT 1668.060 63.280 1668.320 63.540 ;
        RECT 2387.960 63.280 2388.220 63.540 ;
      LAYER met2 ;
        RECT 1669.350 1100.650 1669.630 1104.000 ;
        RECT 1668.120 1100.510 1669.630 1100.650 ;
        RECT 1668.120 63.570 1668.260 1100.510 ;
        RECT 1669.350 1100.000 1669.630 1100.510 ;
        RECT 1668.060 63.250 1668.320 63.570 ;
        RECT 2387.960 63.250 2388.220 63.570 ;
        RECT 2388.020 17.410 2388.160 63.250 ;
        RECT 2387.560 17.270 2388.160 17.410 ;
        RECT 2387.560 2.000 2387.700 17.270 ;
        RECT 2387.350 -4.000 2387.910 2.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1675.850 63.820 1676.170 63.880 ;
        RECT 2401.270 63.820 2401.590 63.880 ;
        RECT 1675.850 63.680 2401.590 63.820 ;
        RECT 1675.850 63.620 1676.170 63.680 ;
        RECT 2401.270 63.620 2401.590 63.680 ;
      LAYER via ;
        RECT 1675.880 63.620 1676.140 63.880 ;
        RECT 2401.300 63.620 2401.560 63.880 ;
      LAYER met2 ;
        RECT 1675.330 1100.650 1675.610 1104.000 ;
        RECT 1675.330 1100.510 1676.080 1100.650 ;
        RECT 1675.330 1100.000 1675.610 1100.510 ;
        RECT 1675.940 63.910 1676.080 1100.510 ;
        RECT 1675.880 63.590 1676.140 63.910 ;
        RECT 2401.300 63.590 2401.560 63.910 ;
        RECT 2401.360 16.730 2401.500 63.590 ;
        RECT 2401.360 16.590 2405.640 16.730 ;
        RECT 2405.500 2.000 2405.640 16.590 ;
        RECT 2405.290 -4.000 2405.850 2.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1120.245 862.665 1120.415 910.775 ;
        RECT 1120.245 476.085 1120.415 497.675 ;
      LAYER mcon ;
        RECT 1120.245 910.605 1120.415 910.775 ;
        RECT 1120.245 497.505 1120.415 497.675 ;
      LAYER met1 ;
        RECT 1120.170 1089.940 1120.490 1090.000 ;
        RECT 1122.930 1089.940 1123.250 1090.000 ;
        RECT 1120.170 1089.800 1123.250 1089.940 ;
        RECT 1120.170 1089.740 1120.490 1089.800 ;
        RECT 1122.930 1089.740 1123.250 1089.800 ;
        RECT 1119.710 931.640 1120.030 931.900 ;
        RECT 1119.800 931.160 1119.940 931.640 ;
        RECT 1120.170 931.160 1120.490 931.220 ;
        RECT 1119.800 931.020 1120.490 931.160 ;
        RECT 1120.170 930.960 1120.490 931.020 ;
        RECT 1120.170 910.760 1120.490 910.820 ;
        RECT 1119.975 910.620 1120.490 910.760 ;
        RECT 1120.170 910.560 1120.490 910.620 ;
        RECT 1120.170 862.820 1120.490 862.880 ;
        RECT 1119.975 862.680 1120.490 862.820 ;
        RECT 1120.170 862.620 1120.490 862.680 ;
        RECT 1120.170 724.780 1120.490 724.840 ;
        RECT 1120.630 724.780 1120.950 724.840 ;
        RECT 1120.170 724.640 1120.950 724.780 ;
        RECT 1120.170 724.580 1120.490 724.640 ;
        RECT 1120.630 724.580 1120.950 724.640 ;
        RECT 1120.170 497.660 1120.490 497.720 ;
        RECT 1119.975 497.520 1120.490 497.660 ;
        RECT 1120.170 497.460 1120.490 497.520 ;
        RECT 1120.185 476.240 1120.475 476.285 ;
        RECT 1120.630 476.240 1120.950 476.300 ;
        RECT 1120.185 476.100 1120.950 476.240 ;
        RECT 1120.185 476.055 1120.475 476.100 ;
        RECT 1120.630 476.040 1120.950 476.100 ;
        RECT 1120.170 427.960 1120.490 428.020 ;
        RECT 1120.630 427.960 1120.950 428.020 ;
        RECT 1120.170 427.820 1120.950 427.960 ;
        RECT 1120.170 427.760 1120.490 427.820 ;
        RECT 1120.630 427.760 1120.950 427.820 ;
        RECT 1120.170 386.820 1120.490 386.880 ;
        RECT 1119.800 386.680 1120.490 386.820 ;
        RECT 1119.800 386.200 1119.940 386.680 ;
        RECT 1120.170 386.620 1120.490 386.680 ;
        RECT 1119.710 385.940 1120.030 386.200 ;
        RECT 1119.710 337.660 1120.030 337.920 ;
        RECT 1119.800 337.520 1119.940 337.660 ;
        RECT 1120.170 337.520 1120.490 337.580 ;
        RECT 1119.800 337.380 1120.490 337.520 ;
        RECT 1120.170 337.320 1120.490 337.380 ;
        RECT 1120.170 255.380 1120.490 255.640 ;
        RECT 1120.260 254.960 1120.400 255.380 ;
        RECT 1120.170 254.700 1120.490 254.960 ;
        RECT 1119.710 96.800 1120.030 96.860 ;
        RECT 1120.170 96.800 1120.490 96.860 ;
        RECT 1119.710 96.660 1120.490 96.800 ;
        RECT 1119.710 96.600 1120.030 96.660 ;
        RECT 1120.170 96.600 1120.490 96.660 ;
        RECT 799.550 28.460 799.870 28.520 ;
        RECT 1120.170 28.460 1120.490 28.520 ;
        RECT 799.550 28.320 1120.490 28.460 ;
        RECT 799.550 28.260 799.870 28.320 ;
        RECT 1120.170 28.260 1120.490 28.320 ;
      LAYER via ;
        RECT 1120.200 1089.740 1120.460 1090.000 ;
        RECT 1122.960 1089.740 1123.220 1090.000 ;
        RECT 1119.740 931.640 1120.000 931.900 ;
        RECT 1120.200 930.960 1120.460 931.220 ;
        RECT 1120.200 910.560 1120.460 910.820 ;
        RECT 1120.200 862.620 1120.460 862.880 ;
        RECT 1120.200 724.580 1120.460 724.840 ;
        RECT 1120.660 724.580 1120.920 724.840 ;
        RECT 1120.200 497.460 1120.460 497.720 ;
        RECT 1120.660 476.040 1120.920 476.300 ;
        RECT 1120.200 427.760 1120.460 428.020 ;
        RECT 1120.660 427.760 1120.920 428.020 ;
        RECT 1120.200 386.620 1120.460 386.880 ;
        RECT 1119.740 385.940 1120.000 386.200 ;
        RECT 1119.740 337.660 1120.000 337.920 ;
        RECT 1120.200 337.320 1120.460 337.580 ;
        RECT 1120.200 255.380 1120.460 255.640 ;
        RECT 1120.200 254.700 1120.460 254.960 ;
        RECT 1119.740 96.600 1120.000 96.860 ;
        RECT 1120.200 96.600 1120.460 96.860 ;
        RECT 799.580 28.260 799.840 28.520 ;
        RECT 1120.200 28.260 1120.460 28.520 ;
      LAYER met2 ;
        RECT 1124.250 1100.650 1124.530 1104.000 ;
        RECT 1123.020 1100.510 1124.530 1100.650 ;
        RECT 1123.020 1090.030 1123.160 1100.510 ;
        RECT 1124.250 1100.000 1124.530 1100.510 ;
        RECT 1120.200 1089.710 1120.460 1090.030 ;
        RECT 1122.960 1089.710 1123.220 1090.030 ;
        RECT 1120.260 980.290 1120.400 1089.710 ;
        RECT 1119.800 980.150 1120.400 980.290 ;
        RECT 1119.800 931.930 1119.940 980.150 ;
        RECT 1119.740 931.610 1120.000 931.930 ;
        RECT 1120.200 930.930 1120.460 931.250 ;
        RECT 1120.260 910.850 1120.400 930.930 ;
        RECT 1120.200 910.530 1120.460 910.850 ;
        RECT 1120.200 862.590 1120.460 862.910 ;
        RECT 1120.260 789.890 1120.400 862.590 ;
        RECT 1120.260 789.750 1121.320 789.890 ;
        RECT 1121.180 772.210 1121.320 789.750 ;
        RECT 1120.720 772.070 1121.320 772.210 ;
        RECT 1120.720 724.870 1120.860 772.070 ;
        RECT 1120.200 724.550 1120.460 724.870 ;
        RECT 1120.660 724.550 1120.920 724.870 ;
        RECT 1120.260 691.970 1120.400 724.550 ;
        RECT 1120.260 691.830 1121.320 691.970 ;
        RECT 1121.180 669.645 1121.320 691.830 ;
        RECT 1120.190 669.275 1120.470 669.645 ;
        RECT 1121.110 669.275 1121.390 669.645 ;
        RECT 1120.260 594.050 1120.400 669.275 ;
        RECT 1120.260 593.910 1120.860 594.050 ;
        RECT 1120.720 589.970 1120.860 593.910 ;
        RECT 1120.260 589.830 1120.860 589.970 ;
        RECT 1120.260 497.750 1120.400 589.830 ;
        RECT 1120.200 497.430 1120.460 497.750 ;
        RECT 1120.660 476.010 1120.920 476.330 ;
        RECT 1120.720 428.050 1120.860 476.010 ;
        RECT 1120.200 427.730 1120.460 428.050 ;
        RECT 1120.660 427.730 1120.920 428.050 ;
        RECT 1120.260 386.910 1120.400 427.730 ;
        RECT 1120.200 386.590 1120.460 386.910 ;
        RECT 1119.740 385.910 1120.000 386.230 ;
        RECT 1119.800 337.950 1119.940 385.910 ;
        RECT 1119.740 337.630 1120.000 337.950 ;
        RECT 1120.200 337.290 1120.460 337.610 ;
        RECT 1120.260 255.670 1120.400 337.290 ;
        RECT 1120.200 255.350 1120.460 255.670 ;
        RECT 1120.200 254.670 1120.460 254.990 ;
        RECT 1120.260 144.570 1120.400 254.670 ;
        RECT 1119.800 144.430 1120.400 144.570 ;
        RECT 1119.800 96.890 1119.940 144.430 ;
        RECT 1119.740 96.570 1120.000 96.890 ;
        RECT 1120.200 96.570 1120.460 96.890 ;
        RECT 1120.260 28.550 1120.400 96.570 ;
        RECT 799.580 28.230 799.840 28.550 ;
        RECT 1120.200 28.230 1120.460 28.550 ;
        RECT 799.640 2.000 799.780 28.230 ;
        RECT 799.430 -4.000 799.990 2.000 ;
      LAYER via2 ;
        RECT 1120.190 669.320 1120.470 669.600 ;
        RECT 1121.110 669.320 1121.390 669.600 ;
      LAYER met3 ;
        RECT 1120.165 669.610 1120.495 669.625 ;
        RECT 1121.085 669.610 1121.415 669.625 ;
        RECT 1120.165 669.310 1121.415 669.610 ;
        RECT 1120.165 669.295 1120.495 669.310 ;
        RECT 1121.085 669.295 1121.415 669.310 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 644.990 34.240 645.310 34.300 ;
        RECT 1069.570 34.240 1069.890 34.300 ;
        RECT 644.990 34.100 1069.890 34.240 ;
        RECT 644.990 34.040 645.310 34.100 ;
        RECT 1069.570 34.040 1069.890 34.100 ;
      LAYER via ;
        RECT 645.020 34.040 645.280 34.300 ;
        RECT 1069.600 34.040 1069.860 34.300 ;
      LAYER met2 ;
        RECT 1071.350 1100.650 1071.630 1104.000 ;
        RECT 1069.660 1100.510 1071.630 1100.650 ;
        RECT 1069.660 34.330 1069.800 1100.510 ;
        RECT 1071.350 1100.000 1071.630 1100.510 ;
        RECT 645.020 34.010 645.280 34.330 ;
        RECT 1069.600 34.010 1069.860 34.330 ;
        RECT 645.080 2.000 645.220 34.010 ;
        RECT 644.870 -4.000 645.430 2.000 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1683.670 1089.260 1683.990 1089.320 ;
        RECT 1688.730 1089.260 1689.050 1089.320 ;
        RECT 1683.670 1089.120 1689.050 1089.260 ;
        RECT 1683.670 1089.060 1683.990 1089.120 ;
        RECT 1688.730 1089.060 1689.050 1089.120 ;
        RECT 1688.730 64.160 1689.050 64.220 ;
        RECT 2428.870 64.160 2429.190 64.220 ;
        RECT 1688.730 64.020 2429.190 64.160 ;
        RECT 1688.730 63.960 1689.050 64.020 ;
        RECT 2428.870 63.960 2429.190 64.020 ;
      LAYER via ;
        RECT 1683.700 1089.060 1683.960 1089.320 ;
        RECT 1688.760 1089.060 1689.020 1089.320 ;
        RECT 1688.760 63.960 1689.020 64.220 ;
        RECT 2428.900 63.960 2429.160 64.220 ;
      LAYER met2 ;
        RECT 1683.610 1100.580 1683.890 1104.000 ;
        RECT 1683.610 1100.000 1683.900 1100.580 ;
        RECT 1683.760 1089.350 1683.900 1100.000 ;
        RECT 1683.700 1089.030 1683.960 1089.350 ;
        RECT 1688.760 1089.030 1689.020 1089.350 ;
        RECT 1688.820 64.250 1688.960 1089.030 ;
        RECT 1688.760 63.930 1689.020 64.250 ;
        RECT 2428.900 63.930 2429.160 64.250 ;
        RECT 2428.960 2.000 2429.100 63.930 ;
        RECT 2428.750 -4.000 2429.310 2.000 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1689.190 64.500 1689.510 64.560 ;
        RECT 2442.670 64.500 2442.990 64.560 ;
        RECT 1689.190 64.360 2442.990 64.500 ;
        RECT 1689.190 64.300 1689.510 64.360 ;
        RECT 2442.670 64.300 2442.990 64.360 ;
      LAYER via ;
        RECT 1689.220 64.300 1689.480 64.560 ;
        RECT 2442.700 64.300 2442.960 64.560 ;
      LAYER met2 ;
        RECT 1689.590 1100.650 1689.870 1104.000 ;
        RECT 1689.280 1100.510 1689.870 1100.650 ;
        RECT 1689.280 64.590 1689.420 1100.510 ;
        RECT 1689.590 1100.000 1689.870 1100.510 ;
        RECT 1689.220 64.270 1689.480 64.590 ;
        RECT 2442.700 64.270 2442.960 64.590 ;
        RECT 2442.760 2.450 2442.900 64.270 ;
        RECT 2442.760 2.310 2447.040 2.450 ;
        RECT 2446.900 2.000 2447.040 2.310 ;
        RECT 2446.690 -4.000 2447.250 2.000 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1696.090 64.840 1696.410 64.900 ;
        RECT 2463.370 64.840 2463.690 64.900 ;
        RECT 1696.090 64.700 2463.690 64.840 ;
        RECT 1696.090 64.640 1696.410 64.700 ;
        RECT 2463.370 64.640 2463.690 64.700 ;
      LAYER via ;
        RECT 1696.120 64.640 1696.380 64.900 ;
        RECT 2463.400 64.640 2463.660 64.900 ;
      LAYER met2 ;
        RECT 1695.570 1100.650 1695.850 1104.000 ;
        RECT 1695.570 1100.510 1696.320 1100.650 ;
        RECT 1695.570 1100.000 1695.850 1100.510 ;
        RECT 1696.180 64.930 1696.320 1100.510 ;
        RECT 1696.120 64.610 1696.380 64.930 ;
        RECT 2463.400 64.610 2463.660 64.930 ;
        RECT 2463.460 2.450 2463.600 64.610 ;
        RECT 2463.460 2.310 2464.980 2.450 ;
        RECT 2464.840 2.000 2464.980 2.310 ;
        RECT 2464.630 -4.000 2465.190 2.000 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1702.530 65.180 1702.850 65.240 ;
        RECT 2477.170 65.180 2477.490 65.240 ;
        RECT 1702.530 65.040 2477.490 65.180 ;
        RECT 1702.530 64.980 1702.850 65.040 ;
        RECT 2477.170 64.980 2477.490 65.040 ;
        RECT 2477.170 2.620 2477.490 2.680 ;
        RECT 2482.690 2.620 2483.010 2.680 ;
        RECT 2477.170 2.480 2483.010 2.620 ;
        RECT 2477.170 2.420 2477.490 2.480 ;
        RECT 2482.690 2.420 2483.010 2.480 ;
      LAYER via ;
        RECT 1702.560 64.980 1702.820 65.240 ;
        RECT 2477.200 64.980 2477.460 65.240 ;
        RECT 2477.200 2.420 2477.460 2.680 ;
        RECT 2482.720 2.420 2482.980 2.680 ;
      LAYER met2 ;
        RECT 1702.010 1100.650 1702.290 1104.000 ;
        RECT 1702.010 1100.510 1702.760 1100.650 ;
        RECT 1702.010 1100.000 1702.290 1100.510 ;
        RECT 1702.620 65.270 1702.760 1100.510 ;
        RECT 1702.560 64.950 1702.820 65.270 ;
        RECT 2477.200 64.950 2477.460 65.270 ;
        RECT 2477.260 2.710 2477.400 64.950 ;
        RECT 2477.200 2.390 2477.460 2.710 ;
        RECT 2482.720 2.390 2482.980 2.710 ;
        RECT 2482.780 2.000 2482.920 2.390 ;
        RECT 2482.570 -4.000 2483.130 2.000 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1709.965 766.105 1710.135 814.215 ;
        RECT 1709.965 703.885 1710.135 710.855 ;
        RECT 1708.585 648.805 1708.755 696.915 ;
        RECT 1709.505 517.565 1709.675 565.335 ;
        RECT 1709.965 366.265 1710.135 373.235 ;
        RECT 1709.505 68.765 1709.675 92.055 ;
      LAYER mcon ;
        RECT 1709.965 814.045 1710.135 814.215 ;
        RECT 1709.965 710.685 1710.135 710.855 ;
        RECT 1708.585 696.745 1708.755 696.915 ;
        RECT 1709.505 565.165 1709.675 565.335 ;
        RECT 1709.965 373.065 1710.135 373.235 ;
        RECT 1709.505 91.885 1709.675 92.055 ;
      LAYER met1 ;
        RECT 1708.970 1055.600 1709.290 1055.660 ;
        RECT 1709.890 1055.600 1710.210 1055.660 ;
        RECT 1708.970 1055.460 1710.210 1055.600 ;
        RECT 1708.970 1055.400 1709.290 1055.460 ;
        RECT 1709.890 1055.400 1710.210 1055.460 ;
        RECT 1709.890 814.200 1710.210 814.260 ;
        RECT 1709.695 814.060 1710.210 814.200 ;
        RECT 1709.890 814.000 1710.210 814.060 ;
        RECT 1709.890 766.260 1710.210 766.320 ;
        RECT 1709.695 766.120 1710.210 766.260 ;
        RECT 1709.890 766.060 1710.210 766.120 ;
        RECT 1709.890 710.840 1710.210 710.900 ;
        RECT 1709.695 710.700 1710.210 710.840 ;
        RECT 1709.890 710.640 1710.210 710.700 ;
        RECT 1709.890 704.040 1710.210 704.100 ;
        RECT 1709.695 703.900 1710.210 704.040 ;
        RECT 1709.890 703.840 1710.210 703.900 ;
        RECT 1708.525 696.900 1708.815 696.945 ;
        RECT 1709.890 696.900 1710.210 696.960 ;
        RECT 1708.525 696.760 1710.210 696.900 ;
        RECT 1708.525 696.715 1708.815 696.760 ;
        RECT 1709.890 696.700 1710.210 696.760 ;
        RECT 1708.510 648.960 1708.830 649.020 ;
        RECT 1708.315 648.820 1708.830 648.960 ;
        RECT 1708.510 648.760 1708.830 648.820 ;
        RECT 1708.970 566.000 1709.290 566.060 ;
        RECT 1709.430 566.000 1709.750 566.060 ;
        RECT 1708.970 565.860 1709.750 566.000 ;
        RECT 1708.970 565.800 1709.290 565.860 ;
        RECT 1709.430 565.800 1709.750 565.860 ;
        RECT 1709.430 565.320 1709.750 565.380 ;
        RECT 1709.235 565.180 1709.750 565.320 ;
        RECT 1709.430 565.120 1709.750 565.180 ;
        RECT 1709.445 517.720 1709.735 517.765 ;
        RECT 1709.890 517.720 1710.210 517.780 ;
        RECT 1709.445 517.580 1710.210 517.720 ;
        RECT 1709.445 517.535 1709.735 517.580 ;
        RECT 1709.890 517.520 1710.210 517.580 ;
        RECT 1709.890 421.640 1710.210 421.900 ;
        RECT 1709.980 421.220 1710.120 421.640 ;
        RECT 1709.890 420.960 1710.210 421.220 ;
        RECT 1709.890 373.220 1710.210 373.280 ;
        RECT 1709.695 373.080 1710.210 373.220 ;
        RECT 1709.890 373.020 1710.210 373.080 ;
        RECT 1709.890 366.420 1710.210 366.480 ;
        RECT 1709.695 366.280 1710.210 366.420 ;
        RECT 1709.890 366.220 1710.210 366.280 ;
        RECT 1709.430 324.400 1709.750 324.660 ;
        RECT 1709.520 323.920 1709.660 324.400 ;
        RECT 1709.890 323.920 1710.210 323.980 ;
        RECT 1709.520 323.780 1710.210 323.920 ;
        RECT 1709.890 323.720 1710.210 323.780 ;
        RECT 1709.890 317.460 1710.210 317.520 ;
        RECT 1709.520 317.320 1710.210 317.460 ;
        RECT 1709.520 317.180 1709.660 317.320 ;
        RECT 1709.890 317.260 1710.210 317.320 ;
        RECT 1709.430 316.920 1709.750 317.180 ;
        RECT 1709.430 227.840 1709.750 228.100 ;
        RECT 1709.520 227.420 1709.660 227.840 ;
        RECT 1709.430 227.160 1709.750 227.420 ;
        RECT 1709.430 92.040 1709.750 92.100 ;
        RECT 1709.235 91.900 1709.750 92.040 ;
        RECT 1709.430 91.840 1709.750 91.900 ;
        RECT 1709.445 68.920 1709.735 68.965 ;
        RECT 2497.870 68.920 2498.190 68.980 ;
        RECT 1709.445 68.780 2498.190 68.920 ;
        RECT 1709.445 68.735 1709.735 68.780 ;
        RECT 2497.870 68.720 2498.190 68.780 ;
      LAYER via ;
        RECT 1709.000 1055.400 1709.260 1055.660 ;
        RECT 1709.920 1055.400 1710.180 1055.660 ;
        RECT 1709.920 814.000 1710.180 814.260 ;
        RECT 1709.920 766.060 1710.180 766.320 ;
        RECT 1709.920 710.640 1710.180 710.900 ;
        RECT 1709.920 703.840 1710.180 704.100 ;
        RECT 1709.920 696.700 1710.180 696.960 ;
        RECT 1708.540 648.760 1708.800 649.020 ;
        RECT 1709.000 565.800 1709.260 566.060 ;
        RECT 1709.460 565.800 1709.720 566.060 ;
        RECT 1709.460 565.120 1709.720 565.380 ;
        RECT 1709.920 517.520 1710.180 517.780 ;
        RECT 1709.920 421.640 1710.180 421.900 ;
        RECT 1709.920 420.960 1710.180 421.220 ;
        RECT 1709.920 373.020 1710.180 373.280 ;
        RECT 1709.920 366.220 1710.180 366.480 ;
        RECT 1709.460 324.400 1709.720 324.660 ;
        RECT 1709.920 323.720 1710.180 323.980 ;
        RECT 1709.920 317.260 1710.180 317.520 ;
        RECT 1709.460 316.920 1709.720 317.180 ;
        RECT 1709.460 227.840 1709.720 228.100 ;
        RECT 1709.460 227.160 1709.720 227.420 ;
        RECT 1709.460 91.840 1709.720 92.100 ;
        RECT 2497.900 68.720 2498.160 68.980 ;
      LAYER met2 ;
        RECT 1707.990 1100.650 1708.270 1104.000 ;
        RECT 1707.990 1100.510 1709.660 1100.650 ;
        RECT 1707.990 1100.000 1708.270 1100.510 ;
        RECT 1709.520 1076.170 1709.660 1100.510 ;
        RECT 1709.520 1076.030 1710.120 1076.170 ;
        RECT 1709.980 1055.690 1710.120 1076.030 ;
        RECT 1709.000 1055.370 1709.260 1055.690 ;
        RECT 1709.920 1055.370 1710.180 1055.690 ;
        RECT 1709.060 1007.605 1709.200 1055.370 ;
        RECT 1708.990 1007.235 1709.270 1007.605 ;
        RECT 1709.910 1007.235 1710.190 1007.605 ;
        RECT 1709.980 980.290 1710.120 1007.235 ;
        RECT 1709.520 980.150 1710.120 980.290 ;
        RECT 1709.520 979.610 1709.660 980.150 ;
        RECT 1709.520 979.470 1710.120 979.610 ;
        RECT 1709.980 835.450 1710.120 979.470 ;
        RECT 1709.520 835.310 1710.120 835.450 ;
        RECT 1709.520 834.770 1709.660 835.310 ;
        RECT 1709.520 834.630 1710.120 834.770 ;
        RECT 1709.980 814.290 1710.120 834.630 ;
        RECT 1709.920 813.970 1710.180 814.290 ;
        RECT 1709.920 766.030 1710.180 766.350 ;
        RECT 1709.980 710.930 1710.120 766.030 ;
        RECT 1709.920 710.610 1710.180 710.930 ;
        RECT 1709.920 703.810 1710.180 704.130 ;
        RECT 1709.980 696.990 1710.120 703.810 ;
        RECT 1709.920 696.670 1710.180 696.990 ;
        RECT 1708.540 648.730 1708.800 649.050 ;
        RECT 1708.600 613.770 1708.740 648.730 ;
        RECT 1708.600 613.630 1709.200 613.770 ;
        RECT 1709.060 566.090 1709.200 613.630 ;
        RECT 1709.000 565.770 1709.260 566.090 ;
        RECT 1709.460 565.770 1709.720 566.090 ;
        RECT 1709.520 565.410 1709.660 565.770 ;
        RECT 1709.460 565.090 1709.720 565.410 ;
        RECT 1709.920 517.490 1710.180 517.810 ;
        RECT 1709.980 421.930 1710.120 517.490 ;
        RECT 1709.920 421.610 1710.180 421.930 ;
        RECT 1709.920 420.930 1710.180 421.250 ;
        RECT 1709.980 373.310 1710.120 420.930 ;
        RECT 1709.920 372.990 1710.180 373.310 ;
        RECT 1709.920 366.250 1710.180 366.510 ;
        RECT 1709.520 366.190 1710.180 366.250 ;
        RECT 1709.520 366.110 1710.120 366.190 ;
        RECT 1709.520 324.690 1709.660 366.110 ;
        RECT 1709.460 324.370 1709.720 324.690 ;
        RECT 1709.920 323.690 1710.180 324.010 ;
        RECT 1709.980 317.550 1710.120 323.690 ;
        RECT 1709.920 317.230 1710.180 317.550 ;
        RECT 1709.460 316.890 1709.720 317.210 ;
        RECT 1709.520 310.605 1709.660 316.890 ;
        RECT 1708.530 310.235 1708.810 310.605 ;
        RECT 1709.450 310.235 1709.730 310.605 ;
        RECT 1708.600 267.650 1708.740 310.235 ;
        RECT 1708.600 267.510 1709.660 267.650 ;
        RECT 1709.520 228.130 1709.660 267.510 ;
        RECT 1709.460 227.810 1709.720 228.130 ;
        RECT 1709.460 227.130 1709.720 227.450 ;
        RECT 1709.520 92.130 1709.660 227.130 ;
        RECT 1709.460 91.810 1709.720 92.130 ;
        RECT 2497.900 68.690 2498.160 69.010 ;
        RECT 2497.960 16.730 2498.100 68.690 ;
        RECT 2497.960 16.590 2500.860 16.730 ;
        RECT 2500.720 2.000 2500.860 16.590 ;
        RECT 2500.510 -4.000 2501.070 2.000 ;
      LAYER via2 ;
        RECT 1708.990 1007.280 1709.270 1007.560 ;
        RECT 1709.910 1007.280 1710.190 1007.560 ;
        RECT 1708.530 310.280 1708.810 310.560 ;
        RECT 1709.450 310.280 1709.730 310.560 ;
      LAYER met3 ;
        RECT 1708.965 1007.570 1709.295 1007.585 ;
        RECT 1709.885 1007.570 1710.215 1007.585 ;
        RECT 1708.965 1007.270 1710.215 1007.570 ;
        RECT 1708.965 1007.255 1709.295 1007.270 ;
        RECT 1709.885 1007.255 1710.215 1007.270 ;
        RECT 1708.505 310.570 1708.835 310.585 ;
        RECT 1709.425 310.570 1709.755 310.585 ;
        RECT 1708.505 310.270 1709.755 310.570 ;
        RECT 1708.505 310.255 1708.835 310.270 ;
        RECT 1709.425 310.255 1709.755 310.270 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1716.405 1027.905 1716.575 1055.615 ;
        RECT 1716.405 703.885 1716.575 793.475 ;
        RECT 1716.405 607.325 1716.575 655.435 ;
        RECT 1716.405 372.725 1716.575 420.835 ;
        RECT 1716.865 142.205 1717.035 186.575 ;
        RECT 1716.405 68.425 1716.575 137.955 ;
      LAYER mcon ;
        RECT 1716.405 1055.445 1716.575 1055.615 ;
        RECT 1716.405 793.305 1716.575 793.475 ;
        RECT 1716.405 655.265 1716.575 655.435 ;
        RECT 1716.405 420.665 1716.575 420.835 ;
        RECT 1716.865 186.405 1717.035 186.575 ;
        RECT 1716.405 137.785 1716.575 137.955 ;
      LAYER met1 ;
        RECT 1716.330 1055.600 1716.650 1055.660 ;
        RECT 1716.135 1055.460 1716.650 1055.600 ;
        RECT 1716.330 1055.400 1716.650 1055.460 ;
        RECT 1716.330 1028.060 1716.650 1028.120 ;
        RECT 1716.135 1027.920 1716.650 1028.060 ;
        RECT 1716.330 1027.860 1716.650 1027.920 ;
        RECT 1714.950 959.040 1715.270 959.100 ;
        RECT 1715.870 959.040 1716.190 959.100 ;
        RECT 1714.950 958.900 1716.190 959.040 ;
        RECT 1714.950 958.840 1715.270 958.900 ;
        RECT 1715.870 958.840 1716.190 958.900 ;
        RECT 1716.330 848.540 1716.650 848.600 ;
        RECT 1716.790 848.540 1717.110 848.600 ;
        RECT 1716.330 848.400 1717.110 848.540 ;
        RECT 1716.330 848.340 1716.650 848.400 ;
        RECT 1716.790 848.340 1717.110 848.400 ;
        RECT 1716.330 793.460 1716.650 793.520 ;
        RECT 1716.135 793.320 1716.650 793.460 ;
        RECT 1716.330 793.260 1716.650 793.320 ;
        RECT 1716.345 704.040 1716.635 704.085 ;
        RECT 1716.790 704.040 1717.110 704.100 ;
        RECT 1716.345 703.900 1717.110 704.040 ;
        RECT 1716.345 703.855 1716.635 703.900 ;
        RECT 1716.790 703.840 1717.110 703.900 ;
        RECT 1716.330 662.560 1716.650 662.620 ;
        RECT 1716.790 662.560 1717.110 662.620 ;
        RECT 1716.330 662.420 1717.110 662.560 ;
        RECT 1716.330 662.360 1716.650 662.420 ;
        RECT 1716.790 662.360 1717.110 662.420 ;
        RECT 1716.330 655.420 1716.650 655.480 ;
        RECT 1716.135 655.280 1716.650 655.420 ;
        RECT 1716.330 655.220 1716.650 655.280 ;
        RECT 1716.330 607.480 1716.650 607.540 ;
        RECT 1716.135 607.340 1716.650 607.480 ;
        RECT 1716.330 607.280 1716.650 607.340 ;
        RECT 1715.410 469.440 1715.730 469.500 ;
        RECT 1715.870 469.440 1716.190 469.500 ;
        RECT 1715.410 469.300 1716.190 469.440 ;
        RECT 1715.410 469.240 1715.730 469.300 ;
        RECT 1715.870 469.240 1716.190 469.300 ;
        RECT 1716.330 420.820 1716.650 420.880 ;
        RECT 1716.135 420.680 1716.650 420.820 ;
        RECT 1716.330 420.620 1716.650 420.680 ;
        RECT 1716.345 372.880 1716.635 372.925 ;
        RECT 1716.790 372.880 1717.110 372.940 ;
        RECT 1716.345 372.740 1717.110 372.880 ;
        RECT 1716.345 372.695 1716.635 372.740 ;
        RECT 1716.790 372.680 1717.110 372.740 ;
        RECT 1715.870 317.460 1716.190 317.520 ;
        RECT 1716.790 317.460 1717.110 317.520 ;
        RECT 1715.870 317.320 1717.110 317.460 ;
        RECT 1715.870 317.260 1716.190 317.320 ;
        RECT 1716.790 317.260 1717.110 317.320 ;
        RECT 1716.790 186.560 1717.110 186.620 ;
        RECT 1716.595 186.420 1717.110 186.560 ;
        RECT 1716.790 186.360 1717.110 186.420 ;
        RECT 1716.790 142.360 1717.110 142.420 ;
        RECT 1716.595 142.220 1717.110 142.360 ;
        RECT 1716.790 142.160 1717.110 142.220 ;
        RECT 1716.345 137.940 1716.635 137.985 ;
        RECT 1716.790 137.940 1717.110 138.000 ;
        RECT 1716.345 137.800 1717.110 137.940 ;
        RECT 1716.345 137.755 1716.635 137.800 ;
        RECT 1716.790 137.740 1717.110 137.800 ;
        RECT 1716.345 68.580 1716.635 68.625 ;
        RECT 2511.670 68.580 2511.990 68.640 ;
        RECT 1716.345 68.440 2511.990 68.580 ;
        RECT 1716.345 68.395 1716.635 68.440 ;
        RECT 2511.670 68.380 2511.990 68.440 ;
        RECT 2511.670 16.900 2511.990 16.960 ;
        RECT 2518.110 16.900 2518.430 16.960 ;
        RECT 2511.670 16.760 2518.430 16.900 ;
        RECT 2511.670 16.700 2511.990 16.760 ;
        RECT 2518.110 16.700 2518.430 16.760 ;
      LAYER via ;
        RECT 1716.360 1055.400 1716.620 1055.660 ;
        RECT 1716.360 1027.860 1716.620 1028.120 ;
        RECT 1714.980 958.840 1715.240 959.100 ;
        RECT 1715.900 958.840 1716.160 959.100 ;
        RECT 1716.360 848.340 1716.620 848.600 ;
        RECT 1716.820 848.340 1717.080 848.600 ;
        RECT 1716.360 793.260 1716.620 793.520 ;
        RECT 1716.820 703.840 1717.080 704.100 ;
        RECT 1716.360 662.360 1716.620 662.620 ;
        RECT 1716.820 662.360 1717.080 662.620 ;
        RECT 1716.360 655.220 1716.620 655.480 ;
        RECT 1716.360 607.280 1716.620 607.540 ;
        RECT 1715.440 469.240 1715.700 469.500 ;
        RECT 1715.900 469.240 1716.160 469.500 ;
        RECT 1716.360 420.620 1716.620 420.880 ;
        RECT 1716.820 372.680 1717.080 372.940 ;
        RECT 1715.900 317.260 1716.160 317.520 ;
        RECT 1716.820 317.260 1717.080 317.520 ;
        RECT 1716.820 186.360 1717.080 186.620 ;
        RECT 1716.820 142.160 1717.080 142.420 ;
        RECT 1716.820 137.740 1717.080 138.000 ;
        RECT 2511.700 68.380 2511.960 68.640 ;
        RECT 2511.700 16.700 2511.960 16.960 ;
        RECT 2518.140 16.700 2518.400 16.960 ;
      LAYER met2 ;
        RECT 1713.970 1100.650 1714.250 1104.000 ;
        RECT 1713.970 1100.510 1716.100 1100.650 ;
        RECT 1713.970 1100.000 1714.250 1100.510 ;
        RECT 1715.960 1076.170 1716.100 1100.510 ;
        RECT 1715.960 1076.030 1716.560 1076.170 ;
        RECT 1716.420 1055.690 1716.560 1076.030 ;
        RECT 1716.360 1055.370 1716.620 1055.690 ;
        RECT 1716.360 1027.830 1716.620 1028.150 ;
        RECT 1716.420 1007.490 1716.560 1027.830 ;
        RECT 1716.420 1007.350 1717.020 1007.490 ;
        RECT 1716.880 966.125 1717.020 1007.350 ;
        RECT 1715.890 965.755 1716.170 966.125 ;
        RECT 1716.810 965.755 1717.090 966.125 ;
        RECT 1715.960 959.130 1716.100 965.755 ;
        RECT 1714.980 958.810 1715.240 959.130 ;
        RECT 1715.900 958.810 1716.160 959.130 ;
        RECT 1715.040 911.045 1715.180 958.810 ;
        RECT 1714.970 910.675 1715.250 911.045 ;
        RECT 1715.890 910.675 1716.170 911.045 ;
        RECT 1715.960 862.765 1716.100 910.675 ;
        RECT 1715.890 862.395 1716.170 862.765 ;
        RECT 1716.810 862.395 1717.090 862.765 ;
        RECT 1716.880 848.630 1717.020 862.395 ;
        RECT 1716.360 848.310 1716.620 848.630 ;
        RECT 1716.820 848.310 1717.080 848.630 ;
        RECT 1716.420 801.565 1716.560 848.310 ;
        RECT 1716.350 801.195 1716.630 801.565 ;
        RECT 1716.350 800.515 1716.630 800.885 ;
        RECT 1716.420 793.550 1716.560 800.515 ;
        RECT 1716.360 793.230 1716.620 793.550 ;
        RECT 1716.820 703.810 1717.080 704.130 ;
        RECT 1716.880 662.650 1717.020 703.810 ;
        RECT 1716.360 662.330 1716.620 662.650 ;
        RECT 1716.820 662.330 1717.080 662.650 ;
        RECT 1716.420 655.510 1716.560 662.330 ;
        RECT 1716.360 655.190 1716.620 655.510 ;
        RECT 1716.360 607.250 1716.620 607.570 ;
        RECT 1716.420 590.650 1716.560 607.250 ;
        RECT 1715.960 590.510 1716.560 590.650 ;
        RECT 1715.960 517.210 1716.100 590.510 ;
        RECT 1715.500 517.070 1716.100 517.210 ;
        RECT 1715.500 469.530 1715.640 517.070 ;
        RECT 1715.440 469.210 1715.700 469.530 ;
        RECT 1715.900 469.210 1716.160 469.530 ;
        RECT 1715.960 434.930 1716.100 469.210 ;
        RECT 1715.960 434.790 1716.560 434.930 ;
        RECT 1716.420 420.910 1716.560 434.790 ;
        RECT 1716.360 420.590 1716.620 420.910 ;
        RECT 1716.820 372.650 1717.080 372.970 ;
        RECT 1716.880 325.565 1717.020 372.650 ;
        RECT 1716.810 325.195 1717.090 325.565 ;
        RECT 1715.890 324.515 1716.170 324.885 ;
        RECT 1715.960 317.550 1716.100 324.515 ;
        RECT 1715.900 317.230 1716.160 317.550 ;
        RECT 1716.820 317.230 1717.080 317.550 ;
        RECT 1716.880 186.650 1717.020 317.230 ;
        RECT 1716.820 186.330 1717.080 186.650 ;
        RECT 1716.820 142.130 1717.080 142.450 ;
        RECT 1716.880 138.030 1717.020 142.130 ;
        RECT 1716.820 137.710 1717.080 138.030 ;
        RECT 2511.700 68.350 2511.960 68.670 ;
        RECT 2511.760 16.990 2511.900 68.350 ;
        RECT 2511.700 16.670 2511.960 16.990 ;
        RECT 2518.140 16.670 2518.400 16.990 ;
        RECT 2518.200 2.000 2518.340 16.670 ;
        RECT 2517.990 -4.000 2518.550 2.000 ;
      LAYER via2 ;
        RECT 1715.890 965.800 1716.170 966.080 ;
        RECT 1716.810 965.800 1717.090 966.080 ;
        RECT 1714.970 910.720 1715.250 911.000 ;
        RECT 1715.890 910.720 1716.170 911.000 ;
        RECT 1715.890 862.440 1716.170 862.720 ;
        RECT 1716.810 862.440 1717.090 862.720 ;
        RECT 1716.350 801.240 1716.630 801.520 ;
        RECT 1716.350 800.560 1716.630 800.840 ;
        RECT 1716.810 325.240 1717.090 325.520 ;
        RECT 1715.890 324.560 1716.170 324.840 ;
      LAYER met3 ;
        RECT 1715.865 966.090 1716.195 966.105 ;
        RECT 1716.785 966.090 1717.115 966.105 ;
        RECT 1715.865 965.790 1717.115 966.090 ;
        RECT 1715.865 965.775 1716.195 965.790 ;
        RECT 1716.785 965.775 1717.115 965.790 ;
        RECT 1714.945 911.010 1715.275 911.025 ;
        RECT 1715.865 911.010 1716.195 911.025 ;
        RECT 1714.945 910.710 1716.195 911.010 ;
        RECT 1714.945 910.695 1715.275 910.710 ;
        RECT 1715.865 910.695 1716.195 910.710 ;
        RECT 1715.865 862.730 1716.195 862.745 ;
        RECT 1716.785 862.730 1717.115 862.745 ;
        RECT 1715.865 862.430 1717.115 862.730 ;
        RECT 1715.865 862.415 1716.195 862.430 ;
        RECT 1716.785 862.415 1717.115 862.430 ;
        RECT 1716.325 801.215 1716.655 801.545 ;
        RECT 1716.340 800.865 1716.640 801.215 ;
        RECT 1716.325 800.535 1716.655 800.865 ;
        RECT 1716.785 325.530 1717.115 325.545 ;
        RECT 1716.110 325.230 1717.115 325.530 ;
        RECT 1716.110 324.865 1716.410 325.230 ;
        RECT 1716.785 325.215 1717.115 325.230 ;
        RECT 1715.865 324.550 1716.410 324.865 ;
        RECT 1715.865 324.535 1716.195 324.550 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1722.845 1027.905 1723.015 1055.615 ;
        RECT 1722.845 814.385 1723.015 837.675 ;
        RECT 1722.385 469.285 1722.555 517.395 ;
        RECT 1722.845 338.045 1723.015 396.695 ;
        RECT 1722.385 276.165 1722.555 324.275 ;
        RECT 1722.845 205.445 1723.015 258.995 ;
        RECT 1723.305 144.925 1723.475 193.035 ;
        RECT 1722.845 68.085 1723.015 137.955 ;
      LAYER mcon ;
        RECT 1722.845 1055.445 1723.015 1055.615 ;
        RECT 1722.845 837.505 1723.015 837.675 ;
        RECT 1722.385 517.225 1722.555 517.395 ;
        RECT 1722.845 396.525 1723.015 396.695 ;
        RECT 1722.385 324.105 1722.555 324.275 ;
        RECT 1722.845 258.825 1723.015 258.995 ;
        RECT 1723.305 192.865 1723.475 193.035 ;
        RECT 1722.845 137.785 1723.015 137.955 ;
      LAYER met1 ;
        RECT 1722.770 1055.600 1723.090 1055.660 ;
        RECT 1722.575 1055.460 1723.090 1055.600 ;
        RECT 1722.770 1055.400 1723.090 1055.460 ;
        RECT 1722.770 1028.060 1723.090 1028.120 ;
        RECT 1722.575 1027.920 1723.090 1028.060 ;
        RECT 1722.770 1027.860 1723.090 1027.920 ;
        RECT 1721.850 918.240 1722.170 918.300 ;
        RECT 1722.770 918.240 1723.090 918.300 ;
        RECT 1721.850 918.100 1723.090 918.240 ;
        RECT 1721.850 918.040 1722.170 918.100 ;
        RECT 1722.770 918.040 1723.090 918.100 ;
        RECT 1722.770 883.020 1723.090 883.280 ;
        RECT 1722.310 882.880 1722.630 882.940 ;
        RECT 1722.860 882.880 1723.000 883.020 ;
        RECT 1722.310 882.740 1723.000 882.880 ;
        RECT 1722.310 882.680 1722.630 882.740 ;
        RECT 1722.785 837.660 1723.075 837.705 ;
        RECT 1723.230 837.660 1723.550 837.720 ;
        RECT 1722.785 837.520 1723.550 837.660 ;
        RECT 1722.785 837.475 1723.075 837.520 ;
        RECT 1723.230 837.460 1723.550 837.520 ;
        RECT 1722.770 814.540 1723.090 814.600 ;
        RECT 1722.575 814.400 1723.090 814.540 ;
        RECT 1722.770 814.340 1723.090 814.400 ;
        RECT 1722.310 759.120 1722.630 759.180 ;
        RECT 1722.770 759.120 1723.090 759.180 ;
        RECT 1722.310 758.980 1723.090 759.120 ;
        RECT 1722.310 758.920 1722.630 758.980 ;
        RECT 1722.770 758.920 1723.090 758.980 ;
        RECT 1721.390 704.040 1721.710 704.100 ;
        RECT 1721.850 704.040 1722.170 704.100 ;
        RECT 1721.390 703.900 1722.170 704.040 ;
        RECT 1721.390 703.840 1721.710 703.900 ;
        RECT 1721.850 703.840 1722.170 703.900 ;
        RECT 1721.390 661.880 1721.710 661.940 ;
        RECT 1722.770 661.880 1723.090 661.940 ;
        RECT 1721.390 661.740 1723.090 661.880 ;
        RECT 1721.390 661.680 1721.710 661.740 ;
        RECT 1722.770 661.680 1723.090 661.740 ;
        RECT 1722.310 613.940 1722.630 614.000 ;
        RECT 1722.770 613.940 1723.090 614.000 ;
        RECT 1722.310 613.800 1723.090 613.940 ;
        RECT 1722.310 613.740 1722.630 613.800 ;
        RECT 1722.770 613.740 1723.090 613.800 ;
        RECT 1722.325 517.380 1722.615 517.425 ;
        RECT 1722.770 517.380 1723.090 517.440 ;
        RECT 1722.325 517.240 1723.090 517.380 ;
        RECT 1722.325 517.195 1722.615 517.240 ;
        RECT 1722.770 517.180 1723.090 517.240 ;
        RECT 1722.310 469.440 1722.630 469.500 ;
        RECT 1722.115 469.300 1722.630 469.440 ;
        RECT 1722.310 469.240 1722.630 469.300 ;
        RECT 1722.770 396.680 1723.090 396.740 ;
        RECT 1722.575 396.540 1723.090 396.680 ;
        RECT 1722.770 396.480 1723.090 396.540 ;
        RECT 1722.770 338.200 1723.090 338.260 ;
        RECT 1722.575 338.060 1723.090 338.200 ;
        RECT 1722.770 338.000 1723.090 338.060 ;
        RECT 1722.325 324.260 1722.615 324.305 ;
        RECT 1722.770 324.260 1723.090 324.320 ;
        RECT 1722.325 324.120 1723.090 324.260 ;
        RECT 1722.325 324.075 1722.615 324.120 ;
        RECT 1722.770 324.060 1723.090 324.120 ;
        RECT 1722.310 276.320 1722.630 276.380 ;
        RECT 1722.115 276.180 1722.630 276.320 ;
        RECT 1722.310 276.120 1722.630 276.180 ;
        RECT 1722.310 258.980 1722.630 259.040 ;
        RECT 1722.785 258.980 1723.075 259.025 ;
        RECT 1722.310 258.840 1723.075 258.980 ;
        RECT 1722.310 258.780 1722.630 258.840 ;
        RECT 1722.785 258.795 1723.075 258.840 ;
        RECT 1722.770 205.600 1723.090 205.660 ;
        RECT 1722.575 205.460 1723.090 205.600 ;
        RECT 1722.770 205.400 1723.090 205.460 ;
        RECT 1723.230 193.020 1723.550 193.080 ;
        RECT 1723.035 192.880 1723.550 193.020 ;
        RECT 1723.230 192.820 1723.550 192.880 ;
        RECT 1723.230 145.080 1723.550 145.140 ;
        RECT 1723.035 144.940 1723.550 145.080 ;
        RECT 1723.230 144.880 1723.550 144.940 ;
        RECT 1722.785 137.940 1723.075 137.985 ;
        RECT 1723.230 137.940 1723.550 138.000 ;
        RECT 1722.785 137.800 1723.550 137.940 ;
        RECT 1722.785 137.755 1723.075 137.800 ;
        RECT 1723.230 137.740 1723.550 137.800 ;
        RECT 1722.785 68.240 1723.075 68.285 ;
        RECT 2532.370 68.240 2532.690 68.300 ;
        RECT 1722.785 68.100 2532.690 68.240 ;
        RECT 1722.785 68.055 1723.075 68.100 ;
        RECT 2532.370 68.040 2532.690 68.100 ;
      LAYER via ;
        RECT 1722.800 1055.400 1723.060 1055.660 ;
        RECT 1722.800 1027.860 1723.060 1028.120 ;
        RECT 1721.880 918.040 1722.140 918.300 ;
        RECT 1722.800 918.040 1723.060 918.300 ;
        RECT 1722.800 883.020 1723.060 883.280 ;
        RECT 1722.340 882.680 1722.600 882.940 ;
        RECT 1723.260 837.460 1723.520 837.720 ;
        RECT 1722.800 814.340 1723.060 814.600 ;
        RECT 1722.340 758.920 1722.600 759.180 ;
        RECT 1722.800 758.920 1723.060 759.180 ;
        RECT 1721.420 703.840 1721.680 704.100 ;
        RECT 1721.880 703.840 1722.140 704.100 ;
        RECT 1721.420 661.680 1721.680 661.940 ;
        RECT 1722.800 661.680 1723.060 661.940 ;
        RECT 1722.340 613.740 1722.600 614.000 ;
        RECT 1722.800 613.740 1723.060 614.000 ;
        RECT 1722.800 517.180 1723.060 517.440 ;
        RECT 1722.340 469.240 1722.600 469.500 ;
        RECT 1722.800 396.480 1723.060 396.740 ;
        RECT 1722.800 338.000 1723.060 338.260 ;
        RECT 1722.800 324.060 1723.060 324.320 ;
        RECT 1722.340 276.120 1722.600 276.380 ;
        RECT 1722.340 258.780 1722.600 259.040 ;
        RECT 1722.800 205.400 1723.060 205.660 ;
        RECT 1723.260 192.820 1723.520 193.080 ;
        RECT 1723.260 144.880 1723.520 145.140 ;
        RECT 1723.260 137.740 1723.520 138.000 ;
        RECT 2532.400 68.040 2532.660 68.300 ;
      LAYER met2 ;
        RECT 1720.410 1100.650 1720.690 1104.000 ;
        RECT 1720.410 1100.510 1721.620 1100.650 ;
        RECT 1720.410 1100.000 1720.690 1100.510 ;
        RECT 1721.480 1088.410 1721.620 1100.510 ;
        RECT 1721.480 1088.270 1722.540 1088.410 ;
        RECT 1722.400 1076.170 1722.540 1088.270 ;
        RECT 1722.400 1076.030 1723.000 1076.170 ;
        RECT 1722.860 1055.690 1723.000 1076.030 ;
        RECT 1722.800 1055.370 1723.060 1055.690 ;
        RECT 1722.800 1027.830 1723.060 1028.150 ;
        RECT 1722.860 1007.490 1723.000 1027.830 ;
        RECT 1722.860 1007.350 1723.460 1007.490 ;
        RECT 1723.320 966.125 1723.460 1007.350 ;
        RECT 1721.870 965.755 1722.150 966.125 ;
        RECT 1723.250 965.755 1723.530 966.125 ;
        RECT 1721.940 918.330 1722.080 965.755 ;
        RECT 1721.880 918.010 1722.140 918.330 ;
        RECT 1722.800 918.010 1723.060 918.330 ;
        RECT 1722.860 883.310 1723.000 918.010 ;
        RECT 1722.800 882.990 1723.060 883.310 ;
        RECT 1722.340 882.650 1722.600 882.970 ;
        RECT 1722.400 862.765 1722.540 882.650 ;
        RECT 1722.330 862.395 1722.610 862.765 ;
        RECT 1723.250 862.395 1723.530 862.765 ;
        RECT 1723.320 837.750 1723.460 862.395 ;
        RECT 1723.260 837.430 1723.520 837.750 ;
        RECT 1722.800 814.310 1723.060 814.630 ;
        RECT 1722.860 759.210 1723.000 814.310 ;
        RECT 1722.340 758.890 1722.600 759.210 ;
        RECT 1722.800 758.890 1723.060 759.210 ;
        RECT 1722.400 711.010 1722.540 758.890 ;
        RECT 1721.940 710.870 1722.540 711.010 ;
        RECT 1721.940 704.130 1722.080 710.870 ;
        RECT 1721.420 703.810 1721.680 704.130 ;
        RECT 1721.880 703.810 1722.140 704.130 ;
        RECT 1721.480 661.970 1721.620 703.810 ;
        RECT 1721.420 661.650 1721.680 661.970 ;
        RECT 1722.800 661.650 1723.060 661.970 ;
        RECT 1722.860 614.030 1723.000 661.650 ;
        RECT 1722.340 613.710 1722.600 614.030 ;
        RECT 1722.800 613.710 1723.060 614.030 ;
        RECT 1722.400 548.490 1722.540 613.710 ;
        RECT 1722.400 548.350 1723.000 548.490 ;
        RECT 1722.860 517.470 1723.000 548.350 ;
        RECT 1722.800 517.150 1723.060 517.470 ;
        RECT 1722.340 469.210 1722.600 469.530 ;
        RECT 1722.400 434.930 1722.540 469.210 ;
        RECT 1722.400 434.790 1723.000 434.930 ;
        RECT 1722.860 396.770 1723.000 434.790 ;
        RECT 1722.800 396.450 1723.060 396.770 ;
        RECT 1722.800 337.970 1723.060 338.290 ;
        RECT 1722.860 324.350 1723.000 337.970 ;
        RECT 1722.800 324.030 1723.060 324.350 ;
        RECT 1722.340 276.090 1722.600 276.410 ;
        RECT 1722.400 259.070 1722.540 276.090 ;
        RECT 1722.340 258.750 1722.600 259.070 ;
        RECT 1722.800 205.370 1723.060 205.690 ;
        RECT 1722.860 193.530 1723.000 205.370 ;
        RECT 1722.860 193.390 1723.460 193.530 ;
        RECT 1723.320 193.110 1723.460 193.390 ;
        RECT 1723.260 192.790 1723.520 193.110 ;
        RECT 1723.260 144.850 1723.520 145.170 ;
        RECT 1723.320 138.030 1723.460 144.850 ;
        RECT 1723.260 137.710 1723.520 138.030 ;
        RECT 2532.400 68.010 2532.660 68.330 ;
        RECT 2532.460 16.730 2532.600 68.010 ;
        RECT 2532.460 16.590 2536.280 16.730 ;
        RECT 2536.140 2.000 2536.280 16.590 ;
        RECT 2535.930 -4.000 2536.490 2.000 ;
      LAYER via2 ;
        RECT 1721.870 965.800 1722.150 966.080 ;
        RECT 1723.250 965.800 1723.530 966.080 ;
        RECT 1722.330 862.440 1722.610 862.720 ;
        RECT 1723.250 862.440 1723.530 862.720 ;
      LAYER met3 ;
        RECT 1721.845 966.090 1722.175 966.105 ;
        RECT 1723.225 966.090 1723.555 966.105 ;
        RECT 1721.845 965.790 1723.555 966.090 ;
        RECT 1721.845 965.775 1722.175 965.790 ;
        RECT 1723.225 965.775 1723.555 965.790 ;
        RECT 1722.305 862.730 1722.635 862.745 ;
        RECT 1723.225 862.730 1723.555 862.745 ;
        RECT 1722.305 862.430 1723.555 862.730 ;
        RECT 1722.305 862.415 1722.635 862.430 ;
        RECT 1723.225 862.415 1723.555 862.430 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1726.450 1088.580 1726.770 1088.640 ;
        RECT 1730.590 1088.580 1730.910 1088.640 ;
        RECT 1726.450 1088.440 1730.910 1088.580 ;
        RECT 1726.450 1088.380 1726.770 1088.440 ;
        RECT 1730.590 1088.380 1730.910 1088.440 ;
        RECT 1730.590 67.900 1730.910 67.960 ;
        RECT 2553.070 67.900 2553.390 67.960 ;
        RECT 1730.590 67.760 2553.390 67.900 ;
        RECT 1730.590 67.700 1730.910 67.760 ;
        RECT 2553.070 67.700 2553.390 67.760 ;
      LAYER via ;
        RECT 1726.480 1088.380 1726.740 1088.640 ;
        RECT 1730.620 1088.380 1730.880 1088.640 ;
        RECT 1730.620 67.700 1730.880 67.960 ;
        RECT 2553.100 67.700 2553.360 67.960 ;
      LAYER met2 ;
        RECT 1726.390 1100.580 1726.670 1104.000 ;
        RECT 1726.390 1100.000 1726.680 1100.580 ;
        RECT 1726.540 1088.670 1726.680 1100.000 ;
        RECT 1726.480 1088.350 1726.740 1088.670 ;
        RECT 1730.620 1088.350 1730.880 1088.670 ;
        RECT 1730.680 67.990 1730.820 1088.350 ;
        RECT 1730.620 67.670 1730.880 67.990 ;
        RECT 2553.100 67.670 2553.360 67.990 ;
        RECT 2553.160 17.410 2553.300 67.670 ;
        RECT 2553.160 17.270 2554.220 17.410 ;
        RECT 2554.080 2.000 2554.220 17.270 ;
        RECT 2553.870 -4.000 2554.430 2.000 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1732.430 1089.260 1732.750 1089.320 ;
        RECT 1737.490 1089.260 1737.810 1089.320 ;
        RECT 1732.430 1089.120 1737.810 1089.260 ;
        RECT 1732.430 1089.060 1732.750 1089.120 ;
        RECT 1737.490 1089.060 1737.810 1089.120 ;
        RECT 1737.490 51.580 1737.810 51.640 ;
        RECT 2566.870 51.580 2567.190 51.640 ;
        RECT 1737.490 51.440 2567.190 51.580 ;
        RECT 1737.490 51.380 1737.810 51.440 ;
        RECT 2566.870 51.380 2567.190 51.440 ;
      LAYER via ;
        RECT 1732.460 1089.060 1732.720 1089.320 ;
        RECT 1737.520 1089.060 1737.780 1089.320 ;
        RECT 1737.520 51.380 1737.780 51.640 ;
        RECT 2566.900 51.380 2567.160 51.640 ;
      LAYER met2 ;
        RECT 1732.370 1100.580 1732.650 1104.000 ;
        RECT 1732.370 1100.000 1732.660 1100.580 ;
        RECT 1732.520 1089.350 1732.660 1100.000 ;
        RECT 1732.460 1089.030 1732.720 1089.350 ;
        RECT 1737.520 1089.030 1737.780 1089.350 ;
        RECT 1737.580 51.670 1737.720 1089.030 ;
        RECT 1737.520 51.350 1737.780 51.670 ;
        RECT 2566.900 51.350 2567.160 51.670 ;
        RECT 2566.960 17.410 2567.100 51.350 ;
        RECT 2566.960 17.270 2572.160 17.410 ;
        RECT 2572.020 2.000 2572.160 17.270 ;
        RECT 2571.810 -4.000 2572.370 2.000 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1737.030 1088.580 1737.350 1088.640 ;
        RECT 1738.410 1088.580 1738.730 1088.640 ;
        RECT 1737.030 1088.440 1738.730 1088.580 ;
        RECT 1737.030 1088.380 1737.350 1088.440 ;
        RECT 1738.410 1088.380 1738.730 1088.440 ;
        RECT 1737.030 67.560 1737.350 67.620 ;
        RECT 2587.570 67.560 2587.890 67.620 ;
        RECT 1737.030 67.420 2587.890 67.560 ;
        RECT 1737.030 67.360 1737.350 67.420 ;
        RECT 2587.570 67.360 2587.890 67.420 ;
      LAYER via ;
        RECT 1737.060 1088.380 1737.320 1088.640 ;
        RECT 1738.440 1088.380 1738.700 1088.640 ;
        RECT 1737.060 67.360 1737.320 67.620 ;
        RECT 2587.600 67.360 2587.860 67.620 ;
      LAYER met2 ;
        RECT 1738.350 1100.580 1738.630 1104.000 ;
        RECT 1738.350 1100.000 1738.640 1100.580 ;
        RECT 1738.500 1088.670 1738.640 1100.000 ;
        RECT 1737.060 1088.350 1737.320 1088.670 ;
        RECT 1738.440 1088.350 1738.700 1088.670 ;
        RECT 1737.120 67.650 1737.260 1088.350 ;
        RECT 1737.060 67.330 1737.320 67.650 ;
        RECT 2587.600 67.330 2587.860 67.650 ;
        RECT 2587.660 17.410 2587.800 67.330 ;
        RECT 2587.660 17.270 2589.640 17.410 ;
        RECT 2589.500 2.000 2589.640 17.270 ;
        RECT 2589.290 -4.000 2589.850 2.000 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 823.470 28.120 823.790 28.180 ;
        RECT 1132.130 28.120 1132.450 28.180 ;
        RECT 823.470 27.980 1132.450 28.120 ;
        RECT 823.470 27.920 823.790 27.980 ;
        RECT 1132.130 27.920 1132.450 27.980 ;
      LAYER via ;
        RECT 823.500 27.920 823.760 28.180 ;
        RECT 1132.160 27.920 1132.420 28.180 ;
      LAYER met2 ;
        RECT 1132.530 1100.650 1132.810 1104.000 ;
        RECT 1132.220 1100.510 1132.810 1100.650 ;
        RECT 1132.220 28.210 1132.360 1100.510 ;
        RECT 1132.530 1100.000 1132.810 1100.510 ;
        RECT 823.500 27.890 823.760 28.210 ;
        RECT 1132.160 27.890 1132.420 28.210 ;
        RECT 823.560 2.000 823.700 27.890 ;
        RECT 823.350 -4.000 823.910 2.000 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1744.390 67.220 1744.710 67.280 ;
        RECT 2601.370 67.220 2601.690 67.280 ;
        RECT 1744.390 67.080 2601.690 67.220 ;
        RECT 1744.390 67.020 1744.710 67.080 ;
        RECT 2601.370 67.020 2601.690 67.080 ;
        RECT 2601.370 18.940 2601.690 19.000 ;
        RECT 2607.350 18.940 2607.670 19.000 ;
        RECT 2601.370 18.800 2607.670 18.940 ;
        RECT 2601.370 18.740 2601.690 18.800 ;
        RECT 2607.350 18.740 2607.670 18.800 ;
      LAYER via ;
        RECT 1744.420 67.020 1744.680 67.280 ;
        RECT 2601.400 67.020 2601.660 67.280 ;
        RECT 2601.400 18.740 2601.660 19.000 ;
        RECT 2607.380 18.740 2607.640 19.000 ;
      LAYER met2 ;
        RECT 1744.790 1100.650 1745.070 1104.000 ;
        RECT 1744.480 1100.510 1745.070 1100.650 ;
        RECT 1744.480 67.310 1744.620 1100.510 ;
        RECT 1744.790 1100.000 1745.070 1100.510 ;
        RECT 1744.420 66.990 1744.680 67.310 ;
        RECT 2601.400 66.990 2601.660 67.310 ;
        RECT 2601.460 19.030 2601.600 66.990 ;
        RECT 2601.400 18.710 2601.660 19.030 ;
        RECT 2607.380 18.710 2607.640 19.030 ;
        RECT 2607.440 2.000 2607.580 18.710 ;
        RECT 2607.230 -4.000 2607.790 2.000 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1751.290 66.880 1751.610 66.940 ;
        RECT 2622.070 66.880 2622.390 66.940 ;
        RECT 1751.290 66.740 2622.390 66.880 ;
        RECT 1751.290 66.680 1751.610 66.740 ;
        RECT 2622.070 66.680 2622.390 66.740 ;
      LAYER via ;
        RECT 1751.320 66.680 1751.580 66.940 ;
        RECT 2622.100 66.680 2622.360 66.940 ;
      LAYER met2 ;
        RECT 1750.770 1100.650 1751.050 1104.000 ;
        RECT 1750.770 1100.510 1751.520 1100.650 ;
        RECT 1750.770 1100.000 1751.050 1100.510 ;
        RECT 1751.380 66.970 1751.520 1100.510 ;
        RECT 1751.320 66.650 1751.580 66.970 ;
        RECT 2622.100 66.650 2622.360 66.970 ;
        RECT 2622.160 2.450 2622.300 66.650 ;
        RECT 2622.160 2.310 2625.520 2.450 ;
        RECT 2625.380 2.000 2625.520 2.310 ;
        RECT 2625.170 -4.000 2625.730 2.000 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1757.730 66.540 1758.050 66.600 ;
        RECT 2642.770 66.540 2643.090 66.600 ;
        RECT 1757.730 66.400 2643.090 66.540 ;
        RECT 1757.730 66.340 1758.050 66.400 ;
        RECT 2642.770 66.340 2643.090 66.400 ;
      LAYER via ;
        RECT 1757.760 66.340 1758.020 66.600 ;
        RECT 2642.800 66.340 2643.060 66.600 ;
      LAYER met2 ;
        RECT 1756.750 1100.650 1757.030 1104.000 ;
        RECT 1756.750 1100.510 1757.960 1100.650 ;
        RECT 1756.750 1100.000 1757.030 1100.510 ;
        RECT 1757.820 66.630 1757.960 1100.510 ;
        RECT 1757.760 66.310 1758.020 66.630 ;
        RECT 2642.800 66.310 2643.060 66.630 ;
        RECT 2642.860 2.450 2643.000 66.310 ;
        RECT 2642.860 2.310 2643.460 2.450 ;
        RECT 2643.320 2.000 2643.460 2.310 ;
        RECT 2643.110 -4.000 2643.670 2.000 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1764.705 58.565 1764.875 96.475 ;
      LAYER mcon ;
        RECT 1764.705 96.305 1764.875 96.475 ;
      LAYER met1 ;
        RECT 1764.170 1014.460 1764.490 1014.520 ;
        RECT 1765.090 1014.460 1765.410 1014.520 ;
        RECT 1764.170 1014.320 1765.410 1014.460 ;
        RECT 1764.170 1014.260 1764.490 1014.320 ;
        RECT 1765.090 1014.260 1765.410 1014.320 ;
        RECT 1764.630 96.460 1764.950 96.520 ;
        RECT 1764.435 96.320 1764.950 96.460 ;
        RECT 1764.630 96.260 1764.950 96.320 ;
        RECT 1764.645 58.720 1764.935 58.765 ;
        RECT 2656.570 58.720 2656.890 58.780 ;
        RECT 1764.645 58.580 2656.890 58.720 ;
        RECT 1764.645 58.535 1764.935 58.580 ;
        RECT 2656.570 58.520 2656.890 58.580 ;
      LAYER via ;
        RECT 1764.200 1014.260 1764.460 1014.520 ;
        RECT 1765.120 1014.260 1765.380 1014.520 ;
        RECT 1764.660 96.260 1764.920 96.520 ;
        RECT 2656.600 58.520 2656.860 58.780 ;
      LAYER met2 ;
        RECT 1763.190 1100.650 1763.470 1104.000 ;
        RECT 1763.190 1100.510 1764.860 1100.650 ;
        RECT 1763.190 1100.000 1763.470 1100.510 ;
        RECT 1764.720 1076.170 1764.860 1100.510 ;
        RECT 1764.720 1076.030 1765.320 1076.170 ;
        RECT 1765.180 1062.685 1765.320 1076.030 ;
        RECT 1764.190 1062.315 1764.470 1062.685 ;
        RECT 1765.110 1062.315 1765.390 1062.685 ;
        RECT 1764.260 1014.550 1764.400 1062.315 ;
        RECT 1764.200 1014.230 1764.460 1014.550 ;
        RECT 1765.120 1014.230 1765.380 1014.550 ;
        RECT 1765.180 980.290 1765.320 1014.230 ;
        RECT 1764.720 980.150 1765.320 980.290 ;
        RECT 1764.720 979.610 1764.860 980.150 ;
        RECT 1764.720 979.470 1765.320 979.610 ;
        RECT 1765.180 835.450 1765.320 979.470 ;
        RECT 1764.720 835.310 1765.320 835.450 ;
        RECT 1764.720 834.770 1764.860 835.310 ;
        RECT 1764.720 834.630 1765.320 834.770 ;
        RECT 1765.180 738.890 1765.320 834.630 ;
        RECT 1764.720 738.750 1765.320 738.890 ;
        RECT 1764.720 738.210 1764.860 738.750 ;
        RECT 1764.720 738.070 1765.320 738.210 ;
        RECT 1765.180 642.330 1765.320 738.070 ;
        RECT 1764.720 642.190 1765.320 642.330 ;
        RECT 1764.720 641.650 1764.860 642.190 ;
        RECT 1764.720 641.510 1765.320 641.650 ;
        RECT 1765.180 545.770 1765.320 641.510 ;
        RECT 1764.720 545.630 1765.320 545.770 ;
        RECT 1764.720 545.090 1764.860 545.630 ;
        RECT 1764.720 544.950 1765.320 545.090 ;
        RECT 1765.180 449.210 1765.320 544.950 ;
        RECT 1764.720 449.070 1765.320 449.210 ;
        RECT 1764.720 448.530 1764.860 449.070 ;
        RECT 1764.720 448.390 1765.320 448.530 ;
        RECT 1765.180 351.970 1765.320 448.390 ;
        RECT 1764.720 351.830 1765.320 351.970 ;
        RECT 1764.720 351.290 1764.860 351.830 ;
        RECT 1764.720 351.150 1765.320 351.290 ;
        RECT 1765.180 255.410 1765.320 351.150 ;
        RECT 1764.720 255.270 1765.320 255.410 ;
        RECT 1764.720 254.730 1764.860 255.270 ;
        RECT 1764.720 254.590 1765.320 254.730 ;
        RECT 1765.180 158.850 1765.320 254.590 ;
        RECT 1764.720 158.710 1765.320 158.850 ;
        RECT 1764.720 96.550 1764.860 158.710 ;
        RECT 1764.660 96.230 1764.920 96.550 ;
        RECT 2656.600 58.490 2656.860 58.810 ;
        RECT 2656.660 2.450 2656.800 58.490 ;
        RECT 2656.660 2.310 2661.400 2.450 ;
        RECT 2661.260 2.000 2661.400 2.310 ;
        RECT 2661.050 -4.000 2661.610 2.000 ;
      LAYER via2 ;
        RECT 1764.190 1062.360 1764.470 1062.640 ;
        RECT 1765.110 1062.360 1765.390 1062.640 ;
      LAYER met3 ;
        RECT 1764.165 1062.650 1764.495 1062.665 ;
        RECT 1765.085 1062.650 1765.415 1062.665 ;
        RECT 1764.165 1062.350 1765.415 1062.650 ;
        RECT 1764.165 1062.335 1764.495 1062.350 ;
        RECT 1765.085 1062.335 1765.415 1062.350 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1771.145 917.405 1771.315 959.055 ;
        RECT 1771.605 882.725 1771.775 910.775 ;
        RECT 1771.605 786.505 1771.775 814.215 ;
        RECT 1772.065 620.925 1772.235 641.835 ;
        RECT 1771.145 565.845 1771.315 573.155 ;
        RECT 1772.065 483.225 1772.235 548.675 ;
        RECT 1771.605 241.825 1771.775 289.595 ;
        RECT 1771.605 205.445 1771.775 241.315 ;
        RECT 1771.605 89.845 1771.775 137.955 ;
      LAYER mcon ;
        RECT 1771.145 958.885 1771.315 959.055 ;
        RECT 1771.605 910.605 1771.775 910.775 ;
        RECT 1771.605 814.045 1771.775 814.215 ;
        RECT 1772.065 641.665 1772.235 641.835 ;
        RECT 1771.145 572.985 1771.315 573.155 ;
        RECT 1772.065 548.505 1772.235 548.675 ;
        RECT 1771.605 289.425 1771.775 289.595 ;
        RECT 1771.605 241.145 1771.775 241.315 ;
        RECT 1771.605 137.785 1771.775 137.955 ;
      LAYER met1 ;
        RECT 1770.610 1055.600 1770.930 1055.660 ;
        RECT 1771.070 1055.600 1771.390 1055.660 ;
        RECT 1770.610 1055.460 1771.390 1055.600 ;
        RECT 1770.610 1055.400 1770.930 1055.460 ;
        RECT 1771.070 1055.400 1771.390 1055.460 ;
        RECT 1771.070 959.040 1771.390 959.100 ;
        RECT 1770.875 958.900 1771.390 959.040 ;
        RECT 1771.070 958.840 1771.390 958.900 ;
        RECT 1771.070 917.560 1771.390 917.620 ;
        RECT 1770.875 917.420 1771.390 917.560 ;
        RECT 1771.070 917.360 1771.390 917.420 ;
        RECT 1771.530 910.760 1771.850 910.820 ;
        RECT 1771.335 910.620 1771.850 910.760 ;
        RECT 1771.530 910.560 1771.850 910.620 ;
        RECT 1771.545 882.880 1771.835 882.925 ;
        RECT 1771.990 882.880 1772.310 882.940 ;
        RECT 1771.545 882.740 1772.310 882.880 ;
        RECT 1771.545 882.695 1771.835 882.740 ;
        RECT 1771.990 882.680 1772.310 882.740 ;
        RECT 1771.530 821.340 1771.850 821.400 ;
        RECT 1771.990 821.340 1772.310 821.400 ;
        RECT 1771.530 821.200 1772.310 821.340 ;
        RECT 1771.530 821.140 1771.850 821.200 ;
        RECT 1771.990 821.140 1772.310 821.200 ;
        RECT 1771.530 814.200 1771.850 814.260 ;
        RECT 1771.335 814.060 1771.850 814.200 ;
        RECT 1771.530 814.000 1771.850 814.060 ;
        RECT 1771.530 786.660 1771.850 786.720 ;
        RECT 1771.335 786.520 1771.850 786.660 ;
        RECT 1771.530 786.460 1771.850 786.520 ;
        RECT 1771.990 738.860 1772.310 739.120 ;
        RECT 1772.080 738.440 1772.220 738.860 ;
        RECT 1771.990 738.180 1772.310 738.440 ;
        RECT 1771.990 641.820 1772.310 641.880 ;
        RECT 1771.795 641.680 1772.310 641.820 ;
        RECT 1771.990 641.620 1772.310 641.680 ;
        RECT 1771.990 621.080 1772.310 621.140 ;
        RECT 1771.795 620.940 1772.310 621.080 ;
        RECT 1771.990 620.880 1772.310 620.940 ;
        RECT 1771.085 573.140 1771.375 573.185 ;
        RECT 1771.990 573.140 1772.310 573.200 ;
        RECT 1771.085 573.000 1772.310 573.140 ;
        RECT 1771.085 572.955 1771.375 573.000 ;
        RECT 1771.990 572.940 1772.310 573.000 ;
        RECT 1771.070 566.000 1771.390 566.060 ;
        RECT 1770.875 565.860 1771.390 566.000 ;
        RECT 1771.070 565.800 1771.390 565.860 ;
        RECT 1771.070 548.660 1771.390 548.720 ;
        RECT 1772.005 548.660 1772.295 548.705 ;
        RECT 1771.070 548.520 1772.295 548.660 ;
        RECT 1771.070 548.460 1771.390 548.520 ;
        RECT 1772.005 548.475 1772.295 548.520 ;
        RECT 1771.990 483.380 1772.310 483.440 ;
        RECT 1771.795 483.240 1772.310 483.380 ;
        RECT 1771.990 483.180 1772.310 483.240 ;
        RECT 1771.990 290.740 1772.310 291.000 ;
        RECT 1772.080 290.320 1772.220 290.740 ;
        RECT 1771.990 290.060 1772.310 290.320 ;
        RECT 1771.545 289.580 1771.835 289.625 ;
        RECT 1771.990 289.580 1772.310 289.640 ;
        RECT 1771.545 289.440 1772.310 289.580 ;
        RECT 1771.545 289.395 1771.835 289.440 ;
        RECT 1771.990 289.380 1772.310 289.440 ;
        RECT 1771.530 241.980 1771.850 242.040 ;
        RECT 1771.335 241.840 1771.850 241.980 ;
        RECT 1771.530 241.780 1771.850 241.840 ;
        RECT 1771.530 241.300 1771.850 241.360 ;
        RECT 1771.335 241.160 1771.850 241.300 ;
        RECT 1771.530 241.100 1771.850 241.160 ;
        RECT 1771.530 205.600 1771.850 205.660 ;
        RECT 1771.335 205.460 1771.850 205.600 ;
        RECT 1771.530 205.400 1771.850 205.460 ;
        RECT 1771.545 137.940 1771.835 137.985 ;
        RECT 1771.990 137.940 1772.310 138.000 ;
        RECT 1771.545 137.800 1772.310 137.940 ;
        RECT 1771.545 137.755 1771.835 137.800 ;
        RECT 1771.990 137.740 1772.310 137.800 ;
        RECT 1771.530 90.000 1771.850 90.060 ;
        RECT 1771.335 89.860 1771.850 90.000 ;
        RECT 1771.530 89.800 1771.850 89.860 ;
        RECT 1771.530 66.200 1771.850 66.260 ;
        RECT 2677.270 66.200 2677.590 66.260 ;
        RECT 1771.530 66.060 2677.590 66.200 ;
        RECT 1771.530 66.000 1771.850 66.060 ;
        RECT 2677.270 66.000 2677.590 66.060 ;
      LAYER via ;
        RECT 1770.640 1055.400 1770.900 1055.660 ;
        RECT 1771.100 1055.400 1771.360 1055.660 ;
        RECT 1771.100 958.840 1771.360 959.100 ;
        RECT 1771.100 917.360 1771.360 917.620 ;
        RECT 1771.560 910.560 1771.820 910.820 ;
        RECT 1772.020 882.680 1772.280 882.940 ;
        RECT 1771.560 821.140 1771.820 821.400 ;
        RECT 1772.020 821.140 1772.280 821.400 ;
        RECT 1771.560 814.000 1771.820 814.260 ;
        RECT 1771.560 786.460 1771.820 786.720 ;
        RECT 1772.020 738.860 1772.280 739.120 ;
        RECT 1772.020 738.180 1772.280 738.440 ;
        RECT 1772.020 641.620 1772.280 641.880 ;
        RECT 1772.020 620.880 1772.280 621.140 ;
        RECT 1772.020 572.940 1772.280 573.200 ;
        RECT 1771.100 565.800 1771.360 566.060 ;
        RECT 1771.100 548.460 1771.360 548.720 ;
        RECT 1772.020 483.180 1772.280 483.440 ;
        RECT 1772.020 290.740 1772.280 291.000 ;
        RECT 1772.020 290.060 1772.280 290.320 ;
        RECT 1772.020 289.380 1772.280 289.640 ;
        RECT 1771.560 241.780 1771.820 242.040 ;
        RECT 1771.560 241.100 1771.820 241.360 ;
        RECT 1771.560 205.400 1771.820 205.660 ;
        RECT 1772.020 137.740 1772.280 138.000 ;
        RECT 1771.560 89.800 1771.820 90.060 ;
        RECT 1771.560 66.000 1771.820 66.260 ;
        RECT 2677.300 66.000 2677.560 66.260 ;
      LAYER met2 ;
        RECT 1769.170 1100.650 1769.450 1104.000 ;
        RECT 1769.170 1100.510 1770.380 1100.650 ;
        RECT 1769.170 1100.000 1769.450 1100.510 ;
        RECT 1770.240 1088.580 1770.380 1100.510 ;
        RECT 1770.240 1088.440 1771.300 1088.580 ;
        RECT 1771.160 1076.170 1771.300 1088.440 ;
        RECT 1771.160 1076.030 1771.760 1076.170 ;
        RECT 1771.620 1062.570 1771.760 1076.030 ;
        RECT 1771.160 1062.430 1771.760 1062.570 ;
        RECT 1771.160 1055.690 1771.300 1062.430 ;
        RECT 1770.640 1055.370 1770.900 1055.690 ;
        RECT 1771.100 1055.370 1771.360 1055.690 ;
        RECT 1770.700 1007.605 1770.840 1055.370 ;
        RECT 1770.630 1007.235 1770.910 1007.605 ;
        RECT 1772.010 1007.235 1772.290 1007.605 ;
        RECT 1772.080 966.125 1772.220 1007.235 ;
        RECT 1771.090 965.755 1771.370 966.125 ;
        RECT 1772.010 965.755 1772.290 966.125 ;
        RECT 1771.160 959.130 1771.300 965.755 ;
        RECT 1771.100 958.810 1771.360 959.130 ;
        RECT 1771.100 917.330 1771.360 917.650 ;
        RECT 1771.160 910.930 1771.300 917.330 ;
        RECT 1771.160 910.850 1771.760 910.930 ;
        RECT 1771.160 910.790 1771.820 910.850 ;
        RECT 1771.560 910.530 1771.820 910.790 ;
        RECT 1772.020 882.650 1772.280 882.970 ;
        RECT 1772.080 821.430 1772.220 882.650 ;
        RECT 1771.560 821.110 1771.820 821.430 ;
        RECT 1772.020 821.110 1772.280 821.430 ;
        RECT 1771.620 814.290 1771.760 821.110 ;
        RECT 1771.560 813.970 1771.820 814.290 ;
        RECT 1771.560 786.430 1771.820 786.750 ;
        RECT 1771.620 766.090 1771.760 786.430 ;
        RECT 1771.620 765.950 1772.220 766.090 ;
        RECT 1772.080 739.150 1772.220 765.950 ;
        RECT 1772.020 738.830 1772.280 739.150 ;
        RECT 1772.020 738.150 1772.280 738.470 ;
        RECT 1772.080 641.910 1772.220 738.150 ;
        RECT 1772.020 641.590 1772.280 641.910 ;
        RECT 1772.020 620.850 1772.280 621.170 ;
        RECT 1772.080 573.230 1772.220 620.850 ;
        RECT 1772.020 572.910 1772.280 573.230 ;
        RECT 1771.100 565.770 1771.360 566.090 ;
        RECT 1771.160 548.750 1771.300 565.770 ;
        RECT 1771.100 548.430 1771.360 548.750 ;
        RECT 1772.020 483.150 1772.280 483.470 ;
        RECT 1772.080 291.030 1772.220 483.150 ;
        RECT 1772.020 290.710 1772.280 291.030 ;
        RECT 1772.020 290.030 1772.280 290.350 ;
        RECT 1772.080 289.670 1772.220 290.030 ;
        RECT 1772.020 289.350 1772.280 289.670 ;
        RECT 1771.560 241.750 1771.820 242.070 ;
        RECT 1771.620 241.390 1771.760 241.750 ;
        RECT 1771.560 241.070 1771.820 241.390 ;
        RECT 1771.560 205.370 1771.820 205.690 ;
        RECT 1771.620 193.530 1771.760 205.370 ;
        RECT 1771.620 193.390 1772.220 193.530 ;
        RECT 1772.080 138.030 1772.220 193.390 ;
        RECT 1772.020 137.710 1772.280 138.030 ;
        RECT 1771.560 89.770 1771.820 90.090 ;
        RECT 1771.620 66.290 1771.760 89.770 ;
        RECT 1771.560 65.970 1771.820 66.290 ;
        RECT 2677.300 65.970 2677.560 66.290 ;
        RECT 2677.360 2.450 2677.500 65.970 ;
        RECT 2677.360 2.310 2678.880 2.450 ;
        RECT 2678.740 2.000 2678.880 2.310 ;
        RECT 2678.530 -4.000 2679.090 2.000 ;
      LAYER via2 ;
        RECT 1770.630 1007.280 1770.910 1007.560 ;
        RECT 1772.010 1007.280 1772.290 1007.560 ;
        RECT 1771.090 965.800 1771.370 966.080 ;
        RECT 1772.010 965.800 1772.290 966.080 ;
      LAYER met3 ;
        RECT 1770.605 1007.570 1770.935 1007.585 ;
        RECT 1771.985 1007.570 1772.315 1007.585 ;
        RECT 1770.605 1007.270 1772.315 1007.570 ;
        RECT 1770.605 1007.255 1770.935 1007.270 ;
        RECT 1771.985 1007.255 1772.315 1007.270 ;
        RECT 1771.065 966.090 1771.395 966.105 ;
        RECT 1771.985 966.090 1772.315 966.105 ;
        RECT 1771.065 965.790 1772.315 966.090 ;
        RECT 1771.065 965.775 1771.395 965.790 ;
        RECT 1771.985 965.775 1772.315 965.790 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1778.045 883.065 1778.215 910.775 ;
        RECT 1778.045 821.185 1778.215 835.295 ;
        RECT 1777.585 766.105 1777.755 814.215 ;
        RECT 1778.505 620.925 1778.675 641.835 ;
        RECT 1778.045 517.565 1778.215 565.675 ;
        RECT 1778.505 421.005 1778.675 469.115 ;
        RECT 1778.045 241.485 1778.215 324.275 ;
        RECT 1777.585 89.845 1777.755 137.955 ;
      LAYER mcon ;
        RECT 1778.045 910.605 1778.215 910.775 ;
        RECT 1778.045 835.125 1778.215 835.295 ;
        RECT 1777.585 814.045 1777.755 814.215 ;
        RECT 1778.505 641.665 1778.675 641.835 ;
        RECT 1778.045 565.505 1778.215 565.675 ;
        RECT 1778.505 468.945 1778.675 469.115 ;
        RECT 1778.045 324.105 1778.215 324.275 ;
        RECT 1777.585 137.785 1777.755 137.955 ;
      LAYER met1 ;
        RECT 1775.210 1089.260 1775.530 1089.320 ;
        RECT 1777.970 1089.260 1778.290 1089.320 ;
        RECT 1775.210 1089.120 1778.290 1089.260 ;
        RECT 1775.210 1089.060 1775.530 1089.120 ;
        RECT 1777.970 1089.060 1778.290 1089.120 ;
        RECT 1777.050 1055.600 1777.370 1055.660 ;
        RECT 1777.970 1055.600 1778.290 1055.660 ;
        RECT 1777.050 1055.460 1778.290 1055.600 ;
        RECT 1777.050 1055.400 1777.370 1055.460 ;
        RECT 1777.970 1055.400 1778.290 1055.460 ;
        RECT 1777.050 959.040 1777.370 959.100 ;
        RECT 1777.510 959.040 1777.830 959.100 ;
        RECT 1777.050 958.900 1777.830 959.040 ;
        RECT 1777.050 958.840 1777.370 958.900 ;
        RECT 1777.510 958.840 1777.830 958.900 ;
        RECT 1777.970 910.760 1778.290 910.820 ;
        RECT 1777.775 910.620 1778.290 910.760 ;
        RECT 1777.970 910.560 1778.290 910.620 ;
        RECT 1777.970 883.220 1778.290 883.280 ;
        RECT 1777.775 883.080 1778.290 883.220 ;
        RECT 1777.970 883.020 1778.290 883.080 ;
        RECT 1777.985 835.280 1778.275 835.325 ;
        RECT 1778.430 835.280 1778.750 835.340 ;
        RECT 1777.985 835.140 1778.750 835.280 ;
        RECT 1777.985 835.095 1778.275 835.140 ;
        RECT 1778.430 835.080 1778.750 835.140 ;
        RECT 1777.970 821.340 1778.290 821.400 ;
        RECT 1777.775 821.200 1778.290 821.340 ;
        RECT 1777.970 821.140 1778.290 821.200 ;
        RECT 1777.525 814.200 1777.815 814.245 ;
        RECT 1777.970 814.200 1778.290 814.260 ;
        RECT 1777.525 814.060 1778.290 814.200 ;
        RECT 1777.525 814.015 1777.815 814.060 ;
        RECT 1777.970 814.000 1778.290 814.060 ;
        RECT 1777.510 766.260 1777.830 766.320 ;
        RECT 1777.315 766.120 1777.830 766.260 ;
        RECT 1777.510 766.060 1777.830 766.120 ;
        RECT 1778.430 641.820 1778.750 641.880 ;
        RECT 1778.235 641.680 1778.750 641.820 ;
        RECT 1778.430 641.620 1778.750 641.680 ;
        RECT 1778.430 621.080 1778.750 621.140 ;
        RECT 1778.235 620.940 1778.750 621.080 ;
        RECT 1778.430 620.880 1778.750 620.940 ;
        RECT 1777.970 565.660 1778.290 565.720 ;
        RECT 1777.775 565.520 1778.290 565.660 ;
        RECT 1777.970 565.460 1778.290 565.520 ;
        RECT 1777.985 517.720 1778.275 517.765 ;
        RECT 1778.430 517.720 1778.750 517.780 ;
        RECT 1777.985 517.580 1778.750 517.720 ;
        RECT 1777.985 517.535 1778.275 517.580 ;
        RECT 1778.430 517.520 1778.750 517.580 ;
        RECT 1778.430 469.100 1778.750 469.160 ;
        RECT 1778.235 468.960 1778.750 469.100 ;
        RECT 1778.430 468.900 1778.750 468.960 ;
        RECT 1778.430 421.160 1778.750 421.220 ;
        RECT 1778.235 421.020 1778.750 421.160 ;
        RECT 1778.430 420.960 1778.750 421.020 ;
        RECT 1777.985 324.260 1778.275 324.305 ;
        RECT 1778.430 324.260 1778.750 324.320 ;
        RECT 1777.985 324.120 1778.750 324.260 ;
        RECT 1777.985 324.075 1778.275 324.120 ;
        RECT 1778.430 324.060 1778.750 324.120 ;
        RECT 1777.970 241.640 1778.290 241.700 ;
        RECT 1777.775 241.500 1778.290 241.640 ;
        RECT 1777.970 241.440 1778.290 241.500 ;
        RECT 1777.525 137.940 1777.815 137.985 ;
        RECT 1778.430 137.940 1778.750 138.000 ;
        RECT 1777.525 137.800 1778.750 137.940 ;
        RECT 1777.525 137.755 1777.815 137.800 ;
        RECT 1778.430 137.740 1778.750 137.800 ;
        RECT 1777.510 90.000 1777.830 90.060 ;
        RECT 1777.315 89.860 1777.830 90.000 ;
        RECT 1777.510 89.800 1777.830 89.860 ;
        RECT 1777.510 65.860 1777.830 65.920 ;
        RECT 2691.070 65.860 2691.390 65.920 ;
        RECT 1777.510 65.720 2691.390 65.860 ;
        RECT 1777.510 65.660 1777.830 65.720 ;
        RECT 2691.070 65.660 2691.390 65.720 ;
        RECT 2691.070 2.620 2691.390 2.680 ;
        RECT 2696.590 2.620 2696.910 2.680 ;
        RECT 2691.070 2.480 2696.910 2.620 ;
        RECT 2691.070 2.420 2691.390 2.480 ;
        RECT 2696.590 2.420 2696.910 2.480 ;
      LAYER via ;
        RECT 1775.240 1089.060 1775.500 1089.320 ;
        RECT 1778.000 1089.060 1778.260 1089.320 ;
        RECT 1777.080 1055.400 1777.340 1055.660 ;
        RECT 1778.000 1055.400 1778.260 1055.660 ;
        RECT 1777.080 958.840 1777.340 959.100 ;
        RECT 1777.540 958.840 1777.800 959.100 ;
        RECT 1778.000 910.560 1778.260 910.820 ;
        RECT 1778.000 883.020 1778.260 883.280 ;
        RECT 1778.460 835.080 1778.720 835.340 ;
        RECT 1778.000 821.140 1778.260 821.400 ;
        RECT 1778.000 814.000 1778.260 814.260 ;
        RECT 1777.540 766.060 1777.800 766.320 ;
        RECT 1778.460 641.620 1778.720 641.880 ;
        RECT 1778.460 620.880 1778.720 621.140 ;
        RECT 1778.000 565.460 1778.260 565.720 ;
        RECT 1778.460 517.520 1778.720 517.780 ;
        RECT 1778.460 468.900 1778.720 469.160 ;
        RECT 1778.460 420.960 1778.720 421.220 ;
        RECT 1778.460 324.060 1778.720 324.320 ;
        RECT 1778.000 241.440 1778.260 241.700 ;
        RECT 1778.460 137.740 1778.720 138.000 ;
        RECT 1777.540 89.800 1777.800 90.060 ;
        RECT 1777.540 65.660 1777.800 65.920 ;
        RECT 2691.100 65.660 2691.360 65.920 ;
        RECT 2691.100 2.420 2691.360 2.680 ;
        RECT 2696.620 2.420 2696.880 2.680 ;
      LAYER met2 ;
        RECT 1775.150 1100.580 1775.430 1104.000 ;
        RECT 1775.150 1100.000 1775.440 1100.580 ;
        RECT 1775.300 1089.350 1775.440 1100.000 ;
        RECT 1775.240 1089.030 1775.500 1089.350 ;
        RECT 1778.000 1089.030 1778.260 1089.350 ;
        RECT 1778.060 1055.690 1778.200 1089.030 ;
        RECT 1777.080 1055.370 1777.340 1055.690 ;
        RECT 1778.000 1055.370 1778.260 1055.690 ;
        RECT 1777.140 1007.605 1777.280 1055.370 ;
        RECT 1777.070 1007.235 1777.350 1007.605 ;
        RECT 1778.450 1007.235 1778.730 1007.605 ;
        RECT 1778.520 966.125 1778.660 1007.235 ;
        RECT 1777.070 965.755 1777.350 966.125 ;
        RECT 1778.450 965.755 1778.730 966.125 ;
        RECT 1777.140 959.130 1777.280 965.755 ;
        RECT 1777.080 958.810 1777.340 959.130 ;
        RECT 1777.540 958.810 1777.800 959.130 ;
        RECT 1777.600 910.930 1777.740 958.810 ;
        RECT 1777.600 910.850 1778.200 910.930 ;
        RECT 1777.600 910.790 1778.260 910.850 ;
        RECT 1778.000 910.530 1778.260 910.790 ;
        RECT 1778.000 882.990 1778.260 883.310 ;
        RECT 1778.060 862.650 1778.200 882.990 ;
        RECT 1778.060 862.510 1778.660 862.650 ;
        RECT 1778.520 835.370 1778.660 862.510 ;
        RECT 1778.460 835.050 1778.720 835.370 ;
        RECT 1778.000 821.110 1778.260 821.430 ;
        RECT 1778.060 814.290 1778.200 821.110 ;
        RECT 1778.000 813.970 1778.260 814.290 ;
        RECT 1777.540 766.030 1777.800 766.350 ;
        RECT 1777.600 724.725 1777.740 766.030 ;
        RECT 1777.530 724.355 1777.810 724.725 ;
        RECT 1778.450 724.355 1778.730 724.725 ;
        RECT 1778.520 641.910 1778.660 724.355 ;
        RECT 1778.460 641.590 1778.720 641.910 ;
        RECT 1778.460 620.850 1778.720 621.170 ;
        RECT 1778.520 572.290 1778.660 620.850 ;
        RECT 1778.060 572.150 1778.660 572.290 ;
        RECT 1778.060 565.750 1778.200 572.150 ;
        RECT 1778.000 565.430 1778.260 565.750 ;
        RECT 1778.460 517.490 1778.720 517.810 ;
        RECT 1778.520 469.190 1778.660 517.490 ;
        RECT 1778.460 468.870 1778.720 469.190 ;
        RECT 1778.460 420.930 1778.720 421.250 ;
        RECT 1778.520 397.530 1778.660 420.930 ;
        RECT 1778.060 397.390 1778.660 397.530 ;
        RECT 1778.060 355.370 1778.200 397.390 ;
        RECT 1778.060 355.230 1778.660 355.370 ;
        RECT 1778.520 324.350 1778.660 355.230 ;
        RECT 1778.460 324.030 1778.720 324.350 ;
        RECT 1778.000 241.410 1778.260 241.730 ;
        RECT 1778.060 193.530 1778.200 241.410 ;
        RECT 1778.060 193.390 1778.660 193.530 ;
        RECT 1778.520 138.030 1778.660 193.390 ;
        RECT 1778.460 137.710 1778.720 138.030 ;
        RECT 1777.540 89.770 1777.800 90.090 ;
        RECT 1777.600 65.950 1777.740 89.770 ;
        RECT 1777.540 65.630 1777.800 65.950 ;
        RECT 2691.100 65.630 2691.360 65.950 ;
        RECT 2691.160 2.710 2691.300 65.630 ;
        RECT 2691.100 2.390 2691.360 2.710 ;
        RECT 2696.620 2.390 2696.880 2.710 ;
        RECT 2696.680 2.000 2696.820 2.390 ;
        RECT 2696.470 -4.000 2697.030 2.000 ;
      LAYER via2 ;
        RECT 1777.070 1007.280 1777.350 1007.560 ;
        RECT 1778.450 1007.280 1778.730 1007.560 ;
        RECT 1777.070 965.800 1777.350 966.080 ;
        RECT 1778.450 965.800 1778.730 966.080 ;
        RECT 1777.530 724.400 1777.810 724.680 ;
        RECT 1778.450 724.400 1778.730 724.680 ;
      LAYER met3 ;
        RECT 1777.045 1007.570 1777.375 1007.585 ;
        RECT 1778.425 1007.570 1778.755 1007.585 ;
        RECT 1777.045 1007.270 1778.755 1007.570 ;
        RECT 1777.045 1007.255 1777.375 1007.270 ;
        RECT 1778.425 1007.255 1778.755 1007.270 ;
        RECT 1777.045 966.090 1777.375 966.105 ;
        RECT 1778.425 966.090 1778.755 966.105 ;
        RECT 1777.045 965.790 1778.755 966.090 ;
        RECT 1777.045 965.775 1777.375 965.790 ;
        RECT 1778.425 965.775 1778.755 965.790 ;
        RECT 1777.505 724.690 1777.835 724.705 ;
        RECT 1778.425 724.690 1778.755 724.705 ;
        RECT 1777.505 724.390 1778.755 724.690 ;
        RECT 1777.505 724.375 1777.835 724.390 ;
        RECT 1778.425 724.375 1778.755 724.390 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1781.650 1088.580 1781.970 1088.640 ;
        RECT 1785.790 1088.580 1786.110 1088.640 ;
        RECT 1781.650 1088.440 1786.110 1088.580 ;
        RECT 1781.650 1088.380 1781.970 1088.440 ;
        RECT 1785.790 1088.380 1786.110 1088.440 ;
        RECT 1785.790 65.520 1786.110 65.580 ;
        RECT 2711.770 65.520 2712.090 65.580 ;
        RECT 1785.790 65.380 2712.090 65.520 ;
        RECT 1785.790 65.320 1786.110 65.380 ;
        RECT 2711.770 65.320 2712.090 65.380 ;
      LAYER via ;
        RECT 1781.680 1088.380 1781.940 1088.640 ;
        RECT 1785.820 1088.380 1786.080 1088.640 ;
        RECT 1785.820 65.320 1786.080 65.580 ;
        RECT 2711.800 65.320 2712.060 65.580 ;
      LAYER met2 ;
        RECT 1781.590 1100.580 1781.870 1104.000 ;
        RECT 1781.590 1100.000 1781.880 1100.580 ;
        RECT 1781.740 1088.670 1781.880 1100.000 ;
        RECT 1781.680 1088.350 1781.940 1088.670 ;
        RECT 1785.820 1088.350 1786.080 1088.670 ;
        RECT 1785.880 65.610 1786.020 1088.350 ;
        RECT 1785.820 65.290 1786.080 65.610 ;
        RECT 2711.800 65.290 2712.060 65.610 ;
        RECT 2711.860 2.450 2712.000 65.290 ;
        RECT 2711.860 2.310 2714.760 2.450 ;
        RECT 2714.620 2.000 2714.760 2.310 ;
        RECT 2714.410 -4.000 2714.970 2.000 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1787.630 1088.580 1787.950 1088.640 ;
        RECT 1792.690 1088.580 1793.010 1088.640 ;
        RECT 1787.630 1088.440 1793.010 1088.580 ;
        RECT 1787.630 1088.380 1787.950 1088.440 ;
        RECT 1792.690 1088.380 1793.010 1088.440 ;
        RECT 1792.690 72.320 1793.010 72.380 ;
        RECT 2732.470 72.320 2732.790 72.380 ;
        RECT 1792.690 72.180 2732.790 72.320 ;
        RECT 1792.690 72.120 1793.010 72.180 ;
        RECT 2732.470 72.120 2732.790 72.180 ;
      LAYER via ;
        RECT 1787.660 1088.380 1787.920 1088.640 ;
        RECT 1792.720 1088.380 1792.980 1088.640 ;
        RECT 1792.720 72.120 1792.980 72.380 ;
        RECT 2732.500 72.120 2732.760 72.380 ;
      LAYER met2 ;
        RECT 1787.570 1100.580 1787.850 1104.000 ;
        RECT 1787.570 1100.000 1787.860 1100.580 ;
        RECT 1787.720 1088.670 1787.860 1100.000 ;
        RECT 1787.660 1088.350 1787.920 1088.670 ;
        RECT 1792.720 1088.350 1792.980 1088.670 ;
        RECT 1792.780 72.410 1792.920 1088.350 ;
        RECT 1792.720 72.090 1792.980 72.410 ;
        RECT 2732.500 72.090 2732.760 72.410 ;
        RECT 2732.560 2.000 2732.700 72.090 ;
        RECT 2732.350 -4.000 2732.910 2.000 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1793.610 1089.940 1793.930 1090.000 ;
        RECT 2349.290 1089.940 2349.610 1090.000 ;
        RECT 1793.610 1089.800 2349.610 1089.940 ;
        RECT 1793.610 1089.740 1793.930 1089.800 ;
        RECT 2349.290 1089.740 2349.610 1089.800 ;
        RECT 2349.290 20.640 2349.610 20.700 ;
        RECT 2750.410 20.640 2750.730 20.700 ;
        RECT 2349.290 20.500 2750.730 20.640 ;
        RECT 2349.290 20.440 2349.610 20.500 ;
        RECT 2750.410 20.440 2750.730 20.500 ;
      LAYER via ;
        RECT 1793.640 1089.740 1793.900 1090.000 ;
        RECT 2349.320 1089.740 2349.580 1090.000 ;
        RECT 2349.320 20.440 2349.580 20.700 ;
        RECT 2750.440 20.440 2750.700 20.700 ;
      LAYER met2 ;
        RECT 1793.550 1100.580 1793.830 1104.000 ;
        RECT 1793.550 1100.000 1793.840 1100.580 ;
        RECT 1793.700 1090.030 1793.840 1100.000 ;
        RECT 1793.640 1089.710 1793.900 1090.030 ;
        RECT 2349.320 1089.710 2349.580 1090.030 ;
        RECT 2349.380 20.730 2349.520 1089.710 ;
        RECT 2349.320 20.410 2349.580 20.730 ;
        RECT 2750.440 20.410 2750.700 20.730 ;
        RECT 2750.500 2.000 2750.640 20.410 ;
        RECT 2750.290 -4.000 2750.850 2.000 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1800.510 18.600 1800.830 18.660 ;
        RECT 2767.890 18.600 2768.210 18.660 ;
        RECT 1800.510 18.460 2768.210 18.600 ;
        RECT 1800.510 18.400 1800.830 18.460 ;
        RECT 2767.890 18.400 2768.210 18.460 ;
      LAYER via ;
        RECT 1800.540 18.400 1800.800 18.660 ;
        RECT 2767.920 18.400 2768.180 18.660 ;
      LAYER met2 ;
        RECT 1799.990 1100.650 1800.270 1104.000 ;
        RECT 1799.990 1100.510 1800.740 1100.650 ;
        RECT 1799.990 1100.000 1800.270 1100.510 ;
        RECT 1800.600 18.690 1800.740 1100.510 ;
        RECT 1800.540 18.370 1800.800 18.690 ;
        RECT 2767.920 18.370 2768.180 18.690 ;
        RECT 2767.980 2.000 2768.120 18.370 ;
        RECT 2767.770 -4.000 2768.330 2.000 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 840.950 27.780 841.270 27.840 ;
        RECT 1139.030 27.780 1139.350 27.840 ;
        RECT 840.950 27.640 1139.350 27.780 ;
        RECT 840.950 27.580 841.270 27.640 ;
        RECT 1139.030 27.580 1139.350 27.640 ;
      LAYER via ;
        RECT 840.980 27.580 841.240 27.840 ;
        RECT 1139.060 27.580 1139.320 27.840 ;
      LAYER met2 ;
        RECT 1138.510 1100.650 1138.790 1104.000 ;
        RECT 1138.510 1100.510 1139.260 1100.650 ;
        RECT 1138.510 1100.000 1138.790 1100.510 ;
        RECT 1139.120 27.870 1139.260 1100.510 ;
        RECT 840.980 27.550 841.240 27.870 ;
        RECT 1139.060 27.550 1139.320 27.870 ;
        RECT 841.040 2.000 841.180 27.550 ;
        RECT 840.830 -4.000 841.390 2.000 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1848.885 1083.665 1849.055 1088.595 ;
      LAYER mcon ;
        RECT 1848.885 1088.425 1849.055 1088.595 ;
      LAYER met1 ;
        RECT 1848.825 1088.580 1849.115 1088.625 ;
        RECT 2369.990 1088.580 2370.310 1088.640 ;
        RECT 1848.825 1088.440 2370.310 1088.580 ;
        RECT 1848.825 1088.395 1849.115 1088.440 ;
        RECT 2369.990 1088.380 2370.310 1088.440 ;
        RECT 1806.030 1083.820 1806.350 1083.880 ;
        RECT 1848.825 1083.820 1849.115 1083.865 ;
        RECT 1806.030 1083.680 1849.115 1083.820 ;
        RECT 1806.030 1083.620 1806.350 1083.680 ;
        RECT 1848.825 1083.635 1849.115 1083.680 ;
        RECT 2369.990 20.300 2370.310 20.360 ;
        RECT 2785.830 20.300 2786.150 20.360 ;
        RECT 2369.990 20.160 2786.150 20.300 ;
        RECT 2369.990 20.100 2370.310 20.160 ;
        RECT 2785.830 20.100 2786.150 20.160 ;
      LAYER via ;
        RECT 2370.020 1088.380 2370.280 1088.640 ;
        RECT 1806.060 1083.620 1806.320 1083.880 ;
        RECT 2370.020 20.100 2370.280 20.360 ;
        RECT 2785.860 20.100 2786.120 20.360 ;
      LAYER met2 ;
        RECT 1805.970 1100.580 1806.250 1104.000 ;
        RECT 1805.970 1100.000 1806.260 1100.580 ;
        RECT 1806.120 1083.910 1806.260 1100.000 ;
        RECT 2370.020 1088.350 2370.280 1088.670 ;
        RECT 1806.060 1083.590 1806.320 1083.910 ;
        RECT 2370.080 20.390 2370.220 1088.350 ;
        RECT 2370.020 20.070 2370.280 20.390 ;
        RECT 2785.860 20.070 2786.120 20.390 ;
        RECT 2785.920 2.000 2786.060 20.070 ;
        RECT 2785.710 -4.000 2786.270 2.000 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1812.010 1088.580 1812.330 1088.640 ;
        RECT 1814.310 1088.580 1814.630 1088.640 ;
        RECT 1812.010 1088.440 1814.630 1088.580 ;
        RECT 1812.010 1088.380 1812.330 1088.440 ;
        RECT 1814.310 1088.380 1814.630 1088.440 ;
        RECT 1814.310 18.260 1814.630 18.320 ;
        RECT 2803.770 18.260 2804.090 18.320 ;
        RECT 1814.310 18.120 2804.090 18.260 ;
        RECT 1814.310 18.060 1814.630 18.120 ;
        RECT 2803.770 18.060 2804.090 18.120 ;
      LAYER via ;
        RECT 1812.040 1088.380 1812.300 1088.640 ;
        RECT 1814.340 1088.380 1814.600 1088.640 ;
        RECT 1814.340 18.060 1814.600 18.320 ;
        RECT 2803.800 18.060 2804.060 18.320 ;
      LAYER met2 ;
        RECT 1811.950 1100.580 1812.230 1104.000 ;
        RECT 1811.950 1100.000 1812.240 1100.580 ;
        RECT 1812.100 1088.670 1812.240 1100.000 ;
        RECT 1812.040 1088.350 1812.300 1088.670 ;
        RECT 1814.340 1088.350 1814.600 1088.670 ;
        RECT 1814.400 18.350 1814.540 1088.350 ;
        RECT 1814.340 18.030 1814.600 18.350 ;
        RECT 2803.800 18.030 2804.060 18.350 ;
        RECT 2803.860 2.000 2804.000 18.030 ;
        RECT 2803.650 -4.000 2804.210 2.000 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1818.450 1089.260 1818.770 1089.320 ;
        RECT 2376.890 1089.260 2377.210 1089.320 ;
        RECT 1818.450 1089.120 2377.210 1089.260 ;
        RECT 1818.450 1089.060 1818.770 1089.120 ;
        RECT 2376.890 1089.060 2377.210 1089.120 ;
        RECT 2376.890 19.960 2377.210 20.020 ;
        RECT 2821.710 19.960 2822.030 20.020 ;
        RECT 2376.890 19.820 2822.030 19.960 ;
        RECT 2376.890 19.760 2377.210 19.820 ;
        RECT 2821.710 19.760 2822.030 19.820 ;
      LAYER via ;
        RECT 1818.480 1089.060 1818.740 1089.320 ;
        RECT 2376.920 1089.060 2377.180 1089.320 ;
        RECT 2376.920 19.760 2377.180 20.020 ;
        RECT 2821.740 19.760 2822.000 20.020 ;
      LAYER met2 ;
        RECT 1818.390 1100.580 1818.670 1104.000 ;
        RECT 1818.390 1100.000 1818.680 1100.580 ;
        RECT 1818.540 1089.350 1818.680 1100.000 ;
        RECT 1818.480 1089.030 1818.740 1089.350 ;
        RECT 2376.920 1089.030 2377.180 1089.350 ;
        RECT 2376.980 20.050 2377.120 1089.030 ;
        RECT 2376.920 19.730 2377.180 20.050 ;
        RECT 2821.740 19.730 2822.000 20.050 ;
        RECT 2821.800 2.000 2821.940 19.730 ;
        RECT 2821.590 -4.000 2822.150 2.000 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1824.430 1088.920 1824.750 1088.980 ;
        RECT 1828.110 1088.920 1828.430 1088.980 ;
        RECT 1824.430 1088.780 1828.430 1088.920 ;
        RECT 1824.430 1088.720 1824.750 1088.780 ;
        RECT 1828.110 1088.720 1828.430 1088.780 ;
        RECT 1828.110 17.920 1828.430 17.980 ;
        RECT 2839.190 17.920 2839.510 17.980 ;
        RECT 1828.110 17.780 2839.510 17.920 ;
        RECT 1828.110 17.720 1828.430 17.780 ;
        RECT 2839.190 17.720 2839.510 17.780 ;
      LAYER via ;
        RECT 1824.460 1088.720 1824.720 1088.980 ;
        RECT 1828.140 1088.720 1828.400 1088.980 ;
        RECT 1828.140 17.720 1828.400 17.980 ;
        RECT 2839.220 17.720 2839.480 17.980 ;
      LAYER met2 ;
        RECT 1824.370 1100.580 1824.650 1104.000 ;
        RECT 1824.370 1100.000 1824.660 1100.580 ;
        RECT 1824.520 1089.010 1824.660 1100.000 ;
        RECT 1824.460 1088.690 1824.720 1089.010 ;
        RECT 1828.140 1088.690 1828.400 1089.010 ;
        RECT 1828.200 18.010 1828.340 1088.690 ;
        RECT 1828.140 17.690 1828.400 18.010 ;
        RECT 2839.220 17.690 2839.480 18.010 ;
        RECT 2839.280 2.000 2839.420 17.690 ;
        RECT 2839.070 -4.000 2839.630 2.000 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1830.410 1089.600 1830.730 1089.660 ;
        RECT 2390.690 1089.600 2391.010 1089.660 ;
        RECT 1830.410 1089.460 2391.010 1089.600 ;
        RECT 1830.410 1089.400 1830.730 1089.460 ;
        RECT 2390.690 1089.400 2391.010 1089.460 ;
        RECT 2390.690 19.620 2391.010 19.680 ;
        RECT 2857.130 19.620 2857.450 19.680 ;
        RECT 2390.690 19.480 2857.450 19.620 ;
        RECT 2390.690 19.420 2391.010 19.480 ;
        RECT 2857.130 19.420 2857.450 19.480 ;
      LAYER via ;
        RECT 1830.440 1089.400 1830.700 1089.660 ;
        RECT 2390.720 1089.400 2390.980 1089.660 ;
        RECT 2390.720 19.420 2390.980 19.680 ;
        RECT 2857.160 19.420 2857.420 19.680 ;
      LAYER met2 ;
        RECT 1830.350 1100.580 1830.630 1104.000 ;
        RECT 1830.350 1100.000 1830.640 1100.580 ;
        RECT 1830.500 1089.690 1830.640 1100.000 ;
        RECT 1830.440 1089.370 1830.700 1089.690 ;
        RECT 2390.720 1089.370 2390.980 1089.690 ;
        RECT 2390.780 19.710 2390.920 1089.370 ;
        RECT 2390.720 19.390 2390.980 19.710 ;
        RECT 2857.160 19.390 2857.420 19.710 ;
        RECT 2857.220 2.000 2857.360 19.390 ;
        RECT 2857.010 -4.000 2857.570 2.000 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1836.390 1088.920 1836.710 1088.980 ;
        RECT 1841.910 1088.920 1842.230 1088.980 ;
        RECT 1836.390 1088.780 1842.230 1088.920 ;
        RECT 1836.390 1088.720 1836.710 1088.780 ;
        RECT 1841.910 1088.720 1842.230 1088.780 ;
        RECT 1841.910 17.580 1842.230 17.640 ;
        RECT 2875.070 17.580 2875.390 17.640 ;
        RECT 1841.910 17.440 2875.390 17.580 ;
        RECT 1841.910 17.380 1842.230 17.440 ;
        RECT 2875.070 17.380 2875.390 17.440 ;
      LAYER via ;
        RECT 1836.420 1088.720 1836.680 1088.980 ;
        RECT 1841.940 1088.720 1842.200 1088.980 ;
        RECT 1841.940 17.380 1842.200 17.640 ;
        RECT 2875.100 17.380 2875.360 17.640 ;
      LAYER met2 ;
        RECT 1836.330 1100.580 1836.610 1104.000 ;
        RECT 1836.330 1100.000 1836.620 1100.580 ;
        RECT 1836.480 1089.010 1836.620 1100.000 ;
        RECT 1836.420 1088.690 1836.680 1089.010 ;
        RECT 1841.940 1088.690 1842.200 1089.010 ;
        RECT 1842.000 17.670 1842.140 1088.690 ;
        RECT 1841.940 17.350 1842.200 17.670 ;
        RECT 2875.100 17.350 2875.360 17.670 ;
        RECT 2875.160 2.000 2875.300 17.350 ;
        RECT 2874.950 -4.000 2875.510 2.000 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1842.830 1088.920 1843.150 1088.980 ;
        RECT 2404.490 1088.920 2404.810 1088.980 ;
        RECT 1842.830 1088.780 2404.810 1088.920 ;
        RECT 1842.830 1088.720 1843.150 1088.780 ;
        RECT 2404.490 1088.720 2404.810 1088.780 ;
        RECT 2404.490 19.280 2404.810 19.340 ;
        RECT 2893.010 19.280 2893.330 19.340 ;
        RECT 2404.490 19.140 2893.330 19.280 ;
        RECT 2404.490 19.080 2404.810 19.140 ;
        RECT 2893.010 19.080 2893.330 19.140 ;
      LAYER via ;
        RECT 1842.860 1088.720 1843.120 1088.980 ;
        RECT 2404.520 1088.720 2404.780 1088.980 ;
        RECT 2404.520 19.080 2404.780 19.340 ;
        RECT 2893.040 19.080 2893.300 19.340 ;
      LAYER met2 ;
        RECT 1842.770 1100.580 1843.050 1104.000 ;
        RECT 1842.770 1100.000 1843.060 1100.580 ;
        RECT 1842.920 1089.010 1843.060 1100.000 ;
        RECT 1842.860 1088.690 1843.120 1089.010 ;
        RECT 2404.520 1088.690 2404.780 1089.010 ;
        RECT 2404.580 19.370 2404.720 1088.690 ;
        RECT 2404.520 19.050 2404.780 19.370 ;
        RECT 2893.040 19.050 2893.300 19.370 ;
        RECT 2893.100 2.000 2893.240 19.050 ;
        RECT 2892.890 -4.000 2893.450 2.000 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1848.810 17.240 1849.130 17.300 ;
        RECT 2910.950 17.240 2911.270 17.300 ;
        RECT 1848.810 17.100 2911.270 17.240 ;
        RECT 1848.810 17.040 1849.130 17.100 ;
        RECT 2910.950 17.040 2911.270 17.100 ;
      LAYER via ;
        RECT 1848.840 17.040 1849.100 17.300 ;
        RECT 2910.980 17.040 2911.240 17.300 ;
      LAYER met2 ;
        RECT 1848.750 1100.580 1849.030 1104.000 ;
        RECT 1848.750 1100.000 1849.040 1100.580 ;
        RECT 1848.900 17.330 1849.040 1100.000 ;
        RECT 1848.840 17.010 1849.100 17.330 ;
        RECT 2910.980 17.010 2911.240 17.330 ;
        RECT 2911.040 2.000 2911.180 17.010 ;
        RECT 2910.830 -4.000 2911.390 2.000 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1139.490 1052.200 1139.810 1052.260 ;
        RECT 1143.170 1052.200 1143.490 1052.260 ;
        RECT 1139.490 1052.060 1143.490 1052.200 ;
        RECT 1139.490 1052.000 1139.810 1052.060 ;
        RECT 1143.170 1052.000 1143.490 1052.060 ;
        RECT 858.890 30.840 859.210 30.900 ;
        RECT 1139.490 30.840 1139.810 30.900 ;
        RECT 858.890 30.700 1139.810 30.840 ;
        RECT 858.890 30.640 859.210 30.700 ;
        RECT 1139.490 30.640 1139.810 30.700 ;
      LAYER via ;
        RECT 1139.520 1052.000 1139.780 1052.260 ;
        RECT 1143.200 1052.000 1143.460 1052.260 ;
        RECT 858.920 30.640 859.180 30.900 ;
        RECT 1139.520 30.640 1139.780 30.900 ;
      LAYER met2 ;
        RECT 1144.490 1100.650 1144.770 1104.000 ;
        RECT 1143.260 1100.510 1144.770 1100.650 ;
        RECT 1143.260 1052.290 1143.400 1100.510 ;
        RECT 1144.490 1100.000 1144.770 1100.510 ;
        RECT 1139.520 1051.970 1139.780 1052.290 ;
        RECT 1143.200 1051.970 1143.460 1052.290 ;
        RECT 1139.580 30.930 1139.720 1051.970 ;
        RECT 858.920 30.610 859.180 30.930 ;
        RECT 1139.520 30.610 1139.780 30.930 ;
        RECT 858.980 2.000 859.120 30.610 ;
        RECT 858.770 -4.000 859.330 2.000 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1145.930 1035.200 1146.250 1035.260 ;
        RECT 1149.150 1035.200 1149.470 1035.260 ;
        RECT 1145.930 1035.060 1149.470 1035.200 ;
        RECT 1145.930 1035.000 1146.250 1035.060 ;
        RECT 1149.150 1035.000 1149.470 1035.060 ;
        RECT 876.830 31.180 877.150 31.240 ;
        RECT 1145.930 31.180 1146.250 31.240 ;
        RECT 876.830 31.040 1146.250 31.180 ;
        RECT 876.830 30.980 877.150 31.040 ;
        RECT 1145.930 30.980 1146.250 31.040 ;
      LAYER via ;
        RECT 1145.960 1035.000 1146.220 1035.260 ;
        RECT 1149.180 1035.000 1149.440 1035.260 ;
        RECT 876.860 30.980 877.120 31.240 ;
        RECT 1145.960 30.980 1146.220 31.240 ;
      LAYER met2 ;
        RECT 1150.930 1100.650 1151.210 1104.000 ;
        RECT 1149.240 1100.510 1151.210 1100.650 ;
        RECT 1149.240 1035.290 1149.380 1100.510 ;
        RECT 1150.930 1100.000 1151.210 1100.510 ;
        RECT 1145.960 1034.970 1146.220 1035.290 ;
        RECT 1149.180 1034.970 1149.440 1035.290 ;
        RECT 1146.020 31.270 1146.160 1034.970 ;
        RECT 876.860 30.950 877.120 31.270 ;
        RECT 1145.960 30.950 1146.220 31.270 ;
        RECT 876.920 2.000 877.060 30.950 ;
        RECT 876.710 -4.000 877.270 2.000 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1152.370 1052.200 1152.690 1052.260 ;
        RECT 1155.590 1052.200 1155.910 1052.260 ;
        RECT 1152.370 1052.060 1155.910 1052.200 ;
        RECT 1152.370 1052.000 1152.690 1052.060 ;
        RECT 1155.590 1052.000 1155.910 1052.060 ;
        RECT 894.770 31.520 895.090 31.580 ;
        RECT 1152.370 31.520 1152.690 31.580 ;
        RECT 894.770 31.380 1152.690 31.520 ;
        RECT 894.770 31.320 895.090 31.380 ;
        RECT 1152.370 31.320 1152.690 31.380 ;
      LAYER via ;
        RECT 1152.400 1052.000 1152.660 1052.260 ;
        RECT 1155.620 1052.000 1155.880 1052.260 ;
        RECT 894.800 31.320 895.060 31.580 ;
        RECT 1152.400 31.320 1152.660 31.580 ;
      LAYER met2 ;
        RECT 1156.910 1100.650 1157.190 1104.000 ;
        RECT 1155.680 1100.510 1157.190 1100.650 ;
        RECT 1155.680 1052.290 1155.820 1100.510 ;
        RECT 1156.910 1100.000 1157.190 1100.510 ;
        RECT 1152.400 1051.970 1152.660 1052.290 ;
        RECT 1155.620 1051.970 1155.880 1052.290 ;
        RECT 1152.460 31.610 1152.600 1051.970 ;
        RECT 894.800 31.290 895.060 31.610 ;
        RECT 1152.400 31.290 1152.660 31.610 ;
        RECT 894.860 2.000 895.000 31.290 ;
        RECT 894.650 -4.000 895.210 2.000 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1161.185 565.845 1161.355 613.955 ;
        RECT 1161.185 379.525 1161.355 386.495 ;
        RECT 1160.265 186.405 1160.435 234.515 ;
      LAYER mcon ;
        RECT 1161.185 613.785 1161.355 613.955 ;
        RECT 1161.185 386.325 1161.355 386.495 ;
        RECT 1160.265 234.345 1160.435 234.515 ;
      LAYER met1 ;
        RECT 1160.650 1014.460 1160.970 1014.520 ;
        RECT 1161.570 1014.460 1161.890 1014.520 ;
        RECT 1160.650 1014.320 1161.890 1014.460 ;
        RECT 1160.650 1014.260 1160.970 1014.320 ;
        RECT 1161.570 1014.260 1161.890 1014.320 ;
        RECT 1160.650 990.660 1160.970 990.720 ;
        RECT 1160.280 990.520 1160.970 990.660 ;
        RECT 1160.280 990.380 1160.420 990.520 ;
        RECT 1160.650 990.460 1160.970 990.520 ;
        RECT 1160.190 990.120 1160.510 990.380 ;
        RECT 1160.650 917.900 1160.970 917.960 ;
        RECT 1161.110 917.900 1161.430 917.960 ;
        RECT 1160.650 917.760 1161.430 917.900 ;
        RECT 1160.650 917.700 1160.970 917.760 ;
        RECT 1161.110 917.700 1161.430 917.760 ;
        RECT 1160.650 869.960 1160.970 870.020 ;
        RECT 1161.110 869.960 1161.430 870.020 ;
        RECT 1160.650 869.820 1161.430 869.960 ;
        RECT 1160.650 869.760 1160.970 869.820 ;
        RECT 1161.110 869.760 1161.430 869.820 ;
        RECT 1160.650 835.420 1160.970 835.680 ;
        RECT 1160.740 835.000 1160.880 835.420 ;
        RECT 1160.650 834.740 1160.970 835.000 ;
        RECT 1160.650 786.320 1160.970 786.380 ;
        RECT 1160.280 786.180 1160.970 786.320 ;
        RECT 1160.280 785.700 1160.420 786.180 ;
        RECT 1160.650 786.120 1160.970 786.180 ;
        RECT 1160.190 785.440 1160.510 785.700 ;
        RECT 1158.810 765.920 1159.130 765.980 ;
        RECT 1160.190 765.920 1160.510 765.980 ;
        RECT 1158.810 765.780 1160.510 765.920 ;
        RECT 1158.810 765.720 1159.130 765.780 ;
        RECT 1160.190 765.720 1160.510 765.780 ;
        RECT 1160.190 696.220 1160.510 696.280 ;
        RECT 1161.570 696.220 1161.890 696.280 ;
        RECT 1160.190 696.080 1161.890 696.220 ;
        RECT 1160.190 696.020 1160.510 696.080 ;
        RECT 1161.570 696.020 1161.890 696.080 ;
        RECT 1161.110 621.080 1161.430 621.140 ;
        RECT 1161.570 621.080 1161.890 621.140 ;
        RECT 1161.110 620.940 1161.890 621.080 ;
        RECT 1161.110 620.880 1161.430 620.940 ;
        RECT 1161.570 620.880 1161.890 620.940 ;
        RECT 1161.125 613.940 1161.415 613.985 ;
        RECT 1161.570 613.940 1161.890 614.000 ;
        RECT 1161.125 613.800 1161.890 613.940 ;
        RECT 1161.125 613.755 1161.415 613.800 ;
        RECT 1161.570 613.740 1161.890 613.800 ;
        RECT 1161.110 566.000 1161.430 566.060 ;
        RECT 1160.915 565.860 1161.430 566.000 ;
        RECT 1161.110 565.800 1161.430 565.860 ;
        RECT 1160.190 483.040 1160.510 483.100 ;
        RECT 1161.110 483.040 1161.430 483.100 ;
        RECT 1160.190 482.900 1161.430 483.040 ;
        RECT 1160.190 482.840 1160.510 482.900 ;
        RECT 1161.110 482.840 1161.430 482.900 ;
        RECT 1161.110 386.480 1161.430 386.540 ;
        RECT 1160.915 386.340 1161.430 386.480 ;
        RECT 1161.110 386.280 1161.430 386.340 ;
        RECT 1161.110 379.680 1161.430 379.740 ;
        RECT 1160.915 379.540 1161.430 379.680 ;
        RECT 1161.110 379.480 1161.430 379.540 ;
        RECT 1160.190 338.200 1160.510 338.260 ;
        RECT 1161.110 338.200 1161.430 338.260 ;
        RECT 1160.190 338.060 1161.430 338.200 ;
        RECT 1160.190 338.000 1160.510 338.060 ;
        RECT 1161.110 338.000 1161.430 338.060 ;
        RECT 1160.650 255.580 1160.970 255.640 ;
        RECT 1160.280 255.440 1160.970 255.580 ;
        RECT 1160.280 255.300 1160.420 255.440 ;
        RECT 1160.650 255.380 1160.970 255.440 ;
        RECT 1160.190 255.040 1160.510 255.300 ;
        RECT 1160.190 234.500 1160.510 234.560 ;
        RECT 1159.995 234.360 1160.510 234.500 ;
        RECT 1160.190 234.300 1160.510 234.360 ;
        RECT 1160.190 186.560 1160.510 186.620 ;
        RECT 1159.995 186.420 1160.510 186.560 ;
        RECT 1160.190 186.360 1160.510 186.420 ;
        RECT 1160.190 145.080 1160.510 145.140 ;
        RECT 1160.650 145.080 1160.970 145.140 ;
        RECT 1160.190 144.940 1160.970 145.080 ;
        RECT 1160.190 144.880 1160.510 144.940 ;
        RECT 1160.650 144.880 1160.970 144.940 ;
        RECT 912.710 31.860 913.030 31.920 ;
        RECT 1160.650 31.860 1160.970 31.920 ;
        RECT 912.710 31.720 1160.970 31.860 ;
        RECT 912.710 31.660 913.030 31.720 ;
        RECT 1160.650 31.660 1160.970 31.720 ;
      LAYER via ;
        RECT 1160.680 1014.260 1160.940 1014.520 ;
        RECT 1161.600 1014.260 1161.860 1014.520 ;
        RECT 1160.680 990.460 1160.940 990.720 ;
        RECT 1160.220 990.120 1160.480 990.380 ;
        RECT 1160.680 917.700 1160.940 917.960 ;
        RECT 1161.140 917.700 1161.400 917.960 ;
        RECT 1160.680 869.760 1160.940 870.020 ;
        RECT 1161.140 869.760 1161.400 870.020 ;
        RECT 1160.680 835.420 1160.940 835.680 ;
        RECT 1160.680 834.740 1160.940 835.000 ;
        RECT 1160.680 786.120 1160.940 786.380 ;
        RECT 1160.220 785.440 1160.480 785.700 ;
        RECT 1158.840 765.720 1159.100 765.980 ;
        RECT 1160.220 765.720 1160.480 765.980 ;
        RECT 1160.220 696.020 1160.480 696.280 ;
        RECT 1161.600 696.020 1161.860 696.280 ;
        RECT 1161.140 620.880 1161.400 621.140 ;
        RECT 1161.600 620.880 1161.860 621.140 ;
        RECT 1161.600 613.740 1161.860 614.000 ;
        RECT 1161.140 565.800 1161.400 566.060 ;
        RECT 1160.220 482.840 1160.480 483.100 ;
        RECT 1161.140 482.840 1161.400 483.100 ;
        RECT 1161.140 386.280 1161.400 386.540 ;
        RECT 1161.140 379.480 1161.400 379.740 ;
        RECT 1160.220 338.000 1160.480 338.260 ;
        RECT 1161.140 338.000 1161.400 338.260 ;
        RECT 1160.680 255.380 1160.940 255.640 ;
        RECT 1160.220 255.040 1160.480 255.300 ;
        RECT 1160.220 234.300 1160.480 234.560 ;
        RECT 1160.220 186.360 1160.480 186.620 ;
        RECT 1160.220 144.880 1160.480 145.140 ;
        RECT 1160.680 144.880 1160.940 145.140 ;
        RECT 912.740 31.660 913.000 31.920 ;
        RECT 1160.680 31.660 1160.940 31.920 ;
      LAYER met2 ;
        RECT 1162.890 1100.650 1163.170 1104.000 ;
        RECT 1161.660 1100.510 1163.170 1100.650 ;
        RECT 1161.660 1081.610 1161.800 1100.510 ;
        RECT 1162.890 1100.000 1163.170 1100.510 ;
        RECT 1160.280 1081.470 1161.800 1081.610 ;
        RECT 1160.280 1062.685 1160.420 1081.470 ;
        RECT 1160.210 1062.315 1160.490 1062.685 ;
        RECT 1161.590 1062.315 1161.870 1062.685 ;
        RECT 1161.660 1014.550 1161.800 1062.315 ;
        RECT 1160.680 1014.230 1160.940 1014.550 ;
        RECT 1161.600 1014.230 1161.860 1014.550 ;
        RECT 1160.740 990.750 1160.880 1014.230 ;
        RECT 1160.680 990.430 1160.940 990.750 ;
        RECT 1160.220 990.090 1160.480 990.410 ;
        RECT 1160.280 966.125 1160.420 990.090 ;
        RECT 1160.210 965.755 1160.490 966.125 ;
        RECT 1161.130 965.755 1161.410 966.125 ;
        RECT 1160.740 917.990 1160.880 918.145 ;
        RECT 1161.200 917.990 1161.340 965.755 ;
        RECT 1160.680 917.730 1160.940 917.990 ;
        RECT 1161.140 917.730 1161.400 917.990 ;
        RECT 1160.680 917.670 1161.400 917.730 ;
        RECT 1160.740 917.590 1161.340 917.670 ;
        RECT 1161.200 870.050 1161.340 917.590 ;
        RECT 1160.680 869.730 1160.940 870.050 ;
        RECT 1161.140 869.730 1161.400 870.050 ;
        RECT 1160.740 835.710 1160.880 869.730 ;
        RECT 1160.680 835.390 1160.940 835.710 ;
        RECT 1160.680 834.710 1160.940 835.030 ;
        RECT 1160.740 786.410 1160.880 834.710 ;
        RECT 1160.680 786.090 1160.940 786.410 ;
        RECT 1160.220 785.410 1160.480 785.730 ;
        RECT 1160.280 766.010 1160.420 785.410 ;
        RECT 1158.840 765.690 1159.100 766.010 ;
        RECT 1160.220 765.690 1160.480 766.010 ;
        RECT 1158.900 717.925 1159.040 765.690 ;
        RECT 1158.830 717.555 1159.110 717.925 ;
        RECT 1160.210 717.555 1160.490 717.925 ;
        RECT 1160.280 696.310 1160.420 717.555 ;
        RECT 1160.220 695.990 1160.480 696.310 ;
        RECT 1161.600 695.990 1161.860 696.310 ;
        RECT 1161.660 621.170 1161.800 695.990 ;
        RECT 1161.140 620.850 1161.400 621.170 ;
        RECT 1161.600 620.850 1161.860 621.170 ;
        RECT 1161.200 620.570 1161.340 620.850 ;
        RECT 1161.200 620.430 1161.800 620.570 ;
        RECT 1161.660 614.030 1161.800 620.430 ;
        RECT 1161.600 613.710 1161.860 614.030 ;
        RECT 1161.140 565.770 1161.400 566.090 ;
        RECT 1161.200 496.130 1161.340 565.770 ;
        RECT 1160.280 495.990 1161.340 496.130 ;
        RECT 1160.280 483.130 1160.420 495.990 ;
        RECT 1160.220 482.810 1160.480 483.130 ;
        RECT 1161.140 482.810 1161.400 483.130 ;
        RECT 1161.200 386.570 1161.340 482.810 ;
        RECT 1161.140 386.250 1161.400 386.570 ;
        RECT 1161.140 379.450 1161.400 379.770 ;
        RECT 1161.200 338.290 1161.340 379.450 ;
        RECT 1160.220 337.970 1160.480 338.290 ;
        RECT 1161.140 337.970 1161.400 338.290 ;
        RECT 1160.280 307.090 1160.420 337.970 ;
        RECT 1160.280 306.950 1161.340 307.090 ;
        RECT 1161.200 303.520 1161.340 306.950 ;
        RECT 1160.740 303.380 1161.340 303.520 ;
        RECT 1160.740 255.670 1160.880 303.380 ;
        RECT 1160.680 255.350 1160.940 255.670 ;
        RECT 1160.220 255.010 1160.480 255.330 ;
        RECT 1160.280 234.590 1160.420 255.010 ;
        RECT 1160.220 234.270 1160.480 234.590 ;
        RECT 1160.220 186.330 1160.480 186.650 ;
        RECT 1160.280 145.170 1160.420 186.330 ;
        RECT 1160.220 144.850 1160.480 145.170 ;
        RECT 1160.680 144.850 1160.940 145.170 ;
        RECT 1160.740 31.950 1160.880 144.850 ;
        RECT 912.740 31.630 913.000 31.950 ;
        RECT 1160.680 31.630 1160.940 31.950 ;
        RECT 912.800 2.000 912.940 31.630 ;
        RECT 912.590 -4.000 913.150 2.000 ;
      LAYER via2 ;
        RECT 1160.210 1062.360 1160.490 1062.640 ;
        RECT 1161.590 1062.360 1161.870 1062.640 ;
        RECT 1160.210 965.800 1160.490 966.080 ;
        RECT 1161.130 965.800 1161.410 966.080 ;
        RECT 1158.830 717.600 1159.110 717.880 ;
        RECT 1160.210 717.600 1160.490 717.880 ;
      LAYER met3 ;
        RECT 1160.185 1062.650 1160.515 1062.665 ;
        RECT 1161.565 1062.650 1161.895 1062.665 ;
        RECT 1160.185 1062.350 1161.895 1062.650 ;
        RECT 1160.185 1062.335 1160.515 1062.350 ;
        RECT 1161.565 1062.335 1161.895 1062.350 ;
        RECT 1160.185 966.090 1160.515 966.105 ;
        RECT 1161.105 966.090 1161.435 966.105 ;
        RECT 1160.185 965.790 1161.435 966.090 ;
        RECT 1160.185 965.775 1160.515 965.790 ;
        RECT 1161.105 965.775 1161.435 965.790 ;
        RECT 1158.805 717.890 1159.135 717.905 ;
        RECT 1160.185 717.890 1160.515 717.905 ;
        RECT 1158.805 717.590 1160.515 717.890 ;
        RECT 1158.805 717.575 1159.135 717.590 ;
        RECT 1160.185 717.575 1160.515 717.590 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 930.190 32.200 930.510 32.260 ;
        RECT 1167.550 32.200 1167.870 32.260 ;
        RECT 930.190 32.060 1167.870 32.200 ;
        RECT 930.190 32.000 930.510 32.060 ;
        RECT 1167.550 32.000 1167.870 32.060 ;
      LAYER via ;
        RECT 930.220 32.000 930.480 32.260 ;
        RECT 1167.580 32.000 1167.840 32.260 ;
      LAYER met2 ;
        RECT 1169.330 1100.650 1169.610 1104.000 ;
        RECT 1167.640 1100.510 1169.610 1100.650 ;
        RECT 1167.640 32.290 1167.780 1100.510 ;
        RECT 1169.330 1100.000 1169.610 1100.510 ;
        RECT 930.220 31.970 930.480 32.290 ;
        RECT 1167.580 31.970 1167.840 32.290 ;
        RECT 930.280 2.000 930.420 31.970 ;
        RECT 930.070 -4.000 930.630 2.000 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1173.070 1051.860 1173.390 1051.920 ;
        RECT 1174.450 1051.860 1174.770 1051.920 ;
        RECT 1173.070 1051.720 1174.770 1051.860 ;
        RECT 1173.070 1051.660 1173.390 1051.720 ;
        RECT 1174.450 1051.660 1174.770 1051.720 ;
        RECT 948.130 18.600 948.450 18.660 ;
        RECT 1173.070 18.600 1173.390 18.660 ;
        RECT 948.130 18.460 1173.390 18.600 ;
        RECT 948.130 18.400 948.450 18.460 ;
        RECT 1173.070 18.400 1173.390 18.460 ;
      LAYER via ;
        RECT 1173.100 1051.660 1173.360 1051.920 ;
        RECT 1174.480 1051.660 1174.740 1051.920 ;
        RECT 948.160 18.400 948.420 18.660 ;
        RECT 1173.100 18.400 1173.360 18.660 ;
      LAYER met2 ;
        RECT 1175.310 1100.650 1175.590 1104.000 ;
        RECT 1174.540 1100.510 1175.590 1100.650 ;
        RECT 1174.540 1051.950 1174.680 1100.510 ;
        RECT 1175.310 1100.000 1175.590 1100.510 ;
        RECT 1173.100 1051.630 1173.360 1051.950 ;
        RECT 1174.480 1051.630 1174.740 1051.950 ;
        RECT 1173.160 18.690 1173.300 1051.630 ;
        RECT 948.160 18.370 948.420 18.690 ;
        RECT 1173.100 18.370 1173.360 18.690 ;
        RECT 948.220 2.000 948.360 18.370 ;
        RECT 948.010 -4.000 948.570 2.000 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1125.765 17.425 1125.935 18.955 ;
      LAYER mcon ;
        RECT 1125.765 18.785 1125.935 18.955 ;
      LAYER met1 ;
        RECT 966.070 18.940 966.390 19.000 ;
        RECT 1125.705 18.940 1125.995 18.985 ;
        RECT 966.070 18.800 1125.995 18.940 ;
        RECT 966.070 18.740 966.390 18.800 ;
        RECT 1125.705 18.755 1125.995 18.800 ;
        RECT 1180.430 17.920 1180.750 17.980 ;
        RECT 1176.840 17.780 1180.750 17.920 ;
        RECT 1125.705 17.580 1125.995 17.625 ;
        RECT 1176.840 17.580 1176.980 17.780 ;
        RECT 1180.430 17.720 1180.750 17.780 ;
        RECT 1125.705 17.440 1176.980 17.580 ;
        RECT 1125.705 17.395 1125.995 17.440 ;
      LAYER via ;
        RECT 966.100 18.740 966.360 19.000 ;
        RECT 1180.460 17.720 1180.720 17.980 ;
      LAYER met2 ;
        RECT 1181.290 1100.650 1181.570 1104.000 ;
        RECT 1180.520 1100.510 1181.570 1100.650 ;
        RECT 966.100 18.710 966.360 19.030 ;
        RECT 966.160 2.000 966.300 18.710 ;
        RECT 1180.520 18.010 1180.660 1100.510 ;
        RECT 1181.290 1100.000 1181.570 1100.510 ;
        RECT 1180.460 17.690 1180.720 18.010 ;
        RECT 965.950 -4.000 966.510 2.000 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1024.490 1087.560 1024.810 1087.620 ;
        RECT 1187.790 1087.560 1188.110 1087.620 ;
        RECT 1024.490 1087.420 1188.110 1087.560 ;
        RECT 1024.490 1087.360 1024.810 1087.420 ;
        RECT 1187.790 1087.360 1188.110 1087.420 ;
        RECT 984.010 16.220 984.330 16.280 ;
        RECT 1024.490 16.220 1024.810 16.280 ;
        RECT 984.010 16.080 1024.810 16.220 ;
        RECT 984.010 16.020 984.330 16.080 ;
        RECT 1024.490 16.020 1024.810 16.080 ;
      LAYER via ;
        RECT 1024.520 1087.360 1024.780 1087.620 ;
        RECT 1187.820 1087.360 1188.080 1087.620 ;
        RECT 984.040 16.020 984.300 16.280 ;
        RECT 1024.520 16.020 1024.780 16.280 ;
      LAYER met2 ;
        RECT 1187.730 1100.580 1188.010 1104.000 ;
        RECT 1187.730 1100.000 1188.020 1100.580 ;
        RECT 1187.880 1087.650 1188.020 1100.000 ;
        RECT 1024.520 1087.330 1024.780 1087.650 ;
        RECT 1187.820 1087.330 1188.080 1087.650 ;
        RECT 1024.580 16.310 1024.720 1087.330 ;
        RECT 984.040 15.990 984.300 16.310 ;
        RECT 1024.520 15.990 1024.780 16.310 ;
        RECT 984.100 2.000 984.240 15.990 ;
        RECT 983.890 -4.000 984.450 2.000 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 662.930 30.500 663.250 30.560 ;
        RECT 1076.470 30.500 1076.790 30.560 ;
        RECT 662.930 30.360 1076.790 30.500 ;
        RECT 662.930 30.300 663.250 30.360 ;
        RECT 1076.470 30.300 1076.790 30.360 ;
      LAYER via ;
        RECT 662.960 30.300 663.220 30.560 ;
        RECT 1076.500 30.300 1076.760 30.560 ;
      LAYER met2 ;
        RECT 1077.330 1100.650 1077.610 1104.000 ;
        RECT 1076.560 1100.510 1077.610 1100.650 ;
        RECT 1076.560 30.590 1076.700 1100.510 ;
        RECT 1077.330 1100.000 1077.610 1100.510 ;
        RECT 662.960 30.270 663.220 30.590 ;
        RECT 1076.500 30.270 1076.760 30.590 ;
        RECT 663.020 2.000 663.160 30.270 ;
        RECT 662.810 -4.000 663.370 2.000 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1007.010 1086.540 1007.330 1086.600 ;
        RECT 1193.770 1086.540 1194.090 1086.600 ;
        RECT 1007.010 1086.400 1194.090 1086.540 ;
        RECT 1007.010 1086.340 1007.330 1086.400 ;
        RECT 1193.770 1086.340 1194.090 1086.400 ;
        RECT 1001.950 15.540 1002.270 15.600 ;
        RECT 1007.010 15.540 1007.330 15.600 ;
        RECT 1001.950 15.400 1007.330 15.540 ;
        RECT 1001.950 15.340 1002.270 15.400 ;
        RECT 1007.010 15.340 1007.330 15.400 ;
      LAYER via ;
        RECT 1007.040 1086.340 1007.300 1086.600 ;
        RECT 1193.800 1086.340 1194.060 1086.600 ;
        RECT 1001.980 15.340 1002.240 15.600 ;
        RECT 1007.040 15.340 1007.300 15.600 ;
      LAYER met2 ;
        RECT 1193.710 1100.580 1193.990 1104.000 ;
        RECT 1193.710 1100.000 1194.000 1100.580 ;
        RECT 1193.860 1086.630 1194.000 1100.000 ;
        RECT 1007.040 1086.310 1007.300 1086.630 ;
        RECT 1193.800 1086.310 1194.060 1086.630 ;
        RECT 1007.100 15.630 1007.240 1086.310 ;
        RECT 1001.980 15.310 1002.240 15.630 ;
        RECT 1007.040 15.310 1007.300 15.630 ;
        RECT 1002.040 2.000 1002.180 15.310 ;
        RECT 1001.830 -4.000 1002.390 2.000 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1020.810 1086.880 1021.130 1086.940 ;
        RECT 1199.750 1086.880 1200.070 1086.940 ;
        RECT 1020.810 1086.740 1200.070 1086.880 ;
        RECT 1020.810 1086.680 1021.130 1086.740 ;
        RECT 1199.750 1086.680 1200.070 1086.740 ;
      LAYER via ;
        RECT 1020.840 1086.680 1021.100 1086.940 ;
        RECT 1199.780 1086.680 1200.040 1086.940 ;
      LAYER met2 ;
        RECT 1199.690 1100.580 1199.970 1104.000 ;
        RECT 1199.690 1100.000 1199.980 1100.580 ;
        RECT 1199.840 1086.970 1199.980 1100.000 ;
        RECT 1020.840 1086.650 1021.100 1086.970 ;
        RECT 1199.780 1086.650 1200.040 1086.970 ;
        RECT 1020.900 2.450 1021.040 1086.650 ;
        RECT 1019.520 2.310 1021.040 2.450 ;
        RECT 1019.520 2.000 1019.660 2.310 ;
        RECT 1019.310 -4.000 1019.870 2.000 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1041.510 1087.900 1041.830 1087.960 ;
        RECT 1205.730 1087.900 1206.050 1087.960 ;
        RECT 1041.510 1087.760 1206.050 1087.900 ;
        RECT 1041.510 1087.700 1041.830 1087.760 ;
        RECT 1205.730 1087.700 1206.050 1087.760 ;
        RECT 1037.370 15.880 1037.690 15.940 ;
        RECT 1041.510 15.880 1041.830 15.940 ;
        RECT 1037.370 15.740 1041.830 15.880 ;
        RECT 1037.370 15.680 1037.690 15.740 ;
        RECT 1041.510 15.680 1041.830 15.740 ;
      LAYER via ;
        RECT 1041.540 1087.700 1041.800 1087.960 ;
        RECT 1205.760 1087.700 1206.020 1087.960 ;
        RECT 1037.400 15.680 1037.660 15.940 ;
        RECT 1041.540 15.680 1041.800 15.940 ;
      LAYER met2 ;
        RECT 1205.670 1100.580 1205.950 1104.000 ;
        RECT 1205.670 1100.000 1205.960 1100.580 ;
        RECT 1205.820 1087.990 1205.960 1100.000 ;
        RECT 1041.540 1087.670 1041.800 1087.990 ;
        RECT 1205.760 1087.670 1206.020 1087.990 ;
        RECT 1041.600 15.970 1041.740 1087.670 ;
        RECT 1037.400 15.650 1037.660 15.970 ;
        RECT 1041.540 15.650 1041.800 15.970 ;
        RECT 1037.460 2.000 1037.600 15.650 ;
        RECT 1037.250 -4.000 1037.810 2.000 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1061.290 1088.240 1061.610 1088.300 ;
        RECT 1212.170 1088.240 1212.490 1088.300 ;
        RECT 1061.290 1088.100 1212.490 1088.240 ;
        RECT 1061.290 1088.040 1061.610 1088.100 ;
        RECT 1212.170 1088.040 1212.490 1088.100 ;
        RECT 1058.990 1083.480 1059.310 1083.540 ;
        RECT 1061.290 1083.480 1061.610 1083.540 ;
        RECT 1058.990 1083.340 1061.610 1083.480 ;
        RECT 1058.990 1083.280 1059.310 1083.340 ;
        RECT 1061.290 1083.280 1061.610 1083.340 ;
        RECT 1055.310 20.640 1055.630 20.700 ;
        RECT 1058.990 20.640 1059.310 20.700 ;
        RECT 1055.310 20.500 1059.310 20.640 ;
        RECT 1055.310 20.440 1055.630 20.500 ;
        RECT 1058.990 20.440 1059.310 20.500 ;
      LAYER via ;
        RECT 1061.320 1088.040 1061.580 1088.300 ;
        RECT 1212.200 1088.040 1212.460 1088.300 ;
        RECT 1059.020 1083.280 1059.280 1083.540 ;
        RECT 1061.320 1083.280 1061.580 1083.540 ;
        RECT 1055.340 20.440 1055.600 20.700 ;
        RECT 1059.020 20.440 1059.280 20.700 ;
      LAYER met2 ;
        RECT 1212.110 1100.580 1212.390 1104.000 ;
        RECT 1212.110 1100.000 1212.400 1100.580 ;
        RECT 1212.260 1088.330 1212.400 1100.000 ;
        RECT 1061.320 1088.010 1061.580 1088.330 ;
        RECT 1212.200 1088.010 1212.460 1088.330 ;
        RECT 1061.380 1083.570 1061.520 1088.010 ;
        RECT 1059.020 1083.250 1059.280 1083.570 ;
        RECT 1061.320 1083.250 1061.580 1083.570 ;
        RECT 1059.080 20.730 1059.220 1083.250 ;
        RECT 1055.340 20.410 1055.600 20.730 ;
        RECT 1059.020 20.410 1059.280 20.730 ;
        RECT 1055.400 2.000 1055.540 20.410 ;
        RECT 1055.190 -4.000 1055.750 2.000 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1076.010 1089.600 1076.330 1089.660 ;
        RECT 1218.150 1089.600 1218.470 1089.660 ;
        RECT 1076.010 1089.460 1218.470 1089.600 ;
        RECT 1076.010 1089.400 1076.330 1089.460 ;
        RECT 1218.150 1089.400 1218.470 1089.460 ;
        RECT 1073.250 20.640 1073.570 20.700 ;
        RECT 1076.010 20.640 1076.330 20.700 ;
        RECT 1073.250 20.500 1076.330 20.640 ;
        RECT 1073.250 20.440 1073.570 20.500 ;
        RECT 1076.010 20.440 1076.330 20.500 ;
      LAYER via ;
        RECT 1076.040 1089.400 1076.300 1089.660 ;
        RECT 1218.180 1089.400 1218.440 1089.660 ;
        RECT 1073.280 20.440 1073.540 20.700 ;
        RECT 1076.040 20.440 1076.300 20.700 ;
      LAYER met2 ;
        RECT 1218.090 1100.580 1218.370 1104.000 ;
        RECT 1218.090 1100.000 1218.380 1100.580 ;
        RECT 1218.240 1089.690 1218.380 1100.000 ;
        RECT 1076.040 1089.370 1076.300 1089.690 ;
        RECT 1218.180 1089.370 1218.440 1089.690 ;
        RECT 1076.100 20.730 1076.240 1089.370 ;
        RECT 1073.280 20.410 1073.540 20.730 ;
        RECT 1076.040 20.410 1076.300 20.730 ;
        RECT 1073.340 2.000 1073.480 20.410 ;
        RECT 1073.130 -4.000 1073.690 2.000 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1196.990 1083.480 1197.310 1083.540 ;
        RECT 1224.130 1083.480 1224.450 1083.540 ;
        RECT 1196.990 1083.340 1224.450 1083.480 ;
        RECT 1196.990 1083.280 1197.310 1083.340 ;
        RECT 1224.130 1083.280 1224.450 1083.340 ;
        RECT 1196.990 16.560 1197.310 16.620 ;
        RECT 1124.860 16.420 1197.310 16.560 ;
        RECT 1090.730 15.880 1091.050 15.940 ;
        RECT 1124.860 15.880 1125.000 16.420 ;
        RECT 1196.990 16.360 1197.310 16.420 ;
        RECT 1090.730 15.740 1125.000 15.880 ;
        RECT 1090.730 15.680 1091.050 15.740 ;
      LAYER via ;
        RECT 1197.020 1083.280 1197.280 1083.540 ;
        RECT 1224.160 1083.280 1224.420 1083.540 ;
        RECT 1090.760 15.680 1091.020 15.940 ;
        RECT 1197.020 16.360 1197.280 16.620 ;
      LAYER met2 ;
        RECT 1224.070 1100.580 1224.350 1104.000 ;
        RECT 1224.070 1100.000 1224.360 1100.580 ;
        RECT 1224.220 1083.570 1224.360 1100.000 ;
        RECT 1197.020 1083.250 1197.280 1083.570 ;
        RECT 1224.160 1083.250 1224.420 1083.570 ;
        RECT 1197.080 16.650 1197.220 1083.250 ;
        RECT 1197.020 16.330 1197.280 16.650 ;
        RECT 1090.760 15.650 1091.020 15.970 ;
        RECT 1090.820 2.000 1090.960 15.650 ;
        RECT 1090.610 -4.000 1091.170 2.000 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1225.050 1083.480 1225.370 1083.540 ;
        RECT 1230.570 1083.480 1230.890 1083.540 ;
        RECT 1225.050 1083.340 1230.890 1083.480 ;
        RECT 1225.050 1083.280 1225.370 1083.340 ;
        RECT 1230.570 1083.280 1230.890 1083.340 ;
        RECT 1108.670 20.640 1108.990 20.700 ;
        RECT 1225.050 20.640 1225.370 20.700 ;
        RECT 1108.670 20.500 1225.370 20.640 ;
        RECT 1108.670 20.440 1108.990 20.500 ;
        RECT 1225.050 20.440 1225.370 20.500 ;
      LAYER via ;
        RECT 1225.080 1083.280 1225.340 1083.540 ;
        RECT 1230.600 1083.280 1230.860 1083.540 ;
        RECT 1108.700 20.440 1108.960 20.700 ;
        RECT 1225.080 20.440 1225.340 20.700 ;
      LAYER met2 ;
        RECT 1230.510 1100.580 1230.790 1104.000 ;
        RECT 1230.510 1100.000 1230.800 1100.580 ;
        RECT 1230.660 1083.570 1230.800 1100.000 ;
        RECT 1225.080 1083.250 1225.340 1083.570 ;
        RECT 1230.600 1083.250 1230.860 1083.570 ;
        RECT 1225.140 20.730 1225.280 1083.250 ;
        RECT 1108.700 20.410 1108.960 20.730 ;
        RECT 1225.080 20.410 1225.340 20.730 ;
        RECT 1108.760 2.000 1108.900 20.410 ;
        RECT 1108.550 -4.000 1109.110 2.000 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1131.210 1085.860 1131.530 1085.920 ;
        RECT 1236.550 1085.860 1236.870 1085.920 ;
        RECT 1131.210 1085.720 1236.870 1085.860 ;
        RECT 1131.210 1085.660 1131.530 1085.720 ;
        RECT 1236.550 1085.660 1236.870 1085.720 ;
        RECT 1126.610 19.620 1126.930 19.680 ;
        RECT 1131.210 19.620 1131.530 19.680 ;
        RECT 1126.610 19.480 1131.530 19.620 ;
        RECT 1126.610 19.420 1126.930 19.480 ;
        RECT 1131.210 19.420 1131.530 19.480 ;
      LAYER via ;
        RECT 1131.240 1085.660 1131.500 1085.920 ;
        RECT 1236.580 1085.660 1236.840 1085.920 ;
        RECT 1126.640 19.420 1126.900 19.680 ;
        RECT 1131.240 19.420 1131.500 19.680 ;
      LAYER met2 ;
        RECT 1236.490 1100.580 1236.770 1104.000 ;
        RECT 1236.490 1100.000 1236.780 1100.580 ;
        RECT 1236.640 1085.950 1236.780 1100.000 ;
        RECT 1131.240 1085.630 1131.500 1085.950 ;
        RECT 1236.580 1085.630 1236.840 1085.950 ;
        RECT 1131.300 19.710 1131.440 1085.630 ;
        RECT 1126.640 19.390 1126.900 19.710 ;
        RECT 1131.240 19.390 1131.500 19.710 ;
        RECT 1126.700 2.000 1126.840 19.390 ;
        RECT 1126.490 -4.000 1127.050 2.000 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1238.390 1083.480 1238.710 1083.540 ;
        RECT 1242.530 1083.480 1242.850 1083.540 ;
        RECT 1238.390 1083.340 1242.850 1083.480 ;
        RECT 1238.390 1083.280 1238.710 1083.340 ;
        RECT 1242.530 1083.280 1242.850 1083.340 ;
        RECT 1144.550 15.880 1144.870 15.940 ;
        RECT 1238.390 15.880 1238.710 15.940 ;
        RECT 1144.550 15.740 1238.710 15.880 ;
        RECT 1144.550 15.680 1144.870 15.740 ;
        RECT 1238.390 15.680 1238.710 15.740 ;
      LAYER via ;
        RECT 1238.420 1083.280 1238.680 1083.540 ;
        RECT 1242.560 1083.280 1242.820 1083.540 ;
        RECT 1144.580 15.680 1144.840 15.940 ;
        RECT 1238.420 15.680 1238.680 15.940 ;
      LAYER met2 ;
        RECT 1242.470 1100.580 1242.750 1104.000 ;
        RECT 1242.470 1100.000 1242.760 1100.580 ;
        RECT 1242.620 1083.570 1242.760 1100.000 ;
        RECT 1238.420 1083.250 1238.680 1083.570 ;
        RECT 1242.560 1083.250 1242.820 1083.570 ;
        RECT 1238.480 15.970 1238.620 1083.250 ;
        RECT 1144.580 15.650 1144.840 15.970 ;
        RECT 1238.420 15.650 1238.680 15.970 ;
        RECT 1144.640 2.000 1144.780 15.650 ;
        RECT 1144.430 -4.000 1144.990 2.000 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1245.750 1083.480 1246.070 1083.540 ;
        RECT 1248.970 1083.480 1249.290 1083.540 ;
        RECT 1245.750 1083.340 1249.290 1083.480 ;
        RECT 1245.750 1083.280 1246.070 1083.340 ;
        RECT 1248.970 1083.280 1249.290 1083.340 ;
        RECT 1162.490 17.240 1162.810 17.300 ;
        RECT 1245.290 17.240 1245.610 17.300 ;
        RECT 1162.490 17.100 1245.610 17.240 ;
        RECT 1162.490 17.040 1162.810 17.100 ;
        RECT 1245.290 17.040 1245.610 17.100 ;
      LAYER via ;
        RECT 1245.780 1083.280 1246.040 1083.540 ;
        RECT 1249.000 1083.280 1249.260 1083.540 ;
        RECT 1162.520 17.040 1162.780 17.300 ;
        RECT 1245.320 17.040 1245.580 17.300 ;
      LAYER met2 ;
        RECT 1248.910 1100.580 1249.190 1104.000 ;
        RECT 1248.910 1100.000 1249.200 1100.580 ;
        RECT 1249.060 1083.570 1249.200 1100.000 ;
        RECT 1245.780 1083.250 1246.040 1083.570 ;
        RECT 1249.000 1083.250 1249.260 1083.570 ;
        RECT 1245.840 1072.090 1245.980 1083.250 ;
        RECT 1245.380 1071.950 1245.980 1072.090 ;
        RECT 1245.380 17.330 1245.520 1071.950 ;
        RECT 1162.520 17.010 1162.780 17.330 ;
        RECT 1245.320 17.010 1245.580 17.330 ;
        RECT 1162.580 2.000 1162.720 17.010 ;
        RECT 1162.370 -4.000 1162.930 2.000 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 680.410 30.160 680.730 30.220 ;
        RECT 1083.830 30.160 1084.150 30.220 ;
        RECT 680.410 30.020 1084.150 30.160 ;
        RECT 680.410 29.960 680.730 30.020 ;
        RECT 1083.830 29.960 1084.150 30.020 ;
      LAYER via ;
        RECT 680.440 29.960 680.700 30.220 ;
        RECT 1083.860 29.960 1084.120 30.220 ;
      LAYER met2 ;
        RECT 1083.310 1100.650 1083.590 1104.000 ;
        RECT 1083.310 1100.510 1084.060 1100.650 ;
        RECT 1083.310 1100.000 1083.590 1100.510 ;
        RECT 1083.920 30.250 1084.060 1100.510 ;
        RECT 680.440 29.930 680.700 30.250 ;
        RECT 1083.860 29.930 1084.120 30.250 ;
        RECT 680.500 2.000 680.640 29.930 ;
        RECT 680.290 -4.000 680.850 2.000 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1179.970 17.580 1180.290 17.640 ;
        RECT 1249.890 17.580 1250.210 17.640 ;
        RECT 1179.970 17.440 1250.210 17.580 ;
        RECT 1179.970 17.380 1180.290 17.440 ;
        RECT 1249.890 17.380 1250.210 17.440 ;
      LAYER via ;
        RECT 1180.000 17.380 1180.260 17.640 ;
        RECT 1249.920 17.380 1250.180 17.640 ;
      LAYER met2 ;
        RECT 1254.890 1100.650 1255.170 1104.000 ;
        RECT 1253.660 1100.510 1255.170 1100.650 ;
        RECT 1253.660 1072.770 1253.800 1100.510 ;
        RECT 1254.890 1100.000 1255.170 1100.510 ;
        RECT 1249.980 1072.630 1253.800 1072.770 ;
        RECT 1249.980 17.670 1250.120 1072.630 ;
        RECT 1180.000 17.350 1180.260 17.670 ;
        RECT 1249.920 17.350 1250.180 17.670 ;
        RECT 1180.060 2.000 1180.200 17.350 ;
        RECT 1179.850 -4.000 1180.410 2.000 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1254.030 1083.820 1254.350 1083.880 ;
        RECT 1260.930 1083.820 1261.250 1083.880 ;
        RECT 1254.030 1083.680 1261.250 1083.820 ;
        RECT 1254.030 1083.620 1254.350 1083.680 ;
        RECT 1260.930 1083.620 1261.250 1083.680 ;
        RECT 1197.910 18.260 1198.230 18.320 ;
        RECT 1252.190 18.260 1252.510 18.320 ;
        RECT 1197.910 18.120 1252.510 18.260 ;
        RECT 1197.910 18.060 1198.230 18.120 ;
        RECT 1252.190 18.060 1252.510 18.120 ;
      LAYER via ;
        RECT 1254.060 1083.620 1254.320 1083.880 ;
        RECT 1260.960 1083.620 1261.220 1083.880 ;
        RECT 1197.940 18.060 1198.200 18.320 ;
        RECT 1252.220 18.060 1252.480 18.320 ;
      LAYER met2 ;
        RECT 1260.870 1100.580 1261.150 1104.000 ;
        RECT 1260.870 1100.000 1261.160 1100.580 ;
        RECT 1261.020 1083.910 1261.160 1100.000 ;
        RECT 1254.060 1083.590 1254.320 1083.910 ;
        RECT 1260.960 1083.590 1261.220 1083.910 ;
        RECT 1254.120 1072.090 1254.260 1083.590 ;
        RECT 1252.280 1071.950 1254.260 1072.090 ;
        RECT 1252.280 18.350 1252.420 1071.950 ;
        RECT 1197.940 18.030 1198.200 18.350 ;
        RECT 1252.220 18.030 1252.480 18.350 ;
        RECT 1198.000 2.000 1198.140 18.030 ;
        RECT 1197.790 -4.000 1198.350 2.000 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1259.090 1083.480 1259.410 1083.540 ;
        RECT 1267.370 1083.480 1267.690 1083.540 ;
        RECT 1259.090 1083.340 1267.690 1083.480 ;
        RECT 1259.090 1083.280 1259.410 1083.340 ;
        RECT 1267.370 1083.280 1267.690 1083.340 ;
        RECT 1215.850 18.600 1216.170 18.660 ;
        RECT 1259.090 18.600 1259.410 18.660 ;
        RECT 1215.850 18.460 1259.410 18.600 ;
        RECT 1215.850 18.400 1216.170 18.460 ;
        RECT 1259.090 18.400 1259.410 18.460 ;
      LAYER via ;
        RECT 1259.120 1083.280 1259.380 1083.540 ;
        RECT 1267.400 1083.280 1267.660 1083.540 ;
        RECT 1215.880 18.400 1216.140 18.660 ;
        RECT 1259.120 18.400 1259.380 18.660 ;
      LAYER met2 ;
        RECT 1267.310 1100.580 1267.590 1104.000 ;
        RECT 1267.310 1100.000 1267.600 1100.580 ;
        RECT 1267.460 1083.570 1267.600 1100.000 ;
        RECT 1259.120 1083.250 1259.380 1083.570 ;
        RECT 1267.400 1083.250 1267.660 1083.570 ;
        RECT 1259.180 18.690 1259.320 1083.250 ;
        RECT 1215.880 18.370 1216.140 18.690 ;
        RECT 1259.120 18.370 1259.380 18.690 ;
        RECT 1215.940 2.000 1216.080 18.370 ;
        RECT 1215.730 -4.000 1216.290 2.000 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1233.790 18.940 1234.110 19.000 ;
        RECT 1270.590 18.940 1270.910 19.000 ;
        RECT 1233.790 18.800 1270.910 18.940 ;
        RECT 1233.790 18.740 1234.110 18.800 ;
        RECT 1270.590 18.740 1270.910 18.800 ;
      LAYER via ;
        RECT 1233.820 18.740 1234.080 19.000 ;
        RECT 1270.620 18.740 1270.880 19.000 ;
      LAYER met2 ;
        RECT 1273.290 1100.650 1273.570 1104.000 ;
        RECT 1272.060 1100.510 1273.570 1100.650 ;
        RECT 1272.060 1076.170 1272.200 1100.510 ;
        RECT 1273.290 1100.000 1273.570 1100.510 ;
        RECT 1271.140 1076.030 1272.200 1076.170 ;
        RECT 1271.140 1028.570 1271.280 1076.030 ;
        RECT 1270.680 1028.430 1271.280 1028.570 ;
        RECT 1270.680 19.030 1270.820 1028.430 ;
        RECT 1233.820 18.710 1234.080 19.030 ;
        RECT 1270.620 18.710 1270.880 19.030 ;
        RECT 1233.880 2.000 1234.020 18.710 ;
        RECT 1233.670 -4.000 1234.230 2.000 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1251.730 16.560 1252.050 16.620 ;
        RECT 1277.950 16.560 1278.270 16.620 ;
        RECT 1251.730 16.420 1278.270 16.560 ;
        RECT 1251.730 16.360 1252.050 16.420 ;
        RECT 1277.950 16.360 1278.270 16.420 ;
      LAYER via ;
        RECT 1251.760 16.360 1252.020 16.620 ;
        RECT 1277.980 16.360 1278.240 16.620 ;
      LAYER met2 ;
        RECT 1279.270 1100.650 1279.550 1104.000 ;
        RECT 1278.040 1100.510 1279.550 1100.650 ;
        RECT 1278.040 16.650 1278.180 1100.510 ;
        RECT 1279.270 1100.000 1279.550 1100.510 ;
        RECT 1251.760 16.330 1252.020 16.650 ;
        RECT 1277.980 16.330 1278.240 16.650 ;
        RECT 1251.820 2.000 1251.960 16.330 ;
        RECT 1251.610 -4.000 1252.170 2.000 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1269.210 16.220 1269.530 16.280 ;
        RECT 1284.390 16.220 1284.710 16.280 ;
        RECT 1269.210 16.080 1284.710 16.220 ;
        RECT 1269.210 16.020 1269.530 16.080 ;
        RECT 1284.390 16.020 1284.710 16.080 ;
      LAYER via ;
        RECT 1269.240 16.020 1269.500 16.280 ;
        RECT 1284.420 16.020 1284.680 16.280 ;
      LAYER met2 ;
        RECT 1285.710 1100.650 1285.990 1104.000 ;
        RECT 1284.480 1100.510 1285.990 1100.650 ;
        RECT 1284.480 16.310 1284.620 1100.510 ;
        RECT 1285.710 1100.000 1285.990 1100.510 ;
        RECT 1269.240 15.990 1269.500 16.310 ;
        RECT 1284.420 15.990 1284.680 16.310 ;
        RECT 1269.300 2.000 1269.440 15.990 ;
        RECT 1269.090 -4.000 1269.650 2.000 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1287.150 20.640 1287.470 20.700 ;
        RECT 1289.910 20.640 1290.230 20.700 ;
        RECT 1287.150 20.500 1290.230 20.640 ;
        RECT 1287.150 20.440 1287.470 20.500 ;
        RECT 1289.910 20.440 1290.230 20.500 ;
      LAYER via ;
        RECT 1287.180 20.440 1287.440 20.700 ;
        RECT 1289.940 20.440 1290.200 20.700 ;
      LAYER met2 ;
        RECT 1291.690 1100.650 1291.970 1104.000 ;
        RECT 1290.460 1100.510 1291.970 1100.650 ;
        RECT 1290.460 1088.410 1290.600 1100.510 ;
        RECT 1291.690 1100.000 1291.970 1100.510 ;
        RECT 1290.000 1088.270 1290.600 1088.410 ;
        RECT 1290.000 20.730 1290.140 1088.270 ;
        RECT 1287.180 20.410 1287.440 20.730 ;
        RECT 1289.940 20.410 1290.200 20.730 ;
        RECT 1287.240 2.000 1287.380 20.410 ;
        RECT 1287.030 -4.000 1287.590 2.000 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1305.625 766.105 1305.795 814.215 ;
        RECT 1305.625 669.545 1305.795 717.655 ;
        RECT 1305.625 572.645 1305.795 620.755 ;
        RECT 1305.625 476.085 1305.795 524.195 ;
        RECT 1304.705 379.525 1304.875 427.635 ;
        RECT 1305.625 89.845 1305.795 137.955 ;
      LAYER mcon ;
        RECT 1305.625 814.045 1305.795 814.215 ;
        RECT 1305.625 717.485 1305.795 717.655 ;
        RECT 1305.625 620.585 1305.795 620.755 ;
        RECT 1305.625 524.025 1305.795 524.195 ;
        RECT 1304.705 427.465 1304.875 427.635 ;
        RECT 1305.625 137.785 1305.795 137.955 ;
      LAYER met1 ;
        RECT 1297.730 1055.940 1298.050 1056.000 ;
        RECT 1305.550 1055.940 1305.870 1056.000 ;
        RECT 1297.730 1055.800 1305.870 1055.940 ;
        RECT 1297.730 1055.740 1298.050 1055.800 ;
        RECT 1305.550 1055.740 1305.870 1055.800 ;
        RECT 1305.550 910.760 1305.870 910.820 ;
        RECT 1306.470 910.760 1306.790 910.820 ;
        RECT 1305.550 910.620 1306.790 910.760 ;
        RECT 1305.550 910.560 1305.870 910.620 ;
        RECT 1306.470 910.560 1306.790 910.620 ;
        RECT 1305.550 814.200 1305.870 814.260 ;
        RECT 1305.355 814.060 1305.870 814.200 ;
        RECT 1305.550 814.000 1305.870 814.060 ;
        RECT 1305.550 766.260 1305.870 766.320 ;
        RECT 1305.355 766.120 1305.870 766.260 ;
        RECT 1305.550 766.060 1305.870 766.120 ;
        RECT 1305.550 717.640 1305.870 717.700 ;
        RECT 1305.355 717.500 1305.870 717.640 ;
        RECT 1305.550 717.440 1305.870 717.500 ;
        RECT 1305.550 669.700 1305.870 669.760 ;
        RECT 1305.355 669.560 1305.870 669.700 ;
        RECT 1305.550 669.500 1305.870 669.560 ;
        RECT 1305.550 620.740 1305.870 620.800 ;
        RECT 1305.355 620.600 1305.870 620.740 ;
        RECT 1305.550 620.540 1305.870 620.600 ;
        RECT 1305.550 572.800 1305.870 572.860 ;
        RECT 1305.355 572.660 1305.870 572.800 ;
        RECT 1305.550 572.600 1305.870 572.660 ;
        RECT 1305.550 524.180 1305.870 524.240 ;
        RECT 1305.355 524.040 1305.870 524.180 ;
        RECT 1305.550 523.980 1305.870 524.040 ;
        RECT 1305.550 476.240 1305.870 476.300 ;
        RECT 1305.355 476.100 1305.870 476.240 ;
        RECT 1305.550 476.040 1305.870 476.100 ;
        RECT 1304.645 427.620 1304.935 427.665 ;
        RECT 1305.550 427.620 1305.870 427.680 ;
        RECT 1304.645 427.480 1305.870 427.620 ;
        RECT 1304.645 427.435 1304.935 427.480 ;
        RECT 1305.550 427.420 1305.870 427.480 ;
        RECT 1304.630 379.680 1304.950 379.740 ;
        RECT 1304.435 379.540 1304.950 379.680 ;
        RECT 1304.630 379.480 1304.950 379.540 ;
        RECT 1305.090 289.580 1305.410 289.640 ;
        RECT 1305.550 289.580 1305.870 289.640 ;
        RECT 1305.090 289.440 1305.870 289.580 ;
        RECT 1305.090 289.380 1305.410 289.440 ;
        RECT 1305.550 289.380 1305.870 289.440 ;
        RECT 1305.090 282.580 1305.410 282.840 ;
        RECT 1305.180 282.440 1305.320 282.580 ;
        RECT 1306.010 282.440 1306.330 282.500 ;
        RECT 1305.180 282.300 1306.330 282.440 ;
        RECT 1306.010 282.240 1306.330 282.300 ;
        RECT 1306.010 234.500 1306.330 234.560 ;
        RECT 1306.470 234.500 1306.790 234.560 ;
        RECT 1306.010 234.360 1306.790 234.500 ;
        RECT 1306.010 234.300 1306.330 234.360 ;
        RECT 1306.470 234.300 1306.790 234.360 ;
        RECT 1305.550 145.080 1305.870 145.140 ;
        RECT 1306.010 145.080 1306.330 145.140 ;
        RECT 1305.550 144.940 1306.330 145.080 ;
        RECT 1305.550 144.880 1305.870 144.940 ;
        RECT 1306.010 144.880 1306.330 144.940 ;
        RECT 1305.550 137.940 1305.870 138.000 ;
        RECT 1305.355 137.800 1305.870 137.940 ;
        RECT 1305.550 137.740 1305.870 137.800 ;
        RECT 1305.550 90.000 1305.870 90.060 ;
        RECT 1305.355 89.860 1305.870 90.000 ;
        RECT 1305.550 89.800 1305.870 89.860 ;
      LAYER via ;
        RECT 1297.760 1055.740 1298.020 1056.000 ;
        RECT 1305.580 1055.740 1305.840 1056.000 ;
        RECT 1305.580 910.560 1305.840 910.820 ;
        RECT 1306.500 910.560 1306.760 910.820 ;
        RECT 1305.580 814.000 1305.840 814.260 ;
        RECT 1305.580 766.060 1305.840 766.320 ;
        RECT 1305.580 717.440 1305.840 717.700 ;
        RECT 1305.580 669.500 1305.840 669.760 ;
        RECT 1305.580 620.540 1305.840 620.800 ;
        RECT 1305.580 572.600 1305.840 572.860 ;
        RECT 1305.580 523.980 1305.840 524.240 ;
        RECT 1305.580 476.040 1305.840 476.300 ;
        RECT 1305.580 427.420 1305.840 427.680 ;
        RECT 1304.660 379.480 1304.920 379.740 ;
        RECT 1305.120 289.380 1305.380 289.640 ;
        RECT 1305.580 289.380 1305.840 289.640 ;
        RECT 1305.120 282.580 1305.380 282.840 ;
        RECT 1306.040 282.240 1306.300 282.500 ;
        RECT 1306.040 234.300 1306.300 234.560 ;
        RECT 1306.500 234.300 1306.760 234.560 ;
        RECT 1305.580 144.880 1305.840 145.140 ;
        RECT 1306.040 144.880 1306.300 145.140 ;
        RECT 1305.580 137.740 1305.840 138.000 ;
        RECT 1305.580 89.800 1305.840 90.060 ;
      LAYER met2 ;
        RECT 1297.670 1100.580 1297.950 1104.000 ;
        RECT 1297.670 1100.000 1297.960 1100.580 ;
        RECT 1297.820 1056.030 1297.960 1100.000 ;
        RECT 1297.760 1055.710 1298.020 1056.030 ;
        RECT 1305.580 1055.710 1305.840 1056.030 ;
        RECT 1305.640 910.850 1305.780 1055.710 ;
        RECT 1305.580 910.530 1305.840 910.850 ;
        RECT 1306.500 910.530 1306.760 910.850 ;
        RECT 1306.560 862.765 1306.700 910.530 ;
        RECT 1305.570 862.395 1305.850 862.765 ;
        RECT 1306.490 862.395 1306.770 862.765 ;
        RECT 1305.640 814.290 1305.780 862.395 ;
        RECT 1305.580 813.970 1305.840 814.290 ;
        RECT 1305.580 766.030 1305.840 766.350 ;
        RECT 1305.640 717.730 1305.780 766.030 ;
        RECT 1305.580 717.410 1305.840 717.730 ;
        RECT 1305.580 669.470 1305.840 669.790 ;
        RECT 1305.640 620.830 1305.780 669.470 ;
        RECT 1305.580 620.510 1305.840 620.830 ;
        RECT 1305.580 572.570 1305.840 572.890 ;
        RECT 1305.640 524.270 1305.780 572.570 ;
        RECT 1305.580 523.950 1305.840 524.270 ;
        RECT 1305.580 476.010 1305.840 476.330 ;
        RECT 1305.640 427.710 1305.780 476.010 ;
        RECT 1305.580 427.390 1305.840 427.710 ;
        RECT 1304.660 379.450 1304.920 379.770 ;
        RECT 1304.720 338.485 1304.860 379.450 ;
        RECT 1304.650 338.115 1304.930 338.485 ;
        RECT 1305.570 338.115 1305.850 338.485 ;
        RECT 1305.640 289.670 1305.780 338.115 ;
        RECT 1305.120 289.350 1305.380 289.670 ;
        RECT 1305.580 289.350 1305.840 289.670 ;
        RECT 1305.180 282.870 1305.320 289.350 ;
        RECT 1305.120 282.550 1305.380 282.870 ;
        RECT 1306.040 282.210 1306.300 282.530 ;
        RECT 1306.100 234.590 1306.240 282.210 ;
        RECT 1306.040 234.270 1306.300 234.590 ;
        RECT 1306.500 234.270 1306.760 234.590 ;
        RECT 1306.560 192.850 1306.700 234.270 ;
        RECT 1306.100 192.710 1306.700 192.850 ;
        RECT 1306.100 145.170 1306.240 192.710 ;
        RECT 1305.580 144.850 1305.840 145.170 ;
        RECT 1306.040 144.850 1306.300 145.170 ;
        RECT 1305.640 138.030 1305.780 144.850 ;
        RECT 1305.580 137.710 1305.840 138.030 ;
        RECT 1305.580 89.770 1305.840 90.090 ;
        RECT 1305.640 62.970 1305.780 89.770 ;
        RECT 1305.640 62.830 1306.240 62.970 ;
        RECT 1306.100 61.610 1306.240 62.830 ;
        RECT 1305.180 61.470 1306.240 61.610 ;
        RECT 1305.180 2.000 1305.320 61.470 ;
        RECT 1304.970 -4.000 1305.530 2.000 ;
      LAYER via2 ;
        RECT 1305.570 862.440 1305.850 862.720 ;
        RECT 1306.490 862.440 1306.770 862.720 ;
        RECT 1304.650 338.160 1304.930 338.440 ;
        RECT 1305.570 338.160 1305.850 338.440 ;
      LAYER met3 ;
        RECT 1305.545 862.730 1305.875 862.745 ;
        RECT 1306.465 862.730 1306.795 862.745 ;
        RECT 1305.545 862.430 1306.795 862.730 ;
        RECT 1305.545 862.415 1305.875 862.430 ;
        RECT 1306.465 862.415 1306.795 862.430 ;
        RECT 1304.625 338.450 1304.955 338.465 ;
        RECT 1305.545 338.450 1305.875 338.465 ;
        RECT 1304.625 338.150 1305.875 338.450 ;
        RECT 1304.625 338.135 1304.955 338.150 ;
        RECT 1305.545 338.135 1305.875 338.150 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1303.710 1088.240 1304.030 1088.300 ;
        RECT 1307.850 1088.240 1308.170 1088.300 ;
        RECT 1303.710 1088.100 1308.170 1088.240 ;
        RECT 1303.710 1088.040 1304.030 1088.100 ;
        RECT 1307.850 1088.040 1308.170 1088.100 ;
        RECT 1323.030 20.640 1323.350 20.700 ;
        RECT 1312.080 20.500 1323.350 20.640 ;
        RECT 1307.850 20.300 1308.170 20.360 ;
        RECT 1312.080 20.300 1312.220 20.500 ;
        RECT 1323.030 20.440 1323.350 20.500 ;
        RECT 1307.850 20.160 1312.220 20.300 ;
        RECT 1307.850 20.100 1308.170 20.160 ;
      LAYER via ;
        RECT 1303.740 1088.040 1304.000 1088.300 ;
        RECT 1307.880 1088.040 1308.140 1088.300 ;
        RECT 1307.880 20.100 1308.140 20.360 ;
        RECT 1323.060 20.440 1323.320 20.700 ;
      LAYER met2 ;
        RECT 1303.650 1100.580 1303.930 1104.000 ;
        RECT 1303.650 1100.000 1303.940 1100.580 ;
        RECT 1303.800 1088.330 1303.940 1100.000 ;
        RECT 1303.740 1088.010 1304.000 1088.330 ;
        RECT 1307.880 1088.010 1308.140 1088.330 ;
        RECT 1307.940 20.390 1308.080 1088.010 ;
        RECT 1323.060 20.410 1323.320 20.730 ;
        RECT 1307.880 20.070 1308.140 20.390 ;
        RECT 1323.120 2.000 1323.260 20.410 ;
        RECT 1322.910 -4.000 1323.470 2.000 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1310.610 18.600 1310.930 18.660 ;
        RECT 1340.510 18.600 1340.830 18.660 ;
        RECT 1310.610 18.460 1340.830 18.600 ;
        RECT 1310.610 18.400 1310.930 18.460 ;
        RECT 1340.510 18.400 1340.830 18.460 ;
      LAYER via ;
        RECT 1310.640 18.400 1310.900 18.660 ;
        RECT 1340.540 18.400 1340.800 18.660 ;
      LAYER met2 ;
        RECT 1310.090 1100.650 1310.370 1104.000 ;
        RECT 1310.090 1100.510 1310.840 1100.650 ;
        RECT 1310.090 1100.000 1310.370 1100.510 ;
        RECT 1310.700 18.690 1310.840 1100.510 ;
        RECT 1310.640 18.370 1310.900 18.690 ;
        RECT 1340.540 18.370 1340.800 18.690 ;
        RECT 1340.600 2.000 1340.740 18.370 ;
        RECT 1340.390 -4.000 1340.950 2.000 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1085.285 1007.505 1085.455 1055.615 ;
        RECT 1086.665 855.525 1086.835 903.975 ;
        RECT 1085.745 758.965 1085.915 807.075 ;
        RECT 1085.285 510.765 1085.455 558.535 ;
        RECT 1086.205 421.005 1086.375 476.935 ;
        RECT 1085.745 331.245 1085.915 379.015 ;
      LAYER mcon ;
        RECT 1085.285 1055.445 1085.455 1055.615 ;
        RECT 1086.665 903.805 1086.835 903.975 ;
        RECT 1085.745 806.905 1085.915 807.075 ;
        RECT 1085.285 558.365 1085.455 558.535 ;
        RECT 1086.205 476.765 1086.375 476.935 ;
        RECT 1085.745 378.845 1085.915 379.015 ;
      LAYER met1 ;
        RECT 1085.210 1055.600 1085.530 1055.660 ;
        RECT 1085.015 1055.460 1085.530 1055.600 ;
        RECT 1085.210 1055.400 1085.530 1055.460 ;
        RECT 1085.225 1007.660 1085.515 1007.705 ;
        RECT 1085.670 1007.660 1085.990 1007.720 ;
        RECT 1085.225 1007.520 1085.990 1007.660 ;
        RECT 1085.225 1007.475 1085.515 1007.520 ;
        RECT 1085.670 1007.460 1085.990 1007.520 ;
        RECT 1085.670 965.840 1085.990 965.900 ;
        RECT 1086.130 965.840 1086.450 965.900 ;
        RECT 1085.670 965.700 1086.450 965.840 ;
        RECT 1085.670 965.640 1085.990 965.700 ;
        RECT 1086.130 965.640 1086.450 965.700 ;
        RECT 1086.590 903.960 1086.910 904.020 ;
        RECT 1086.395 903.820 1086.910 903.960 ;
        RECT 1086.590 903.760 1086.910 903.820 ;
        RECT 1086.605 855.680 1086.895 855.725 ;
        RECT 1087.050 855.680 1087.370 855.740 ;
        RECT 1086.605 855.540 1087.370 855.680 ;
        RECT 1086.605 855.495 1086.895 855.540 ;
        RECT 1087.050 855.480 1087.370 855.540 ;
        RECT 1086.130 821.340 1086.450 821.400 ;
        RECT 1087.050 821.340 1087.370 821.400 ;
        RECT 1086.130 821.200 1087.370 821.340 ;
        RECT 1086.130 821.140 1086.450 821.200 ;
        RECT 1087.050 821.140 1087.370 821.200 ;
        RECT 1085.685 807.060 1085.975 807.105 ;
        RECT 1086.130 807.060 1086.450 807.120 ;
        RECT 1085.685 806.920 1086.450 807.060 ;
        RECT 1085.685 806.875 1085.975 806.920 ;
        RECT 1086.130 806.860 1086.450 806.920 ;
        RECT 1085.670 759.120 1085.990 759.180 ;
        RECT 1085.475 758.980 1085.990 759.120 ;
        RECT 1085.670 758.920 1085.990 758.980 ;
        RECT 1085.670 738.180 1085.990 738.440 ;
        RECT 1085.760 738.040 1085.900 738.180 ;
        RECT 1086.130 738.040 1086.450 738.100 ;
        RECT 1085.760 737.900 1086.450 738.040 ;
        RECT 1086.130 737.840 1086.450 737.900 ;
        RECT 1085.670 669.700 1085.990 669.760 ;
        RECT 1086.130 669.700 1086.450 669.760 ;
        RECT 1085.670 669.560 1086.450 669.700 ;
        RECT 1085.670 669.500 1085.990 669.560 ;
        RECT 1086.130 669.500 1086.450 669.560 ;
        RECT 1085.210 559.200 1085.530 559.260 ;
        RECT 1086.130 559.200 1086.450 559.260 ;
        RECT 1085.210 559.060 1086.450 559.200 ;
        RECT 1085.210 559.000 1085.530 559.060 ;
        RECT 1086.130 559.000 1086.450 559.060 ;
        RECT 1085.210 558.520 1085.530 558.580 ;
        RECT 1085.015 558.380 1085.530 558.520 ;
        RECT 1085.210 558.320 1085.530 558.380 ;
        RECT 1085.225 510.920 1085.515 510.965 ;
        RECT 1086.130 510.920 1086.450 510.980 ;
        RECT 1085.225 510.780 1086.450 510.920 ;
        RECT 1085.225 510.735 1085.515 510.780 ;
        RECT 1086.130 510.720 1086.450 510.780 ;
        RECT 1086.130 476.920 1086.450 476.980 ;
        RECT 1085.935 476.780 1086.450 476.920 ;
        RECT 1086.130 476.720 1086.450 476.780 ;
        RECT 1086.130 421.160 1086.450 421.220 ;
        RECT 1085.935 421.020 1086.450 421.160 ;
        RECT 1086.130 420.960 1086.450 421.020 ;
        RECT 1085.670 379.680 1085.990 379.740 ;
        RECT 1086.590 379.680 1086.910 379.740 ;
        RECT 1085.670 379.540 1086.910 379.680 ;
        RECT 1085.670 379.480 1085.990 379.540 ;
        RECT 1086.590 379.480 1086.910 379.540 ;
        RECT 1085.670 379.000 1085.990 379.060 ;
        RECT 1085.475 378.860 1085.990 379.000 ;
        RECT 1085.670 378.800 1085.990 378.860 ;
        RECT 1085.685 331.400 1085.975 331.445 ;
        RECT 1086.130 331.400 1086.450 331.460 ;
        RECT 1085.685 331.260 1086.450 331.400 ;
        RECT 1085.685 331.215 1085.975 331.260 ;
        RECT 1086.130 331.200 1086.450 331.260 ;
        RECT 1085.670 186.560 1085.990 186.620 ;
        RECT 1086.130 186.560 1086.450 186.620 ;
        RECT 1085.670 186.420 1086.450 186.560 ;
        RECT 1085.670 186.360 1085.990 186.420 ;
        RECT 1086.130 186.360 1086.450 186.420 ;
        RECT 1085.670 110.540 1085.990 110.800 ;
        RECT 1085.760 110.120 1085.900 110.540 ;
        RECT 1085.670 109.860 1085.990 110.120 ;
        RECT 698.350 29.820 698.670 29.880 ;
        RECT 1085.670 29.820 1085.990 29.880 ;
        RECT 698.350 29.680 1085.990 29.820 ;
        RECT 698.350 29.620 698.670 29.680 ;
        RECT 1085.670 29.620 1085.990 29.680 ;
      LAYER via ;
        RECT 1085.240 1055.400 1085.500 1055.660 ;
        RECT 1085.700 1007.460 1085.960 1007.720 ;
        RECT 1085.700 965.640 1085.960 965.900 ;
        RECT 1086.160 965.640 1086.420 965.900 ;
        RECT 1086.620 903.760 1086.880 904.020 ;
        RECT 1087.080 855.480 1087.340 855.740 ;
        RECT 1086.160 821.140 1086.420 821.400 ;
        RECT 1087.080 821.140 1087.340 821.400 ;
        RECT 1086.160 806.860 1086.420 807.120 ;
        RECT 1085.700 758.920 1085.960 759.180 ;
        RECT 1085.700 738.180 1085.960 738.440 ;
        RECT 1086.160 737.840 1086.420 738.100 ;
        RECT 1085.700 669.500 1085.960 669.760 ;
        RECT 1086.160 669.500 1086.420 669.760 ;
        RECT 1085.240 559.000 1085.500 559.260 ;
        RECT 1086.160 559.000 1086.420 559.260 ;
        RECT 1085.240 558.320 1085.500 558.580 ;
        RECT 1086.160 510.720 1086.420 510.980 ;
        RECT 1086.160 476.720 1086.420 476.980 ;
        RECT 1086.160 420.960 1086.420 421.220 ;
        RECT 1085.700 379.480 1085.960 379.740 ;
        RECT 1086.620 379.480 1086.880 379.740 ;
        RECT 1085.700 378.800 1085.960 379.060 ;
        RECT 1086.160 331.200 1086.420 331.460 ;
        RECT 1085.700 186.360 1085.960 186.620 ;
        RECT 1086.160 186.360 1086.420 186.620 ;
        RECT 1085.700 110.540 1085.960 110.800 ;
        RECT 1085.700 109.860 1085.960 110.120 ;
        RECT 698.380 29.620 698.640 29.880 ;
        RECT 1085.700 29.620 1085.960 29.880 ;
      LAYER met2 ;
        RECT 1089.750 1100.580 1090.030 1104.000 ;
        RECT 1089.750 1100.000 1090.040 1100.580 ;
        RECT 1089.900 1055.885 1090.040 1100.000 ;
        RECT 1085.230 1055.515 1085.510 1055.885 ;
        RECT 1089.830 1055.515 1090.110 1055.885 ;
        RECT 1085.240 1055.370 1085.500 1055.515 ;
        RECT 1085.700 1007.430 1085.960 1007.750 ;
        RECT 1085.760 965.930 1085.900 1007.430 ;
        RECT 1085.700 965.610 1085.960 965.930 ;
        RECT 1086.160 965.610 1086.420 965.930 ;
        RECT 1086.220 934.730 1086.360 965.610 ;
        RECT 1086.220 934.590 1087.280 934.730 ;
        RECT 1087.140 910.930 1087.280 934.590 ;
        RECT 1086.680 910.790 1087.280 910.930 ;
        RECT 1086.680 904.050 1086.820 910.790 ;
        RECT 1086.620 903.730 1086.880 904.050 ;
        RECT 1087.080 855.450 1087.340 855.770 ;
        RECT 1087.140 821.430 1087.280 855.450 ;
        RECT 1086.160 821.110 1086.420 821.430 ;
        RECT 1087.080 821.110 1087.340 821.430 ;
        RECT 1086.220 807.150 1086.360 821.110 ;
        RECT 1086.160 806.830 1086.420 807.150 ;
        RECT 1085.700 758.890 1085.960 759.210 ;
        RECT 1085.760 738.470 1085.900 758.890 ;
        RECT 1085.700 738.150 1085.960 738.470 ;
        RECT 1086.160 737.810 1086.420 738.130 ;
        RECT 1086.220 669.790 1086.360 737.810 ;
        RECT 1085.700 669.470 1085.960 669.790 ;
        RECT 1086.160 669.470 1086.420 669.790 ;
        RECT 1085.760 621.250 1085.900 669.470 ;
        RECT 1085.760 621.110 1086.360 621.250 ;
        RECT 1086.220 559.290 1086.360 621.110 ;
        RECT 1085.240 558.970 1085.500 559.290 ;
        RECT 1086.160 558.970 1086.420 559.290 ;
        RECT 1085.300 558.610 1085.440 558.970 ;
        RECT 1085.240 558.290 1085.500 558.610 ;
        RECT 1086.160 510.690 1086.420 511.010 ;
        RECT 1086.220 477.010 1086.360 510.690 ;
        RECT 1086.160 476.690 1086.420 477.010 ;
        RECT 1086.160 420.930 1086.420 421.250 ;
        RECT 1086.220 400.930 1086.360 420.930 ;
        RECT 1086.220 400.790 1086.820 400.930 ;
        RECT 1086.680 379.770 1086.820 400.790 ;
        RECT 1085.700 379.450 1085.960 379.770 ;
        RECT 1086.620 379.450 1086.880 379.770 ;
        RECT 1085.760 379.090 1085.900 379.450 ;
        RECT 1085.700 378.770 1085.960 379.090 ;
        RECT 1086.160 331.170 1086.420 331.490 ;
        RECT 1086.220 283.290 1086.360 331.170 ;
        RECT 1085.760 283.150 1086.360 283.290 ;
        RECT 1085.760 258.810 1085.900 283.150 ;
        RECT 1085.760 258.670 1086.360 258.810 ;
        RECT 1086.220 186.650 1086.360 258.670 ;
        RECT 1085.700 186.330 1085.960 186.650 ;
        RECT 1086.160 186.330 1086.420 186.650 ;
        RECT 1085.760 110.830 1085.900 186.330 ;
        RECT 1085.700 110.510 1085.960 110.830 ;
        RECT 1085.700 109.830 1085.960 110.150 ;
        RECT 1085.760 29.910 1085.900 109.830 ;
        RECT 698.380 29.590 698.640 29.910 ;
        RECT 1085.700 29.590 1085.960 29.910 ;
        RECT 698.440 2.000 698.580 29.590 ;
        RECT 698.230 -4.000 698.790 2.000 ;
      LAYER via2 ;
        RECT 1085.230 1055.560 1085.510 1055.840 ;
        RECT 1089.830 1055.560 1090.110 1055.840 ;
      LAYER met3 ;
        RECT 1085.205 1055.850 1085.535 1055.865 ;
        RECT 1089.805 1055.850 1090.135 1055.865 ;
        RECT 1085.205 1055.550 1090.135 1055.850 ;
        RECT 1085.205 1055.535 1085.535 1055.550 ;
        RECT 1089.805 1055.535 1090.135 1055.550 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1316.590 17.240 1316.910 17.300 ;
        RECT 1358.450 17.240 1358.770 17.300 ;
        RECT 1316.590 17.100 1358.770 17.240 ;
        RECT 1316.590 17.040 1316.910 17.100 ;
        RECT 1358.450 17.040 1358.770 17.100 ;
      LAYER via ;
        RECT 1316.620 17.040 1316.880 17.300 ;
        RECT 1358.480 17.040 1358.740 17.300 ;
      LAYER met2 ;
        RECT 1316.070 1100.650 1316.350 1104.000 ;
        RECT 1316.070 1100.510 1316.820 1100.650 ;
        RECT 1316.070 1100.000 1316.350 1100.510 ;
        RECT 1316.680 17.330 1316.820 1100.510 ;
        RECT 1316.620 17.010 1316.880 17.330 ;
        RECT 1358.480 17.010 1358.740 17.330 ;
        RECT 1358.540 2.000 1358.680 17.010 ;
        RECT 1358.330 -4.000 1358.890 2.000 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1322.110 1088.240 1322.430 1088.300 ;
        RECT 1362.590 1088.240 1362.910 1088.300 ;
        RECT 1322.110 1088.100 1362.910 1088.240 ;
        RECT 1322.110 1088.040 1322.430 1088.100 ;
        RECT 1362.590 1088.040 1362.910 1088.100 ;
        RECT 1362.590 17.580 1362.910 17.640 ;
        RECT 1376.390 17.580 1376.710 17.640 ;
        RECT 1362.590 17.440 1376.710 17.580 ;
        RECT 1362.590 17.380 1362.910 17.440 ;
        RECT 1376.390 17.380 1376.710 17.440 ;
      LAYER via ;
        RECT 1322.140 1088.040 1322.400 1088.300 ;
        RECT 1362.620 1088.040 1362.880 1088.300 ;
        RECT 1362.620 17.380 1362.880 17.640 ;
        RECT 1376.420 17.380 1376.680 17.640 ;
      LAYER met2 ;
        RECT 1322.050 1100.580 1322.330 1104.000 ;
        RECT 1322.050 1100.000 1322.340 1100.580 ;
        RECT 1322.200 1088.330 1322.340 1100.000 ;
        RECT 1322.140 1088.010 1322.400 1088.330 ;
        RECT 1362.620 1088.010 1362.880 1088.330 ;
        RECT 1362.680 17.670 1362.820 1088.010 ;
        RECT 1362.620 17.350 1362.880 17.670 ;
        RECT 1376.420 17.350 1376.680 17.670 ;
        RECT 1376.480 2.000 1376.620 17.350 ;
        RECT 1376.270 -4.000 1376.830 2.000 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1365.885 18.105 1366.055 19.295 ;
      LAYER mcon ;
        RECT 1365.885 19.125 1366.055 19.295 ;
      LAYER met1 ;
        RECT 1365.825 19.280 1366.115 19.325 ;
        RECT 1365.825 19.140 1371.560 19.280 ;
        RECT 1365.825 19.095 1366.115 19.140 ;
        RECT 1371.420 18.940 1371.560 19.140 ;
        RECT 1394.330 18.940 1394.650 19.000 ;
        RECT 1371.420 18.800 1394.650 18.940 ;
        RECT 1394.330 18.740 1394.650 18.800 ;
        RECT 1330.850 18.260 1331.170 18.320 ;
        RECT 1365.825 18.260 1366.115 18.305 ;
        RECT 1330.850 18.120 1366.115 18.260 ;
        RECT 1330.850 18.060 1331.170 18.120 ;
        RECT 1365.825 18.075 1366.115 18.120 ;
      LAYER via ;
        RECT 1394.360 18.740 1394.620 19.000 ;
        RECT 1330.880 18.060 1331.140 18.320 ;
      LAYER met2 ;
        RECT 1328.490 1100.650 1328.770 1104.000 ;
        RECT 1328.490 1100.510 1329.700 1100.650 ;
        RECT 1328.490 1100.000 1328.770 1100.510 ;
        RECT 1329.560 1088.410 1329.700 1100.510 ;
        RECT 1329.560 1088.270 1330.620 1088.410 ;
        RECT 1330.480 1076.170 1330.620 1088.270 ;
        RECT 1330.480 1076.030 1331.080 1076.170 ;
        RECT 1330.940 18.350 1331.080 1076.030 ;
        RECT 1394.360 18.710 1394.620 19.030 ;
        RECT 1330.880 18.030 1331.140 18.350 ;
        RECT 1394.420 2.000 1394.560 18.710 ;
        RECT 1394.210 -4.000 1394.770 2.000 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1379.225 1089.785 1379.855 1089.955 ;
      LAYER mcon ;
        RECT 1379.685 1089.785 1379.855 1089.955 ;
      LAYER met1 ;
        RECT 1334.530 1089.940 1334.850 1090.000 ;
        RECT 1379.165 1089.940 1379.455 1089.985 ;
        RECT 1334.530 1089.800 1379.455 1089.940 ;
        RECT 1334.530 1089.740 1334.850 1089.800 ;
        RECT 1379.165 1089.755 1379.455 1089.800 ;
        RECT 1379.625 1089.940 1379.915 1089.985 ;
        RECT 1397.090 1089.940 1397.410 1090.000 ;
        RECT 1379.625 1089.800 1397.410 1089.940 ;
        RECT 1379.625 1089.755 1379.915 1089.800 ;
        RECT 1397.090 1089.740 1397.410 1089.800 ;
        RECT 1397.090 20.640 1397.410 20.700 ;
        RECT 1412.270 20.640 1412.590 20.700 ;
        RECT 1397.090 20.500 1412.590 20.640 ;
        RECT 1397.090 20.440 1397.410 20.500 ;
        RECT 1412.270 20.440 1412.590 20.500 ;
      LAYER via ;
        RECT 1334.560 1089.740 1334.820 1090.000 ;
        RECT 1397.120 1089.740 1397.380 1090.000 ;
        RECT 1397.120 20.440 1397.380 20.700 ;
        RECT 1412.300 20.440 1412.560 20.700 ;
      LAYER met2 ;
        RECT 1334.470 1100.580 1334.750 1104.000 ;
        RECT 1334.470 1100.000 1334.760 1100.580 ;
        RECT 1334.620 1090.030 1334.760 1100.000 ;
        RECT 1334.560 1089.710 1334.820 1090.030 ;
        RECT 1397.120 1089.710 1397.380 1090.030 ;
        RECT 1397.180 20.730 1397.320 1089.710 ;
        RECT 1397.120 20.410 1397.380 20.730 ;
        RECT 1412.300 20.410 1412.560 20.730 ;
        RECT 1412.360 2.000 1412.500 20.410 ;
        RECT 1412.150 -4.000 1412.710 2.000 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1343.805 89.845 1343.975 137.955 ;
      LAYER mcon ;
        RECT 1343.805 137.785 1343.975 137.955 ;
      LAYER met1 ;
        RECT 1343.730 137.940 1344.050 138.000 ;
        RECT 1343.535 137.800 1344.050 137.940 ;
        RECT 1343.730 137.740 1344.050 137.800 ;
        RECT 1343.730 90.000 1344.050 90.060 ;
        RECT 1343.535 89.860 1344.050 90.000 ;
        RECT 1343.730 89.800 1344.050 89.860 ;
        RECT 1429.750 19.960 1430.070 20.020 ;
        RECT 1390.280 19.820 1430.070 19.960 ;
        RECT 1343.730 19.620 1344.050 19.680 ;
        RECT 1390.280 19.620 1390.420 19.820 ;
        RECT 1429.750 19.760 1430.070 19.820 ;
        RECT 1343.730 19.480 1390.420 19.620 ;
        RECT 1343.730 19.420 1344.050 19.480 ;
      LAYER via ;
        RECT 1343.760 137.740 1344.020 138.000 ;
        RECT 1343.760 89.800 1344.020 90.060 ;
        RECT 1343.760 19.420 1344.020 19.680 ;
        RECT 1429.780 19.760 1430.040 20.020 ;
      LAYER met2 ;
        RECT 1340.450 1100.650 1340.730 1104.000 ;
        RECT 1340.450 1100.510 1342.580 1100.650 ;
        RECT 1340.450 1100.000 1340.730 1100.510 ;
        RECT 1342.440 1076.170 1342.580 1100.510 ;
        RECT 1342.440 1076.030 1343.500 1076.170 ;
        RECT 1343.360 979.610 1343.500 1076.030 ;
        RECT 1343.360 979.470 1343.960 979.610 ;
        RECT 1343.820 835.450 1343.960 979.470 ;
        RECT 1343.360 835.310 1343.960 835.450 ;
        RECT 1343.360 834.770 1343.500 835.310 ;
        RECT 1343.360 834.630 1343.960 834.770 ;
        RECT 1343.820 738.890 1343.960 834.630 ;
        RECT 1343.360 738.750 1343.960 738.890 ;
        RECT 1343.360 738.210 1343.500 738.750 ;
        RECT 1343.360 738.070 1343.960 738.210 ;
        RECT 1343.820 642.330 1343.960 738.070 ;
        RECT 1343.360 642.190 1343.960 642.330 ;
        RECT 1343.360 641.650 1343.500 642.190 ;
        RECT 1343.360 641.510 1343.960 641.650 ;
        RECT 1343.820 545.770 1343.960 641.510 ;
        RECT 1343.360 545.630 1343.960 545.770 ;
        RECT 1343.360 545.090 1343.500 545.630 ;
        RECT 1343.360 544.950 1343.960 545.090 ;
        RECT 1343.820 449.210 1343.960 544.950 ;
        RECT 1343.360 449.070 1343.960 449.210 ;
        RECT 1343.360 448.530 1343.500 449.070 ;
        RECT 1343.360 448.390 1343.960 448.530 ;
        RECT 1343.820 351.970 1343.960 448.390 ;
        RECT 1343.360 351.830 1343.960 351.970 ;
        RECT 1343.360 351.290 1343.500 351.830 ;
        RECT 1343.360 351.150 1343.960 351.290 ;
        RECT 1343.820 255.410 1343.960 351.150 ;
        RECT 1343.360 255.270 1343.960 255.410 ;
        RECT 1343.360 254.730 1343.500 255.270 ;
        RECT 1343.360 254.590 1343.960 254.730 ;
        RECT 1343.820 146.045 1343.960 254.590 ;
        RECT 1343.750 145.675 1344.030 146.045 ;
        RECT 1343.750 144.995 1344.030 145.365 ;
        RECT 1343.820 138.030 1343.960 144.995 ;
        RECT 1343.760 137.710 1344.020 138.030 ;
        RECT 1343.760 89.770 1344.020 90.090 ;
        RECT 1343.820 19.710 1343.960 89.770 ;
        RECT 1429.780 19.730 1430.040 20.050 ;
        RECT 1343.760 19.390 1344.020 19.710 ;
        RECT 1429.840 2.000 1429.980 19.730 ;
        RECT 1429.630 -4.000 1430.190 2.000 ;
      LAYER via2 ;
        RECT 1343.750 145.720 1344.030 146.000 ;
        RECT 1343.750 145.040 1344.030 145.320 ;
      LAYER met3 ;
        RECT 1343.725 146.010 1344.055 146.025 ;
        RECT 1343.725 145.710 1344.730 146.010 ;
        RECT 1343.725 145.695 1344.055 145.710 ;
        RECT 1343.725 145.330 1344.055 145.345 ;
        RECT 1344.430 145.330 1344.730 145.710 ;
        RECT 1343.725 145.030 1344.730 145.330 ;
        RECT 1343.725 145.015 1344.055 145.030 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1346.950 1087.220 1347.270 1087.280 ;
        RECT 1351.090 1087.220 1351.410 1087.280 ;
        RECT 1346.950 1087.080 1351.410 1087.220 ;
        RECT 1346.950 1087.020 1347.270 1087.080 ;
        RECT 1351.090 1087.020 1351.410 1087.080 ;
        RECT 1351.090 14.860 1351.410 14.920 ;
        RECT 1447.690 14.860 1448.010 14.920 ;
        RECT 1351.090 14.720 1448.010 14.860 ;
        RECT 1351.090 14.660 1351.410 14.720 ;
        RECT 1447.690 14.660 1448.010 14.720 ;
      LAYER via ;
        RECT 1346.980 1087.020 1347.240 1087.280 ;
        RECT 1351.120 1087.020 1351.380 1087.280 ;
        RECT 1351.120 14.660 1351.380 14.920 ;
        RECT 1447.720 14.660 1447.980 14.920 ;
      LAYER met2 ;
        RECT 1346.890 1100.580 1347.170 1104.000 ;
        RECT 1346.890 1100.000 1347.180 1100.580 ;
        RECT 1347.040 1087.310 1347.180 1100.000 ;
        RECT 1346.980 1086.990 1347.240 1087.310 ;
        RECT 1351.120 1086.990 1351.380 1087.310 ;
        RECT 1351.180 14.950 1351.320 1086.990 ;
        RECT 1351.120 14.630 1351.380 14.950 ;
        RECT 1447.720 14.630 1447.980 14.950 ;
        RECT 1447.780 2.000 1447.920 14.630 ;
        RECT 1447.570 -4.000 1448.130 2.000 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1378.765 15.725 1378.935 17.595 ;
      LAYER mcon ;
        RECT 1378.765 17.425 1378.935 17.595 ;
      LAYER met1 ;
        RECT 1352.930 1088.580 1353.250 1088.640 ;
        RECT 1358.910 1088.580 1359.230 1088.640 ;
        RECT 1352.930 1088.440 1359.230 1088.580 ;
        RECT 1352.930 1088.380 1353.250 1088.440 ;
        RECT 1358.910 1088.380 1359.230 1088.440 ;
        RECT 1378.705 17.580 1378.995 17.625 ;
        RECT 1378.705 17.440 1383.980 17.580 ;
        RECT 1378.705 17.395 1378.995 17.440 ;
        RECT 1383.840 17.240 1383.980 17.440 ;
        RECT 1465.630 17.240 1465.950 17.300 ;
        RECT 1383.840 17.100 1465.950 17.240 ;
        RECT 1465.630 17.040 1465.950 17.100 ;
        RECT 1358.910 15.880 1359.230 15.940 ;
        RECT 1378.705 15.880 1378.995 15.925 ;
        RECT 1358.910 15.740 1378.995 15.880 ;
        RECT 1358.910 15.680 1359.230 15.740 ;
        RECT 1378.705 15.695 1378.995 15.740 ;
      LAYER via ;
        RECT 1352.960 1088.380 1353.220 1088.640 ;
        RECT 1358.940 1088.380 1359.200 1088.640 ;
        RECT 1465.660 17.040 1465.920 17.300 ;
        RECT 1358.940 15.680 1359.200 15.940 ;
      LAYER met2 ;
        RECT 1352.870 1100.580 1353.150 1104.000 ;
        RECT 1352.870 1100.000 1353.160 1100.580 ;
        RECT 1353.020 1088.670 1353.160 1100.000 ;
        RECT 1352.960 1088.350 1353.220 1088.670 ;
        RECT 1358.940 1088.350 1359.200 1088.670 ;
        RECT 1359.000 15.970 1359.140 1088.350 ;
        RECT 1465.660 17.010 1465.920 17.330 ;
        RECT 1358.940 15.650 1359.200 15.970 ;
        RECT 1465.720 2.000 1465.860 17.010 ;
        RECT 1465.510 -4.000 1466.070 2.000 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1415.565 1084.005 1415.735 1089.615 ;
        RECT 1459.725 1075.845 1459.895 1084.175 ;
        RECT 1459.725 724.965 1459.895 772.735 ;
        RECT 1459.725 572.645 1459.895 620.755 ;
        RECT 1459.265 48.365 1459.435 96.475 ;
      LAYER mcon ;
        RECT 1415.565 1089.445 1415.735 1089.615 ;
        RECT 1459.725 1084.005 1459.895 1084.175 ;
        RECT 1459.725 772.565 1459.895 772.735 ;
        RECT 1459.725 620.585 1459.895 620.755 ;
        RECT 1459.265 96.305 1459.435 96.475 ;
      LAYER met1 ;
        RECT 1358.910 1089.600 1359.230 1089.660 ;
        RECT 1415.505 1089.600 1415.795 1089.645 ;
        RECT 1358.910 1089.460 1415.795 1089.600 ;
        RECT 1358.910 1089.400 1359.230 1089.460 ;
        RECT 1415.505 1089.415 1415.795 1089.460 ;
        RECT 1415.505 1084.160 1415.795 1084.205 ;
        RECT 1459.665 1084.160 1459.955 1084.205 ;
        RECT 1415.505 1084.020 1459.955 1084.160 ;
        RECT 1415.505 1083.975 1415.795 1084.020 ;
        RECT 1459.665 1083.975 1459.955 1084.020 ;
        RECT 1459.650 1076.000 1459.970 1076.060 ;
        RECT 1459.455 1075.860 1459.970 1076.000 ;
        RECT 1459.650 1075.800 1459.970 1075.860 ;
        RECT 1458.270 917.900 1458.590 917.960 ;
        RECT 1459.650 917.900 1459.970 917.960 ;
        RECT 1458.270 917.760 1459.970 917.900 ;
        RECT 1458.270 917.700 1458.590 917.760 ;
        RECT 1459.650 917.700 1459.970 917.760 ;
        RECT 1459.650 883.700 1459.970 883.960 ;
        RECT 1459.740 882.940 1459.880 883.700 ;
        RECT 1459.650 882.680 1459.970 882.940 ;
        RECT 1459.650 786.460 1459.970 786.720 ;
        RECT 1459.740 786.040 1459.880 786.460 ;
        RECT 1459.650 785.780 1459.970 786.040 ;
        RECT 1459.650 772.720 1459.970 772.780 ;
        RECT 1459.455 772.580 1459.970 772.720 ;
        RECT 1459.650 772.520 1459.970 772.580 ;
        RECT 1459.650 725.120 1459.970 725.180 ;
        RECT 1459.455 724.980 1459.970 725.120 ;
        RECT 1459.650 724.920 1459.970 724.980 ;
        RECT 1459.190 717.640 1459.510 717.700 ;
        RECT 1459.650 717.640 1459.970 717.700 ;
        RECT 1459.190 717.500 1459.970 717.640 ;
        RECT 1459.190 717.440 1459.510 717.500 ;
        RECT 1459.650 717.440 1459.970 717.500 ;
        RECT 1458.730 669.360 1459.050 669.420 ;
        RECT 1459.650 669.360 1459.970 669.420 ;
        RECT 1458.730 669.220 1459.970 669.360 ;
        RECT 1458.730 669.160 1459.050 669.220 ;
        RECT 1459.650 669.160 1459.970 669.220 ;
        RECT 1459.650 620.740 1459.970 620.800 ;
        RECT 1459.455 620.600 1459.970 620.740 ;
        RECT 1459.650 620.540 1459.970 620.600 ;
        RECT 1459.650 572.800 1459.970 572.860 ;
        RECT 1459.455 572.660 1459.970 572.800 ;
        RECT 1459.650 572.600 1459.970 572.660 ;
        RECT 1459.650 483.380 1459.970 483.440 ;
        RECT 1460.110 483.380 1460.430 483.440 ;
        RECT 1459.650 483.240 1460.430 483.380 ;
        RECT 1459.650 483.180 1459.970 483.240 ;
        RECT 1460.110 483.180 1460.430 483.240 ;
        RECT 1459.650 400.420 1459.970 400.480 ;
        RECT 1459.280 400.280 1459.970 400.420 ;
        RECT 1459.280 400.140 1459.420 400.280 ;
        RECT 1459.650 400.220 1459.970 400.280 ;
        RECT 1459.190 399.880 1459.510 400.140 ;
        RECT 1459.650 331.060 1459.970 331.120 ;
        RECT 1459.650 330.920 1460.340 331.060 ;
        RECT 1459.650 330.860 1459.970 330.920 ;
        RECT 1460.200 330.780 1460.340 330.920 ;
        RECT 1460.110 330.520 1460.430 330.780 ;
        RECT 1459.190 255.240 1459.510 255.300 ;
        RECT 1460.110 255.240 1460.430 255.300 ;
        RECT 1459.190 255.100 1460.430 255.240 ;
        RECT 1459.190 255.040 1459.510 255.100 ;
        RECT 1460.110 255.040 1460.430 255.100 ;
        RECT 1458.730 240.960 1459.050 241.020 ;
        RECT 1459.190 240.960 1459.510 241.020 ;
        RECT 1458.730 240.820 1459.510 240.960 ;
        RECT 1458.730 240.760 1459.050 240.820 ;
        RECT 1459.190 240.760 1459.510 240.820 ;
        RECT 1459.190 158.820 1459.510 159.080 ;
        RECT 1459.280 158.680 1459.420 158.820 ;
        RECT 1459.650 158.680 1459.970 158.740 ;
        RECT 1459.280 158.540 1459.970 158.680 ;
        RECT 1459.650 158.480 1459.970 158.540 ;
        RECT 1459.650 110.540 1459.970 110.800 ;
        RECT 1459.740 110.120 1459.880 110.540 ;
        RECT 1459.650 109.860 1459.970 110.120 ;
        RECT 1459.205 96.460 1459.495 96.505 ;
        RECT 1459.650 96.460 1459.970 96.520 ;
        RECT 1459.205 96.320 1459.970 96.460 ;
        RECT 1459.205 96.275 1459.495 96.320 ;
        RECT 1459.650 96.260 1459.970 96.320 ;
        RECT 1459.190 48.520 1459.510 48.580 ;
        RECT 1458.995 48.380 1459.510 48.520 ;
        RECT 1459.190 48.320 1459.510 48.380 ;
        RECT 1459.190 4.660 1459.510 4.720 ;
        RECT 1483.570 4.660 1483.890 4.720 ;
        RECT 1459.190 4.520 1483.890 4.660 ;
        RECT 1459.190 4.460 1459.510 4.520 ;
        RECT 1483.570 4.460 1483.890 4.520 ;
      LAYER via ;
        RECT 1358.940 1089.400 1359.200 1089.660 ;
        RECT 1459.680 1075.800 1459.940 1076.060 ;
        RECT 1458.300 917.700 1458.560 917.960 ;
        RECT 1459.680 917.700 1459.940 917.960 ;
        RECT 1459.680 883.700 1459.940 883.960 ;
        RECT 1459.680 882.680 1459.940 882.940 ;
        RECT 1459.680 786.460 1459.940 786.720 ;
        RECT 1459.680 785.780 1459.940 786.040 ;
        RECT 1459.680 772.520 1459.940 772.780 ;
        RECT 1459.680 724.920 1459.940 725.180 ;
        RECT 1459.220 717.440 1459.480 717.700 ;
        RECT 1459.680 717.440 1459.940 717.700 ;
        RECT 1458.760 669.160 1459.020 669.420 ;
        RECT 1459.680 669.160 1459.940 669.420 ;
        RECT 1459.680 620.540 1459.940 620.800 ;
        RECT 1459.680 572.600 1459.940 572.860 ;
        RECT 1459.680 483.180 1459.940 483.440 ;
        RECT 1460.140 483.180 1460.400 483.440 ;
        RECT 1459.680 400.220 1459.940 400.480 ;
        RECT 1459.220 399.880 1459.480 400.140 ;
        RECT 1459.680 330.860 1459.940 331.120 ;
        RECT 1460.140 330.520 1460.400 330.780 ;
        RECT 1459.220 255.040 1459.480 255.300 ;
        RECT 1460.140 255.040 1460.400 255.300 ;
        RECT 1458.760 240.760 1459.020 241.020 ;
        RECT 1459.220 240.760 1459.480 241.020 ;
        RECT 1459.220 158.820 1459.480 159.080 ;
        RECT 1459.680 158.480 1459.940 158.740 ;
        RECT 1459.680 110.540 1459.940 110.800 ;
        RECT 1459.680 109.860 1459.940 110.120 ;
        RECT 1459.680 96.260 1459.940 96.520 ;
        RECT 1459.220 48.320 1459.480 48.580 ;
        RECT 1459.220 4.460 1459.480 4.720 ;
        RECT 1483.600 4.460 1483.860 4.720 ;
      LAYER met2 ;
        RECT 1358.850 1100.580 1359.130 1104.000 ;
        RECT 1358.850 1100.000 1359.140 1100.580 ;
        RECT 1359.000 1089.690 1359.140 1100.000 ;
        RECT 1358.940 1089.370 1359.200 1089.690 ;
        RECT 1459.680 1075.770 1459.940 1076.090 ;
        RECT 1459.740 980.290 1459.880 1075.770 ;
        RECT 1459.280 980.150 1459.880 980.290 ;
        RECT 1459.280 966.125 1459.420 980.150 ;
        RECT 1458.290 965.755 1458.570 966.125 ;
        RECT 1459.210 965.755 1459.490 966.125 ;
        RECT 1458.360 917.990 1458.500 965.755 ;
        RECT 1458.300 917.670 1458.560 917.990 ;
        RECT 1459.680 917.670 1459.940 917.990 ;
        RECT 1459.740 883.990 1459.880 917.670 ;
        RECT 1459.680 883.670 1459.940 883.990 ;
        RECT 1459.680 882.650 1459.940 882.970 ;
        RECT 1459.740 786.750 1459.880 882.650 ;
        RECT 1459.680 786.430 1459.940 786.750 ;
        RECT 1459.680 785.750 1459.940 786.070 ;
        RECT 1459.740 772.810 1459.880 785.750 ;
        RECT 1459.680 772.490 1459.940 772.810 ;
        RECT 1459.680 724.890 1459.940 725.210 ;
        RECT 1459.740 717.730 1459.880 724.890 ;
        RECT 1459.220 717.410 1459.480 717.730 ;
        RECT 1459.680 717.410 1459.940 717.730 ;
        RECT 1459.280 670.325 1459.420 717.410 ;
        RECT 1459.210 669.955 1459.490 670.325 ;
        RECT 1458.760 669.130 1459.020 669.450 ;
        RECT 1459.670 669.275 1459.950 669.645 ;
        RECT 1459.680 669.130 1459.940 669.275 ;
        RECT 1458.820 621.365 1458.960 669.130 ;
        RECT 1458.750 620.995 1459.030 621.365 ;
        RECT 1459.670 620.995 1459.950 621.365 ;
        RECT 1459.740 620.830 1459.880 620.995 ;
        RECT 1459.680 620.510 1459.940 620.830 ;
        RECT 1459.680 572.570 1459.940 572.890 ;
        RECT 1459.740 496.810 1459.880 572.570 ;
        RECT 1459.740 496.670 1460.340 496.810 ;
        RECT 1460.200 483.470 1460.340 496.670 ;
        RECT 1459.680 483.150 1459.940 483.470 ;
        RECT 1460.140 483.150 1460.400 483.470 ;
        RECT 1459.740 400.510 1459.880 483.150 ;
        RECT 1459.680 400.190 1459.940 400.510 ;
        RECT 1459.220 399.850 1459.480 400.170 ;
        RECT 1459.280 386.650 1459.420 399.850 ;
        RECT 1459.280 386.510 1459.880 386.650 ;
        RECT 1459.740 331.150 1459.880 386.510 ;
        RECT 1459.680 330.830 1459.940 331.150 ;
        RECT 1460.140 330.490 1460.400 330.810 ;
        RECT 1460.200 255.330 1460.340 330.490 ;
        RECT 1459.220 255.010 1459.480 255.330 ;
        RECT 1460.140 255.010 1460.400 255.330 ;
        RECT 1459.280 241.050 1459.420 255.010 ;
        RECT 1458.760 240.730 1459.020 241.050 ;
        RECT 1459.220 240.730 1459.480 241.050 ;
        RECT 1458.820 216.650 1458.960 240.730 ;
        RECT 1458.820 216.510 1459.420 216.650 ;
        RECT 1459.280 159.110 1459.420 216.510 ;
        RECT 1459.220 158.790 1459.480 159.110 ;
        RECT 1459.680 158.450 1459.940 158.770 ;
        RECT 1459.740 110.830 1459.880 158.450 ;
        RECT 1459.680 110.510 1459.940 110.830 ;
        RECT 1459.680 109.830 1459.940 110.150 ;
        RECT 1459.740 96.550 1459.880 109.830 ;
        RECT 1459.680 96.230 1459.940 96.550 ;
        RECT 1459.220 48.290 1459.480 48.610 ;
        RECT 1459.280 4.750 1459.420 48.290 ;
        RECT 1459.220 4.430 1459.480 4.750 ;
        RECT 1483.600 4.430 1483.860 4.750 ;
        RECT 1483.660 2.000 1483.800 4.430 ;
        RECT 1483.450 -4.000 1484.010 2.000 ;
      LAYER via2 ;
        RECT 1458.290 965.800 1458.570 966.080 ;
        RECT 1459.210 965.800 1459.490 966.080 ;
        RECT 1459.210 670.000 1459.490 670.280 ;
        RECT 1459.670 669.320 1459.950 669.600 ;
        RECT 1458.750 621.040 1459.030 621.320 ;
        RECT 1459.670 621.040 1459.950 621.320 ;
      LAYER met3 ;
        RECT 1458.265 966.090 1458.595 966.105 ;
        RECT 1459.185 966.090 1459.515 966.105 ;
        RECT 1458.265 965.790 1459.515 966.090 ;
        RECT 1458.265 965.775 1458.595 965.790 ;
        RECT 1459.185 965.775 1459.515 965.790 ;
        RECT 1459.185 670.290 1459.515 670.305 ;
        RECT 1459.185 669.975 1459.730 670.290 ;
        RECT 1459.430 669.625 1459.730 669.975 ;
        RECT 1459.430 669.310 1459.975 669.625 ;
        RECT 1459.645 669.295 1459.975 669.310 ;
        RECT 1458.725 621.330 1459.055 621.345 ;
        RECT 1459.645 621.330 1459.975 621.345 ;
        RECT 1458.725 621.030 1459.975 621.330 ;
        RECT 1458.725 621.015 1459.055 621.030 ;
        RECT 1459.645 621.015 1459.975 621.030 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1365.810 773.200 1366.130 773.460 ;
        RECT 1365.900 772.780 1366.040 773.200 ;
        RECT 1365.810 772.520 1366.130 772.780 ;
        RECT 1501.510 15.880 1501.830 15.940 ;
        RECT 1390.740 15.740 1501.830 15.880 ;
        RECT 1365.810 15.540 1366.130 15.600 ;
        RECT 1390.740 15.540 1390.880 15.740 ;
        RECT 1501.510 15.680 1501.830 15.740 ;
        RECT 1365.810 15.400 1390.880 15.540 ;
        RECT 1365.810 15.340 1366.130 15.400 ;
      LAYER via ;
        RECT 1365.840 773.200 1366.100 773.460 ;
        RECT 1365.840 772.520 1366.100 772.780 ;
        RECT 1365.840 15.340 1366.100 15.600 ;
        RECT 1501.540 15.680 1501.800 15.940 ;
      LAYER met2 ;
        RECT 1365.290 1100.650 1365.570 1104.000 ;
        RECT 1365.290 1100.510 1366.040 1100.650 ;
        RECT 1365.290 1100.000 1365.570 1100.510 ;
        RECT 1365.900 773.490 1366.040 1100.510 ;
        RECT 1365.840 773.170 1366.100 773.490 ;
        RECT 1365.840 772.490 1366.100 772.810 ;
        RECT 1365.900 15.630 1366.040 772.490 ;
        RECT 1501.540 15.650 1501.800 15.970 ;
        RECT 1365.840 15.310 1366.100 15.630 ;
        RECT 1501.600 2.000 1501.740 15.650 ;
        RECT 1501.390 -4.000 1501.950 2.000 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1389.345 14.875 1389.515 15.215 ;
        RECT 1390.265 15.045 1391.355 15.215 ;
        RECT 1401.765 15.045 1401.935 16.235 ;
        RECT 1390.265 14.875 1390.435 15.045 ;
        RECT 1389.345 14.705 1390.435 14.875 ;
        RECT 1485.945 14.705 1486.115 16.235 ;
      LAYER mcon ;
        RECT 1401.765 16.065 1401.935 16.235 ;
        RECT 1389.345 15.045 1389.515 15.215 ;
        RECT 1391.185 15.045 1391.355 15.215 ;
        RECT 1485.945 16.065 1486.115 16.235 ;
      LAYER met1 ;
        RECT 1401.705 16.220 1401.995 16.265 ;
        RECT 1485.885 16.220 1486.175 16.265 ;
        RECT 1401.705 16.080 1486.175 16.220 ;
        RECT 1401.705 16.035 1401.995 16.080 ;
        RECT 1485.885 16.035 1486.175 16.080 ;
        RECT 1372.710 15.200 1373.030 15.260 ;
        RECT 1389.285 15.200 1389.575 15.245 ;
        RECT 1372.710 15.060 1389.575 15.200 ;
        RECT 1372.710 15.000 1373.030 15.060 ;
        RECT 1389.285 15.015 1389.575 15.060 ;
        RECT 1391.125 15.200 1391.415 15.245 ;
        RECT 1401.705 15.200 1401.995 15.245 ;
        RECT 1391.125 15.060 1401.995 15.200 ;
        RECT 1391.125 15.015 1391.415 15.060 ;
        RECT 1401.705 15.015 1401.995 15.060 ;
        RECT 1485.885 14.860 1486.175 14.905 ;
        RECT 1518.990 14.860 1519.310 14.920 ;
        RECT 1485.885 14.720 1519.310 14.860 ;
        RECT 1485.885 14.675 1486.175 14.720 ;
        RECT 1518.990 14.660 1519.310 14.720 ;
      LAYER via ;
        RECT 1372.740 15.000 1373.000 15.260 ;
        RECT 1519.020 14.660 1519.280 14.920 ;
      LAYER met2 ;
        RECT 1371.270 1100.650 1371.550 1104.000 ;
        RECT 1371.270 1100.510 1372.940 1100.650 ;
        RECT 1371.270 1100.000 1371.550 1100.510 ;
        RECT 1372.800 15.290 1372.940 1100.510 ;
        RECT 1372.740 14.970 1373.000 15.290 ;
        RECT 1519.020 14.630 1519.280 14.950 ;
        RECT 1519.080 2.000 1519.220 14.630 ;
        RECT 1518.870 -4.000 1519.430 2.000 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1090.270 1052.200 1090.590 1052.260 ;
        RECT 1093.950 1052.200 1094.270 1052.260 ;
        RECT 1090.270 1052.060 1094.270 1052.200 ;
        RECT 1090.270 1052.000 1090.590 1052.060 ;
        RECT 1093.950 1052.000 1094.270 1052.060 ;
        RECT 716.290 29.480 716.610 29.540 ;
        RECT 1090.270 29.480 1090.590 29.540 ;
        RECT 716.290 29.340 1090.590 29.480 ;
        RECT 716.290 29.280 716.610 29.340 ;
        RECT 1090.270 29.280 1090.590 29.340 ;
      LAYER via ;
        RECT 1090.300 1052.000 1090.560 1052.260 ;
        RECT 1093.980 1052.000 1094.240 1052.260 ;
        RECT 716.320 29.280 716.580 29.540 ;
        RECT 1090.300 29.280 1090.560 29.540 ;
      LAYER met2 ;
        RECT 1095.730 1100.650 1096.010 1104.000 ;
        RECT 1094.040 1100.510 1096.010 1100.650 ;
        RECT 1094.040 1052.290 1094.180 1100.510 ;
        RECT 1095.730 1100.000 1096.010 1100.510 ;
        RECT 1090.300 1051.970 1090.560 1052.290 ;
        RECT 1093.980 1051.970 1094.240 1052.290 ;
        RECT 1090.360 29.570 1090.500 1051.970 ;
        RECT 716.320 29.250 716.580 29.570 ;
        RECT 1090.300 29.250 1090.560 29.570 ;
        RECT 716.380 2.000 716.520 29.250 ;
        RECT 716.170 -4.000 716.730 2.000 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1379.225 855.525 1379.395 903.975 ;
        RECT 1379.225 669.545 1379.395 717.655 ;
        RECT 1379.225 476.085 1379.395 524.195 ;
        RECT 1378.765 269.025 1378.935 317.475 ;
        RECT 1379.225 166.005 1379.395 193.035 ;
        RECT 1379.685 89.845 1379.855 137.955 ;
      LAYER mcon ;
        RECT 1379.225 903.805 1379.395 903.975 ;
        RECT 1379.225 717.485 1379.395 717.655 ;
        RECT 1379.225 524.025 1379.395 524.195 ;
        RECT 1378.765 317.305 1378.935 317.475 ;
        RECT 1379.225 192.865 1379.395 193.035 ;
        RECT 1379.685 137.785 1379.855 137.955 ;
      LAYER met1 ;
        RECT 1379.150 1048.800 1379.470 1048.860 ;
        RECT 1380.530 1048.800 1380.850 1048.860 ;
        RECT 1379.150 1048.660 1380.850 1048.800 ;
        RECT 1379.150 1048.600 1379.470 1048.660 ;
        RECT 1380.530 1048.600 1380.850 1048.660 ;
        RECT 1379.150 976.380 1379.470 976.440 ;
        RECT 1380.530 976.380 1380.850 976.440 ;
        RECT 1379.150 976.240 1380.850 976.380 ;
        RECT 1379.150 976.180 1379.470 976.240 ;
        RECT 1380.530 976.180 1380.850 976.240 ;
        RECT 1379.150 918.040 1379.470 918.300 ;
        RECT 1379.240 917.620 1379.380 918.040 ;
        RECT 1379.150 917.360 1379.470 917.620 ;
        RECT 1379.150 903.960 1379.470 904.020 ;
        RECT 1378.955 903.820 1379.470 903.960 ;
        RECT 1379.150 903.760 1379.470 903.820 ;
        RECT 1379.165 855.680 1379.455 855.725 ;
        RECT 1379.610 855.680 1379.930 855.740 ;
        RECT 1379.165 855.540 1379.930 855.680 ;
        RECT 1379.165 855.495 1379.455 855.540 ;
        RECT 1379.610 855.480 1379.930 855.540 ;
        RECT 1379.150 814.200 1379.470 814.260 ;
        RECT 1379.610 814.200 1379.930 814.260 ;
        RECT 1379.150 814.060 1379.930 814.200 ;
        RECT 1379.150 814.000 1379.470 814.060 ;
        RECT 1379.610 814.000 1379.930 814.060 ;
        RECT 1379.165 717.640 1379.455 717.685 ;
        RECT 1379.610 717.640 1379.930 717.700 ;
        RECT 1379.165 717.500 1379.930 717.640 ;
        RECT 1379.165 717.455 1379.455 717.500 ;
        RECT 1379.610 717.440 1379.930 717.500 ;
        RECT 1379.150 669.700 1379.470 669.760 ;
        RECT 1378.955 669.560 1379.470 669.700 ;
        RECT 1379.150 669.500 1379.470 669.560 ;
        RECT 1379.610 620.740 1379.930 620.800 ;
        RECT 1380.070 620.740 1380.390 620.800 ;
        RECT 1379.610 620.600 1380.390 620.740 ;
        RECT 1379.610 620.540 1379.930 620.600 ;
        RECT 1380.070 620.540 1380.390 620.600 ;
        RECT 1379.165 524.180 1379.455 524.225 ;
        RECT 1379.610 524.180 1379.930 524.240 ;
        RECT 1379.165 524.040 1379.930 524.180 ;
        RECT 1379.165 523.995 1379.455 524.040 ;
        RECT 1379.610 523.980 1379.930 524.040 ;
        RECT 1379.150 476.240 1379.470 476.300 ;
        RECT 1378.955 476.100 1379.470 476.240 ;
        RECT 1379.150 476.040 1379.470 476.100 ;
        RECT 1378.690 420.820 1379.010 420.880 ;
        RECT 1379.610 420.820 1379.930 420.880 ;
        RECT 1378.690 420.680 1379.930 420.820 ;
        RECT 1378.690 420.620 1379.010 420.680 ;
        RECT 1379.610 420.620 1379.930 420.680 ;
        RECT 1379.150 330.860 1379.470 331.120 ;
        RECT 1379.240 330.720 1379.380 330.860 ;
        RECT 1380.070 330.720 1380.390 330.780 ;
        RECT 1379.240 330.580 1380.390 330.720 ;
        RECT 1380.070 330.520 1380.390 330.580 ;
        RECT 1378.705 317.460 1378.995 317.505 ;
        RECT 1379.610 317.460 1379.930 317.520 ;
        RECT 1378.705 317.320 1379.930 317.460 ;
        RECT 1378.705 317.275 1378.995 317.320 ;
        RECT 1379.610 317.260 1379.930 317.320 ;
        RECT 1378.690 269.180 1379.010 269.240 ;
        RECT 1378.495 269.040 1379.010 269.180 ;
        RECT 1378.690 268.980 1379.010 269.040 ;
        RECT 1378.690 265.780 1379.010 265.840 ;
        RECT 1379.610 265.780 1379.930 265.840 ;
        RECT 1378.690 265.640 1379.930 265.780 ;
        RECT 1378.690 265.580 1379.010 265.640 ;
        RECT 1379.610 265.580 1379.930 265.640 ;
        RECT 1379.150 241.300 1379.470 241.360 ;
        RECT 1379.610 241.300 1379.930 241.360 ;
        RECT 1379.150 241.160 1379.930 241.300 ;
        RECT 1379.150 241.100 1379.470 241.160 ;
        RECT 1379.610 241.100 1379.930 241.160 ;
        RECT 1379.150 193.020 1379.470 193.080 ;
        RECT 1378.955 192.880 1379.470 193.020 ;
        RECT 1379.150 192.820 1379.470 192.880 ;
        RECT 1379.165 166.160 1379.455 166.205 ;
        RECT 1379.610 166.160 1379.930 166.220 ;
        RECT 1379.165 166.020 1379.930 166.160 ;
        RECT 1379.165 165.975 1379.455 166.020 ;
        RECT 1379.610 165.960 1379.930 166.020 ;
        RECT 1379.610 137.940 1379.930 138.000 ;
        RECT 1379.415 137.800 1379.930 137.940 ;
        RECT 1379.610 137.740 1379.930 137.800 ;
        RECT 1379.610 90.000 1379.930 90.060 ;
        RECT 1379.415 89.860 1379.930 90.000 ;
        RECT 1379.610 89.800 1379.930 89.860 ;
        RECT 1536.930 16.560 1537.250 16.620 ;
        RECT 1401.320 16.420 1537.250 16.560 ;
        RECT 1379.610 16.220 1379.930 16.280 ;
        RECT 1401.320 16.220 1401.460 16.420 ;
        RECT 1536.930 16.360 1537.250 16.420 ;
        RECT 1379.610 16.080 1401.460 16.220 ;
        RECT 1379.610 16.020 1379.930 16.080 ;
      LAYER via ;
        RECT 1379.180 1048.600 1379.440 1048.860 ;
        RECT 1380.560 1048.600 1380.820 1048.860 ;
        RECT 1379.180 976.180 1379.440 976.440 ;
        RECT 1380.560 976.180 1380.820 976.440 ;
        RECT 1379.180 918.040 1379.440 918.300 ;
        RECT 1379.180 917.360 1379.440 917.620 ;
        RECT 1379.180 903.760 1379.440 904.020 ;
        RECT 1379.640 855.480 1379.900 855.740 ;
        RECT 1379.180 814.000 1379.440 814.260 ;
        RECT 1379.640 814.000 1379.900 814.260 ;
        RECT 1379.640 717.440 1379.900 717.700 ;
        RECT 1379.180 669.500 1379.440 669.760 ;
        RECT 1379.640 620.540 1379.900 620.800 ;
        RECT 1380.100 620.540 1380.360 620.800 ;
        RECT 1379.640 523.980 1379.900 524.240 ;
        RECT 1379.180 476.040 1379.440 476.300 ;
        RECT 1378.720 420.620 1378.980 420.880 ;
        RECT 1379.640 420.620 1379.900 420.880 ;
        RECT 1379.180 330.860 1379.440 331.120 ;
        RECT 1380.100 330.520 1380.360 330.780 ;
        RECT 1379.640 317.260 1379.900 317.520 ;
        RECT 1378.720 268.980 1378.980 269.240 ;
        RECT 1378.720 265.580 1378.980 265.840 ;
        RECT 1379.640 265.580 1379.900 265.840 ;
        RECT 1379.180 241.100 1379.440 241.360 ;
        RECT 1379.640 241.100 1379.900 241.360 ;
        RECT 1379.180 192.820 1379.440 193.080 ;
        RECT 1379.640 165.960 1379.900 166.220 ;
        RECT 1379.640 137.740 1379.900 138.000 ;
        RECT 1379.640 89.800 1379.900 90.060 ;
        RECT 1379.640 16.020 1379.900 16.280 ;
        RECT 1536.960 16.360 1537.220 16.620 ;
      LAYER met2 ;
        RECT 1377.250 1100.580 1377.530 1104.000 ;
        RECT 1377.250 1100.000 1377.540 1100.580 ;
        RECT 1377.400 1098.045 1377.540 1100.000 ;
        RECT 1377.330 1097.675 1377.610 1098.045 ;
        RECT 1379.170 1096.995 1379.450 1097.365 ;
        RECT 1379.240 1048.890 1379.380 1096.995 ;
        RECT 1379.180 1048.570 1379.440 1048.890 ;
        RECT 1380.560 1048.570 1380.820 1048.890 ;
        RECT 1380.620 976.470 1380.760 1048.570 ;
        RECT 1379.180 976.150 1379.440 976.470 ;
        RECT 1380.560 976.150 1380.820 976.470 ;
        RECT 1379.240 918.330 1379.380 976.150 ;
        RECT 1379.180 918.010 1379.440 918.330 ;
        RECT 1379.180 917.330 1379.440 917.650 ;
        RECT 1379.240 904.050 1379.380 917.330 ;
        RECT 1379.180 903.730 1379.440 904.050 ;
        RECT 1379.640 855.450 1379.900 855.770 ;
        RECT 1379.700 814.290 1379.840 855.450 ;
        RECT 1379.180 813.970 1379.440 814.290 ;
        RECT 1379.640 813.970 1379.900 814.290 ;
        RECT 1379.240 724.610 1379.380 813.970 ;
        RECT 1379.240 724.470 1379.840 724.610 ;
        RECT 1379.700 717.730 1379.840 724.470 ;
        RECT 1379.640 717.410 1379.900 717.730 ;
        RECT 1379.180 669.470 1379.440 669.790 ;
        RECT 1379.240 651.850 1379.380 669.470 ;
        RECT 1379.240 651.710 1379.840 651.850 ;
        RECT 1379.700 620.830 1379.840 651.710 ;
        RECT 1379.640 620.510 1379.900 620.830 ;
        RECT 1380.100 620.510 1380.360 620.830 ;
        RECT 1380.160 554.610 1380.300 620.510 ;
        RECT 1379.700 554.470 1380.300 554.610 ;
        RECT 1379.700 524.270 1379.840 554.470 ;
        RECT 1379.640 523.950 1379.900 524.270 ;
        RECT 1379.180 476.010 1379.440 476.330 ;
        RECT 1379.240 448.360 1379.380 476.010 ;
        RECT 1379.240 448.220 1379.840 448.360 ;
        RECT 1379.700 420.910 1379.840 448.220 ;
        RECT 1378.720 420.590 1378.980 420.910 ;
        RECT 1379.640 420.590 1379.900 420.910 ;
        RECT 1378.780 373.050 1378.920 420.590 ;
        RECT 1378.780 372.910 1379.380 373.050 ;
        RECT 1379.240 331.150 1379.380 372.910 ;
        RECT 1379.180 330.830 1379.440 331.150 ;
        RECT 1380.100 330.490 1380.360 330.810 ;
        RECT 1380.160 324.770 1380.300 330.490 ;
        RECT 1379.700 324.630 1380.300 324.770 ;
        RECT 1379.700 317.550 1379.840 324.630 ;
        RECT 1379.640 317.230 1379.900 317.550 ;
        RECT 1378.720 268.950 1378.980 269.270 ;
        RECT 1378.780 265.870 1378.920 268.950 ;
        RECT 1378.720 265.550 1378.980 265.870 ;
        RECT 1379.640 265.550 1379.900 265.870 ;
        RECT 1379.700 241.390 1379.840 265.550 ;
        RECT 1379.180 241.070 1379.440 241.390 ;
        RECT 1379.640 241.070 1379.900 241.390 ;
        RECT 1379.240 193.110 1379.380 241.070 ;
        RECT 1379.180 192.790 1379.440 193.110 ;
        RECT 1379.640 165.930 1379.900 166.250 ;
        RECT 1379.700 138.030 1379.840 165.930 ;
        RECT 1379.640 137.710 1379.900 138.030 ;
        RECT 1379.640 89.770 1379.900 90.090 ;
        RECT 1379.700 16.310 1379.840 89.770 ;
        RECT 1536.960 16.330 1537.220 16.650 ;
        RECT 1379.640 15.990 1379.900 16.310 ;
        RECT 1537.020 2.000 1537.160 16.330 ;
        RECT 1536.810 -4.000 1537.370 2.000 ;
      LAYER via2 ;
        RECT 1377.330 1097.720 1377.610 1098.000 ;
        RECT 1379.170 1097.040 1379.450 1097.320 ;
      LAYER met3 ;
        RECT 1377.305 1098.010 1377.635 1098.025 ;
        RECT 1377.305 1097.710 1379.690 1098.010 ;
        RECT 1377.305 1097.695 1377.635 1097.710 ;
        RECT 1379.390 1097.345 1379.690 1097.710 ;
        RECT 1379.145 1097.030 1379.690 1097.345 ;
        RECT 1379.145 1097.015 1379.475 1097.030 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1386.125 917.745 1386.295 1000.535 ;
        RECT 1385.665 862.665 1385.835 910.775 ;
        RECT 1386.125 620.925 1386.295 669.375 ;
        RECT 1386.125 572.645 1386.295 593.895 ;
        RECT 1386.125 524.705 1386.295 572.135 ;
        RECT 1385.665 476.085 1385.835 524.195 ;
        RECT 1385.665 241.485 1385.835 317.475 ;
        RECT 1385.665 48.365 1385.835 137.955 ;
        RECT 1430.285 20.145 1431.375 20.315 ;
      LAYER mcon ;
        RECT 1386.125 1000.365 1386.295 1000.535 ;
        RECT 1385.665 910.605 1385.835 910.775 ;
        RECT 1386.125 669.205 1386.295 669.375 ;
        RECT 1386.125 593.725 1386.295 593.895 ;
        RECT 1386.125 571.965 1386.295 572.135 ;
        RECT 1385.665 524.025 1385.835 524.195 ;
        RECT 1385.665 317.305 1385.835 317.475 ;
        RECT 1385.665 137.785 1385.835 137.955 ;
        RECT 1431.205 20.145 1431.375 20.315 ;
      LAYER met1 ;
        RECT 1386.050 1000.520 1386.370 1000.580 ;
        RECT 1385.855 1000.380 1386.370 1000.520 ;
        RECT 1386.050 1000.320 1386.370 1000.380 ;
        RECT 1386.050 917.900 1386.370 917.960 ;
        RECT 1385.855 917.760 1386.370 917.900 ;
        RECT 1386.050 917.700 1386.370 917.760 ;
        RECT 1385.605 910.760 1385.895 910.805 ;
        RECT 1386.050 910.760 1386.370 910.820 ;
        RECT 1385.605 910.620 1386.370 910.760 ;
        RECT 1385.605 910.575 1385.895 910.620 ;
        RECT 1386.050 910.560 1386.370 910.620 ;
        RECT 1385.590 862.820 1385.910 862.880 ;
        RECT 1385.395 862.680 1385.910 862.820 ;
        RECT 1385.590 862.620 1385.910 862.680 ;
        RECT 1385.130 765.920 1385.450 765.980 ;
        RECT 1385.590 765.920 1385.910 765.980 ;
        RECT 1385.130 765.780 1385.910 765.920 ;
        RECT 1385.130 765.720 1385.450 765.780 ;
        RECT 1385.590 765.720 1385.910 765.780 ;
        RECT 1386.050 669.360 1386.370 669.420 ;
        RECT 1385.855 669.220 1386.370 669.360 ;
        RECT 1386.050 669.160 1386.370 669.220 ;
        RECT 1386.050 621.080 1386.370 621.140 ;
        RECT 1385.855 620.940 1386.370 621.080 ;
        RECT 1386.050 620.880 1386.370 620.940 ;
        RECT 1386.050 593.880 1386.370 593.940 ;
        RECT 1385.855 593.740 1386.370 593.880 ;
        RECT 1386.050 593.680 1386.370 593.740 ;
        RECT 1386.065 572.615 1386.355 572.845 ;
        RECT 1386.140 572.165 1386.280 572.615 ;
        RECT 1386.065 571.935 1386.355 572.165 ;
        RECT 1386.050 524.860 1386.370 524.920 ;
        RECT 1385.855 524.720 1386.370 524.860 ;
        RECT 1386.050 524.660 1386.370 524.720 ;
        RECT 1385.605 524.180 1385.895 524.225 ;
        RECT 1386.050 524.180 1386.370 524.240 ;
        RECT 1385.605 524.040 1386.370 524.180 ;
        RECT 1385.605 523.995 1385.895 524.040 ;
        RECT 1386.050 523.980 1386.370 524.040 ;
        RECT 1385.590 476.240 1385.910 476.300 ;
        RECT 1385.395 476.100 1385.910 476.240 ;
        RECT 1385.590 476.040 1385.910 476.100 ;
        RECT 1385.590 373.220 1385.910 373.280 ;
        RECT 1386.050 373.220 1386.370 373.280 ;
        RECT 1385.590 373.080 1386.370 373.220 ;
        RECT 1385.590 373.020 1385.910 373.080 ;
        RECT 1386.050 373.020 1386.370 373.080 ;
        RECT 1385.605 317.460 1385.895 317.505 ;
        RECT 1386.050 317.460 1386.370 317.520 ;
        RECT 1385.605 317.320 1386.370 317.460 ;
        RECT 1385.605 317.275 1385.895 317.320 ;
        RECT 1386.050 317.260 1386.370 317.320 ;
        RECT 1385.605 241.640 1385.895 241.685 ;
        RECT 1386.050 241.640 1386.370 241.700 ;
        RECT 1385.605 241.500 1386.370 241.640 ;
        RECT 1385.605 241.455 1385.895 241.500 ;
        RECT 1386.050 241.440 1386.370 241.500 ;
        RECT 1385.605 137.940 1385.895 137.985 ;
        RECT 1386.050 137.940 1386.370 138.000 ;
        RECT 1385.605 137.800 1386.370 137.940 ;
        RECT 1385.605 137.755 1385.895 137.800 ;
        RECT 1386.050 137.740 1386.370 137.800 ;
        RECT 1385.605 48.520 1385.895 48.565 ;
        RECT 1386.050 48.520 1386.370 48.580 ;
        RECT 1385.605 48.380 1386.370 48.520 ;
        RECT 1385.605 48.335 1385.895 48.380 ;
        RECT 1386.050 48.320 1386.370 48.380 ;
        RECT 1386.050 20.980 1386.370 21.040 ;
        RECT 1386.050 20.840 1389.040 20.980 ;
        RECT 1386.050 20.780 1386.370 20.840 ;
        RECT 1388.900 20.640 1389.040 20.840 ;
        RECT 1388.900 20.500 1391.340 20.640 ;
        RECT 1391.200 20.300 1391.340 20.500 ;
        RECT 1430.225 20.300 1430.515 20.345 ;
        RECT 1391.200 20.160 1430.515 20.300 ;
        RECT 1430.225 20.115 1430.515 20.160 ;
        RECT 1431.145 20.300 1431.435 20.345 ;
        RECT 1554.870 20.300 1555.190 20.360 ;
        RECT 1431.145 20.160 1555.190 20.300 ;
        RECT 1431.145 20.115 1431.435 20.160 ;
        RECT 1554.870 20.100 1555.190 20.160 ;
      LAYER via ;
        RECT 1386.080 1000.320 1386.340 1000.580 ;
        RECT 1386.080 917.700 1386.340 917.960 ;
        RECT 1386.080 910.560 1386.340 910.820 ;
        RECT 1385.620 862.620 1385.880 862.880 ;
        RECT 1385.160 765.720 1385.420 765.980 ;
        RECT 1385.620 765.720 1385.880 765.980 ;
        RECT 1386.080 669.160 1386.340 669.420 ;
        RECT 1386.080 620.880 1386.340 621.140 ;
        RECT 1386.080 593.680 1386.340 593.940 ;
        RECT 1386.080 524.660 1386.340 524.920 ;
        RECT 1386.080 523.980 1386.340 524.240 ;
        RECT 1385.620 476.040 1385.880 476.300 ;
        RECT 1385.620 373.020 1385.880 373.280 ;
        RECT 1386.080 373.020 1386.340 373.280 ;
        RECT 1386.080 317.260 1386.340 317.520 ;
        RECT 1386.080 241.440 1386.340 241.700 ;
        RECT 1386.080 137.740 1386.340 138.000 ;
        RECT 1386.080 48.320 1386.340 48.580 ;
        RECT 1386.080 20.780 1386.340 21.040 ;
        RECT 1554.900 20.100 1555.160 20.360 ;
      LAYER met2 ;
        RECT 1383.230 1101.330 1383.510 1104.000 ;
        RECT 1383.230 1101.190 1385.360 1101.330 ;
        RECT 1383.230 1100.000 1383.510 1101.190 ;
        RECT 1385.220 1062.570 1385.360 1101.190 ;
        RECT 1384.760 1062.430 1385.360 1062.570 ;
        RECT 1384.760 1007.605 1384.900 1062.430 ;
        RECT 1384.690 1007.235 1384.970 1007.605 ;
        RECT 1386.070 1007.235 1386.350 1007.605 ;
        RECT 1386.140 1000.610 1386.280 1007.235 ;
        RECT 1386.080 1000.290 1386.340 1000.610 ;
        RECT 1386.080 917.670 1386.340 917.990 ;
        RECT 1386.140 910.850 1386.280 917.670 ;
        RECT 1386.080 910.530 1386.340 910.850 ;
        RECT 1385.620 862.590 1385.880 862.910 ;
        RECT 1385.680 838.170 1385.820 862.590 ;
        RECT 1385.220 838.030 1385.820 838.170 ;
        RECT 1385.220 814.485 1385.360 838.030 ;
        RECT 1385.150 814.115 1385.430 814.485 ;
        RECT 1385.160 765.690 1385.420 766.010 ;
        RECT 1385.610 765.835 1385.890 766.205 ;
        RECT 1385.620 765.690 1385.880 765.835 ;
        RECT 1385.220 717.925 1385.360 765.690 ;
        RECT 1385.150 717.555 1385.430 717.925 ;
        RECT 1386.070 717.555 1386.350 717.925 ;
        RECT 1386.140 669.450 1386.280 717.555 ;
        RECT 1386.080 669.130 1386.340 669.450 ;
        RECT 1386.080 620.850 1386.340 621.170 ;
        RECT 1386.140 593.970 1386.280 620.850 ;
        RECT 1386.080 593.650 1386.340 593.970 ;
        RECT 1386.080 524.630 1386.340 524.950 ;
        RECT 1386.140 524.270 1386.280 524.630 ;
        RECT 1386.080 523.950 1386.340 524.270 ;
        RECT 1385.620 476.010 1385.880 476.330 ;
        RECT 1385.680 448.530 1385.820 476.010 ;
        RECT 1385.680 448.390 1386.280 448.530 ;
        RECT 1386.140 373.310 1386.280 448.390 ;
        RECT 1385.620 372.990 1385.880 373.310 ;
        RECT 1386.080 372.990 1386.340 373.310 ;
        RECT 1385.680 348.570 1385.820 372.990 ;
        RECT 1385.680 348.430 1386.280 348.570 ;
        RECT 1386.140 317.550 1386.280 348.430 ;
        RECT 1386.080 317.230 1386.340 317.550 ;
        RECT 1386.080 241.410 1386.340 241.730 ;
        RECT 1386.140 193.530 1386.280 241.410 ;
        RECT 1385.680 193.390 1386.280 193.530 ;
        RECT 1385.680 157.490 1385.820 193.390 ;
        RECT 1385.680 157.350 1386.280 157.490 ;
        RECT 1386.140 138.030 1386.280 157.350 ;
        RECT 1386.080 137.710 1386.340 138.030 ;
        RECT 1386.080 48.290 1386.340 48.610 ;
        RECT 1386.140 21.070 1386.280 48.290 ;
        RECT 1386.080 20.750 1386.340 21.070 ;
        RECT 1554.900 20.070 1555.160 20.390 ;
        RECT 1554.960 2.000 1555.100 20.070 ;
        RECT 1554.750 -4.000 1555.310 2.000 ;
      LAYER via2 ;
        RECT 1384.690 1007.280 1384.970 1007.560 ;
        RECT 1386.070 1007.280 1386.350 1007.560 ;
        RECT 1385.150 814.160 1385.430 814.440 ;
        RECT 1385.610 765.880 1385.890 766.160 ;
        RECT 1385.150 717.600 1385.430 717.880 ;
        RECT 1386.070 717.600 1386.350 717.880 ;
      LAYER met3 ;
        RECT 1384.665 1007.570 1384.995 1007.585 ;
        RECT 1386.045 1007.570 1386.375 1007.585 ;
        RECT 1384.665 1007.270 1386.375 1007.570 ;
        RECT 1384.665 1007.255 1384.995 1007.270 ;
        RECT 1386.045 1007.255 1386.375 1007.270 ;
        RECT 1385.125 814.450 1385.455 814.465 ;
        RECT 1385.125 814.150 1386.130 814.450 ;
        RECT 1385.125 814.135 1385.455 814.150 ;
        RECT 1385.830 813.780 1386.130 814.150 ;
        RECT 1385.790 813.460 1386.170 813.780 ;
        RECT 1385.585 766.180 1385.915 766.185 ;
        RECT 1385.585 766.170 1386.170 766.180 ;
        RECT 1385.360 765.870 1386.170 766.170 ;
        RECT 1385.585 765.860 1386.170 765.870 ;
        RECT 1385.585 765.855 1385.915 765.860 ;
        RECT 1385.125 717.890 1385.455 717.905 ;
        RECT 1386.045 717.890 1386.375 717.905 ;
        RECT 1385.125 717.590 1386.375 717.890 ;
        RECT 1385.125 717.575 1385.455 717.590 ;
        RECT 1386.045 717.575 1386.375 717.590 ;
      LAYER via3 ;
        RECT 1385.820 813.460 1386.140 813.780 ;
        RECT 1385.820 765.860 1386.140 766.180 ;
      LAYER met4 ;
        RECT 1385.815 813.455 1386.145 813.785 ;
        RECT 1385.830 766.185 1386.130 813.455 ;
        RECT 1385.815 765.855 1386.145 766.185 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1438.565 18.445 1438.735 19.975 ;
      LAYER mcon ;
        RECT 1438.565 19.805 1438.735 19.975 ;
      LAYER met1 ;
        RECT 1389.730 1088.580 1390.050 1088.640 ;
        RECT 1393.410 1088.580 1393.730 1088.640 ;
        RECT 1389.730 1088.440 1393.730 1088.580 ;
        RECT 1389.730 1088.380 1390.050 1088.440 ;
        RECT 1393.410 1088.380 1393.730 1088.440 ;
        RECT 1438.505 19.960 1438.795 20.005 ;
        RECT 1572.810 19.960 1573.130 20.020 ;
        RECT 1438.505 19.820 1573.130 19.960 ;
        RECT 1438.505 19.775 1438.795 19.820 ;
        RECT 1572.810 19.760 1573.130 19.820 ;
        RECT 1393.410 18.600 1393.730 18.660 ;
        RECT 1438.505 18.600 1438.795 18.645 ;
        RECT 1393.410 18.460 1438.795 18.600 ;
        RECT 1393.410 18.400 1393.730 18.460 ;
        RECT 1438.505 18.415 1438.795 18.460 ;
      LAYER via ;
        RECT 1389.760 1088.380 1390.020 1088.640 ;
        RECT 1393.440 1088.380 1393.700 1088.640 ;
        RECT 1572.840 19.760 1573.100 20.020 ;
        RECT 1393.440 18.400 1393.700 18.660 ;
      LAYER met2 ;
        RECT 1389.670 1100.580 1389.950 1104.000 ;
        RECT 1389.670 1100.000 1389.960 1100.580 ;
        RECT 1389.820 1088.670 1389.960 1100.000 ;
        RECT 1389.760 1088.350 1390.020 1088.670 ;
        RECT 1393.440 1088.350 1393.700 1088.670 ;
        RECT 1393.500 18.690 1393.640 1088.350 ;
        RECT 1572.840 19.730 1573.100 20.050 ;
        RECT 1393.440 18.370 1393.700 18.690 ;
        RECT 1572.900 2.000 1573.040 19.730 ;
        RECT 1572.690 -4.000 1573.250 2.000 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1395.710 1088.580 1396.030 1088.640 ;
        RECT 1400.310 1088.580 1400.630 1088.640 ;
        RECT 1395.710 1088.440 1400.630 1088.580 ;
        RECT 1395.710 1088.380 1396.030 1088.440 ;
        RECT 1400.310 1088.380 1400.630 1088.440 ;
        RECT 1590.290 19.620 1590.610 19.680 ;
        RECT 1438.580 19.480 1590.610 19.620 ;
        RECT 1400.310 18.940 1400.630 19.000 ;
        RECT 1438.580 18.940 1438.720 19.480 ;
        RECT 1590.290 19.420 1590.610 19.480 ;
        RECT 1400.310 18.800 1438.720 18.940 ;
        RECT 1400.310 18.740 1400.630 18.800 ;
      LAYER via ;
        RECT 1395.740 1088.380 1396.000 1088.640 ;
        RECT 1400.340 1088.380 1400.600 1088.640 ;
        RECT 1400.340 18.740 1400.600 19.000 ;
        RECT 1590.320 19.420 1590.580 19.680 ;
      LAYER met2 ;
        RECT 1395.650 1100.580 1395.930 1104.000 ;
        RECT 1395.650 1100.000 1395.940 1100.580 ;
        RECT 1395.800 1088.670 1395.940 1100.000 ;
        RECT 1395.740 1088.350 1396.000 1088.670 ;
        RECT 1400.340 1088.350 1400.600 1088.670 ;
        RECT 1400.400 19.030 1400.540 1088.350 ;
        RECT 1590.320 19.390 1590.580 19.710 ;
        RECT 1400.340 18.710 1400.600 19.030 ;
        RECT 1590.380 2.000 1590.520 19.390 ;
        RECT 1590.170 -4.000 1590.730 2.000 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1401.690 1088.580 1402.010 1088.640 ;
        RECT 1407.210 1088.580 1407.530 1088.640 ;
        RECT 1401.690 1088.440 1407.530 1088.580 ;
        RECT 1401.690 1088.380 1402.010 1088.440 ;
        RECT 1407.210 1088.380 1407.530 1088.440 ;
        RECT 1608.230 19.280 1608.550 19.340 ;
        RECT 1439.040 19.140 1608.550 19.280 ;
        RECT 1407.210 18.260 1407.530 18.320 ;
        RECT 1439.040 18.260 1439.180 19.140 ;
        RECT 1608.230 19.080 1608.550 19.140 ;
        RECT 1407.210 18.120 1439.180 18.260 ;
        RECT 1407.210 18.060 1407.530 18.120 ;
      LAYER via ;
        RECT 1401.720 1088.380 1401.980 1088.640 ;
        RECT 1407.240 1088.380 1407.500 1088.640 ;
        RECT 1407.240 18.060 1407.500 18.320 ;
        RECT 1608.260 19.080 1608.520 19.340 ;
      LAYER met2 ;
        RECT 1401.630 1100.580 1401.910 1104.000 ;
        RECT 1401.630 1100.000 1401.920 1100.580 ;
        RECT 1401.780 1088.670 1401.920 1100.000 ;
        RECT 1401.720 1088.350 1401.980 1088.670 ;
        RECT 1407.240 1088.350 1407.500 1088.670 ;
        RECT 1407.300 18.350 1407.440 1088.350 ;
        RECT 1608.260 19.050 1608.520 19.370 ;
        RECT 1407.240 18.030 1407.500 18.350 ;
        RECT 1608.320 2.000 1608.460 19.050 ;
        RECT 1608.110 -4.000 1608.670 2.000 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1408.130 1087.560 1408.450 1087.620 ;
        RECT 1548.890 1087.560 1549.210 1087.620 ;
        RECT 1408.130 1087.420 1549.210 1087.560 ;
        RECT 1408.130 1087.360 1408.450 1087.420 ;
        RECT 1548.890 1087.360 1549.210 1087.420 ;
        RECT 1626.170 16.900 1626.490 16.960 ;
        RECT 1567.380 16.760 1626.490 16.900 ;
        RECT 1548.430 16.560 1548.750 16.620 ;
        RECT 1567.380 16.560 1567.520 16.760 ;
        RECT 1626.170 16.700 1626.490 16.760 ;
        RECT 1548.430 16.420 1567.520 16.560 ;
        RECT 1548.430 16.360 1548.750 16.420 ;
      LAYER via ;
        RECT 1408.160 1087.360 1408.420 1087.620 ;
        RECT 1548.920 1087.360 1549.180 1087.620 ;
        RECT 1548.460 16.360 1548.720 16.620 ;
        RECT 1626.200 16.700 1626.460 16.960 ;
      LAYER met2 ;
        RECT 1408.070 1100.580 1408.350 1104.000 ;
        RECT 1408.070 1100.000 1408.360 1100.580 ;
        RECT 1408.220 1087.650 1408.360 1100.000 ;
        RECT 1408.160 1087.330 1408.420 1087.650 ;
        RECT 1548.920 1087.330 1549.180 1087.650 ;
        RECT 1548.980 34.410 1549.120 1087.330 ;
        RECT 1548.520 34.270 1549.120 34.410 ;
        RECT 1548.520 16.650 1548.660 34.270 ;
        RECT 1626.200 16.670 1626.460 16.990 ;
        RECT 1548.460 16.330 1548.720 16.650 ;
        RECT 1626.260 2.000 1626.400 16.670 ;
        RECT 1626.050 -4.000 1626.610 2.000 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1449.145 1083.325 1449.315 1084.515 ;
        RECT 1496.985 1083.325 1497.155 1084.175 ;
        RECT 1510.785 1084.005 1510.955 1085.535 ;
      LAYER mcon ;
        RECT 1510.785 1085.365 1510.955 1085.535 ;
        RECT 1449.145 1084.345 1449.315 1084.515 ;
        RECT 1496.985 1084.005 1497.155 1084.175 ;
      LAYER met1 ;
        RECT 1510.725 1085.520 1511.015 1085.565 ;
        RECT 1583.390 1085.520 1583.710 1085.580 ;
        RECT 1510.725 1085.380 1583.710 1085.520 ;
        RECT 1510.725 1085.335 1511.015 1085.380 ;
        RECT 1583.390 1085.320 1583.710 1085.380 ;
        RECT 1414.110 1084.500 1414.430 1084.560 ;
        RECT 1449.085 1084.500 1449.375 1084.545 ;
        RECT 1414.110 1084.360 1449.375 1084.500 ;
        RECT 1414.110 1084.300 1414.430 1084.360 ;
        RECT 1449.085 1084.315 1449.375 1084.360 ;
        RECT 1496.925 1084.160 1497.215 1084.205 ;
        RECT 1510.725 1084.160 1511.015 1084.205 ;
        RECT 1496.925 1084.020 1511.015 1084.160 ;
        RECT 1496.925 1083.975 1497.215 1084.020 ;
        RECT 1510.725 1083.975 1511.015 1084.020 ;
        RECT 1449.085 1083.480 1449.375 1083.525 ;
        RECT 1496.925 1083.480 1497.215 1083.525 ;
        RECT 1449.085 1083.340 1497.215 1083.480 ;
        RECT 1449.085 1083.295 1449.375 1083.340 ;
        RECT 1496.925 1083.295 1497.215 1083.340 ;
        RECT 1583.390 19.960 1583.710 20.020 ;
        RECT 1644.110 19.960 1644.430 20.020 ;
        RECT 1583.390 19.820 1644.430 19.960 ;
        RECT 1583.390 19.760 1583.710 19.820 ;
        RECT 1644.110 19.760 1644.430 19.820 ;
      LAYER via ;
        RECT 1583.420 1085.320 1583.680 1085.580 ;
        RECT 1414.140 1084.300 1414.400 1084.560 ;
        RECT 1583.420 19.760 1583.680 20.020 ;
        RECT 1644.140 19.760 1644.400 20.020 ;
      LAYER met2 ;
        RECT 1414.050 1100.580 1414.330 1104.000 ;
        RECT 1414.050 1100.000 1414.340 1100.580 ;
        RECT 1414.200 1084.590 1414.340 1100.000 ;
        RECT 1583.420 1085.290 1583.680 1085.610 ;
        RECT 1414.140 1084.270 1414.400 1084.590 ;
        RECT 1583.480 20.050 1583.620 1085.290 ;
        RECT 1583.420 19.730 1583.680 20.050 ;
        RECT 1644.140 19.730 1644.400 20.050 ;
        RECT 1644.200 2.000 1644.340 19.730 ;
        RECT 1643.990 -4.000 1644.550 2.000 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1421.010 193.500 1421.330 193.760 ;
        RECT 1421.100 193.080 1421.240 193.500 ;
        RECT 1421.010 192.820 1421.330 193.080 ;
      LAYER via ;
        RECT 1421.040 193.500 1421.300 193.760 ;
        RECT 1421.040 192.820 1421.300 193.080 ;
      LAYER met2 ;
        RECT 1420.030 1100.650 1420.310 1104.000 ;
        RECT 1420.030 1100.510 1421.240 1100.650 ;
        RECT 1420.030 1100.000 1420.310 1100.510 ;
        RECT 1421.100 193.790 1421.240 1100.510 ;
        RECT 1421.040 193.470 1421.300 193.790 ;
        RECT 1421.040 192.790 1421.300 193.110 ;
        RECT 1421.100 16.845 1421.240 192.790 ;
        RECT 1421.030 16.475 1421.310 16.845 ;
        RECT 1662.070 16.475 1662.350 16.845 ;
        RECT 1662.140 2.000 1662.280 16.475 ;
        RECT 1661.930 -4.000 1662.490 2.000 ;
      LAYER via2 ;
        RECT 1421.030 16.520 1421.310 16.800 ;
        RECT 1662.070 16.520 1662.350 16.800 ;
      LAYER met3 ;
        RECT 1421.005 16.810 1421.335 16.825 ;
        RECT 1662.045 16.810 1662.375 16.825 ;
        RECT 1421.005 16.510 1662.375 16.810 ;
        RECT 1421.005 16.495 1421.335 16.510 ;
        RECT 1662.045 16.495 1662.375 16.510 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1427.910 19.620 1428.230 19.680 ;
        RECT 1438.030 19.620 1438.350 19.680 ;
        RECT 1427.910 19.480 1438.350 19.620 ;
        RECT 1427.910 19.420 1428.230 19.480 ;
        RECT 1438.030 19.420 1438.350 19.480 ;
        RECT 1439.870 18.940 1440.190 19.000 ;
        RECT 1679.530 18.940 1679.850 19.000 ;
        RECT 1439.870 18.800 1679.850 18.940 ;
        RECT 1439.870 18.740 1440.190 18.800 ;
        RECT 1679.530 18.740 1679.850 18.800 ;
      LAYER via ;
        RECT 1427.940 19.420 1428.200 19.680 ;
        RECT 1438.060 19.420 1438.320 19.680 ;
        RECT 1439.900 18.740 1440.160 19.000 ;
        RECT 1679.560 18.740 1679.820 19.000 ;
      LAYER met2 ;
        RECT 1426.470 1100.650 1426.750 1104.000 ;
        RECT 1426.470 1100.510 1428.140 1100.650 ;
        RECT 1426.470 1100.000 1426.750 1100.510 ;
        RECT 1428.000 19.710 1428.140 1100.510 ;
        RECT 1427.940 19.390 1428.200 19.710 ;
        RECT 1438.060 19.450 1438.320 19.710 ;
        RECT 1438.060 19.390 1440.100 19.450 ;
        RECT 1438.120 19.310 1440.100 19.390 ;
        RECT 1439.960 19.030 1440.100 19.310 ;
        RECT 1439.900 18.710 1440.160 19.030 ;
        RECT 1679.560 18.710 1679.820 19.030 ;
        RECT 1679.620 2.000 1679.760 18.710 ;
        RECT 1679.410 -4.000 1679.970 2.000 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1439.485 18.445 1439.655 20.655 ;
      LAYER mcon ;
        RECT 1439.485 20.485 1439.655 20.655 ;
      LAYER met1 ;
        RECT 1432.510 1089.600 1432.830 1089.660 ;
        RECT 1434.810 1089.600 1435.130 1089.660 ;
        RECT 1432.510 1089.460 1435.130 1089.600 ;
        RECT 1432.510 1089.400 1432.830 1089.460 ;
        RECT 1434.810 1089.400 1435.130 1089.460 ;
        RECT 1434.810 20.640 1435.130 20.700 ;
        RECT 1439.425 20.640 1439.715 20.685 ;
        RECT 1434.810 20.500 1439.715 20.640 ;
        RECT 1434.810 20.440 1435.130 20.500 ;
        RECT 1439.425 20.455 1439.715 20.500 ;
        RECT 1439.425 18.600 1439.715 18.645 ;
        RECT 1697.470 18.600 1697.790 18.660 ;
        RECT 1439.425 18.460 1697.790 18.600 ;
        RECT 1439.425 18.415 1439.715 18.460 ;
        RECT 1697.470 18.400 1697.790 18.460 ;
      LAYER via ;
        RECT 1432.540 1089.400 1432.800 1089.660 ;
        RECT 1434.840 1089.400 1435.100 1089.660 ;
        RECT 1434.840 20.440 1435.100 20.700 ;
        RECT 1697.500 18.400 1697.760 18.660 ;
      LAYER met2 ;
        RECT 1432.450 1100.580 1432.730 1104.000 ;
        RECT 1432.450 1100.000 1432.740 1100.580 ;
        RECT 1432.600 1089.690 1432.740 1100.000 ;
        RECT 1432.540 1089.370 1432.800 1089.690 ;
        RECT 1434.840 1089.370 1435.100 1089.690 ;
        RECT 1434.900 20.730 1435.040 1089.370 ;
        RECT 1434.840 20.410 1435.100 20.730 ;
        RECT 1697.500 18.370 1697.760 18.690 ;
        RECT 1697.560 2.000 1697.700 18.370 ;
        RECT 1697.350 -4.000 1697.910 2.000 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1099.085 1014.305 1099.255 1028.415 ;
        RECT 1099.085 517.905 1099.255 565.675 ;
        RECT 1098.625 469.285 1098.795 517.395 ;
        RECT 1098.625 331.245 1098.795 352.495 ;
        RECT 1099.085 179.605 1099.255 212.415 ;
      LAYER mcon ;
        RECT 1099.085 1028.245 1099.255 1028.415 ;
        RECT 1099.085 565.505 1099.255 565.675 ;
        RECT 1098.625 517.225 1098.795 517.395 ;
        RECT 1098.625 352.325 1098.795 352.495 ;
        RECT 1099.085 212.245 1099.255 212.415 ;
      LAYER met1 ;
        RECT 1099.010 1078.720 1099.330 1078.780 ;
        RECT 1101.770 1078.720 1102.090 1078.780 ;
        RECT 1099.010 1078.580 1102.090 1078.720 ;
        RECT 1099.010 1078.520 1099.330 1078.580 ;
        RECT 1101.770 1078.520 1102.090 1078.580 ;
        RECT 1099.010 1028.400 1099.330 1028.460 ;
        RECT 1098.815 1028.260 1099.330 1028.400 ;
        RECT 1099.010 1028.200 1099.330 1028.260 ;
        RECT 1099.010 1014.460 1099.330 1014.520 ;
        RECT 1098.815 1014.320 1099.330 1014.460 ;
        RECT 1099.010 1014.260 1099.330 1014.320 ;
        RECT 1099.010 980.120 1099.330 980.180 ;
        RECT 1098.640 979.980 1099.330 980.120 ;
        RECT 1098.640 979.840 1098.780 979.980 ;
        RECT 1099.010 979.920 1099.330 979.980 ;
        RECT 1098.550 979.580 1098.870 979.840 ;
        RECT 1099.010 869.620 1099.330 869.680 ;
        RECT 1099.930 869.620 1100.250 869.680 ;
        RECT 1099.010 869.480 1100.250 869.620 ;
        RECT 1099.010 869.420 1099.330 869.480 ;
        RECT 1099.930 869.420 1100.250 869.480 ;
        RECT 1099.025 565.660 1099.315 565.705 ;
        RECT 1099.470 565.660 1099.790 565.720 ;
        RECT 1099.025 565.520 1099.790 565.660 ;
        RECT 1099.025 565.475 1099.315 565.520 ;
        RECT 1099.470 565.460 1099.790 565.520 ;
        RECT 1099.010 518.060 1099.330 518.120 ;
        RECT 1098.815 517.920 1099.330 518.060 ;
        RECT 1099.010 517.860 1099.330 517.920 ;
        RECT 1098.565 517.380 1098.855 517.425 ;
        RECT 1099.010 517.380 1099.330 517.440 ;
        RECT 1098.565 517.240 1099.330 517.380 ;
        RECT 1098.565 517.195 1098.855 517.240 ;
        RECT 1099.010 517.180 1099.330 517.240 ;
        RECT 1098.550 469.440 1098.870 469.500 ;
        RECT 1098.355 469.300 1098.870 469.440 ;
        RECT 1098.550 469.240 1098.870 469.300 ;
        RECT 1097.630 421.160 1097.950 421.220 ;
        RECT 1099.010 421.160 1099.330 421.220 ;
        RECT 1097.630 421.020 1099.330 421.160 ;
        RECT 1097.630 420.960 1097.950 421.020 ;
        RECT 1099.010 420.960 1099.330 421.020 ;
        RECT 1098.565 352.480 1098.855 352.525 ;
        RECT 1099.010 352.480 1099.330 352.540 ;
        RECT 1098.565 352.340 1099.330 352.480 ;
        RECT 1098.565 352.295 1098.855 352.340 ;
        RECT 1099.010 352.280 1099.330 352.340 ;
        RECT 1098.550 331.400 1098.870 331.460 ;
        RECT 1098.355 331.260 1098.870 331.400 ;
        RECT 1098.550 331.200 1098.870 331.260 ;
        RECT 1098.550 283.120 1098.870 283.180 ;
        RECT 1099.010 283.120 1099.330 283.180 ;
        RECT 1098.550 282.980 1099.330 283.120 ;
        RECT 1098.550 282.920 1098.870 282.980 ;
        RECT 1099.010 282.920 1099.330 282.980 ;
        RECT 1099.010 212.400 1099.330 212.460 ;
        RECT 1098.815 212.260 1099.330 212.400 ;
        RECT 1099.010 212.200 1099.330 212.260 ;
        RECT 1099.025 179.760 1099.315 179.805 ;
        RECT 1099.930 179.760 1100.250 179.820 ;
        RECT 1099.025 179.620 1100.250 179.760 ;
        RECT 1099.025 179.575 1099.315 179.620 ;
        RECT 1099.930 179.560 1100.250 179.620 ;
        RECT 1099.010 138.280 1099.330 138.340 ;
        RECT 1099.930 138.280 1100.250 138.340 ;
        RECT 1099.010 138.140 1100.250 138.280 ;
        RECT 1099.010 138.080 1099.330 138.140 ;
        RECT 1099.930 138.080 1100.250 138.140 ;
        RECT 1098.550 90.340 1098.870 90.400 ;
        RECT 1098.550 90.200 1099.240 90.340 ;
        RECT 1098.550 90.140 1098.870 90.200 ;
        RECT 1099.100 90.060 1099.240 90.200 ;
        RECT 1099.010 89.800 1099.330 90.060 ;
        RECT 734.230 29.140 734.550 29.200 ;
        RECT 1099.010 29.140 1099.330 29.200 ;
        RECT 734.230 29.000 1099.330 29.140 ;
        RECT 734.230 28.940 734.550 29.000 ;
        RECT 1099.010 28.940 1099.330 29.000 ;
      LAYER via ;
        RECT 1099.040 1078.520 1099.300 1078.780 ;
        RECT 1101.800 1078.520 1102.060 1078.780 ;
        RECT 1099.040 1028.200 1099.300 1028.460 ;
        RECT 1099.040 1014.260 1099.300 1014.520 ;
        RECT 1099.040 979.920 1099.300 980.180 ;
        RECT 1098.580 979.580 1098.840 979.840 ;
        RECT 1099.040 869.420 1099.300 869.680 ;
        RECT 1099.960 869.420 1100.220 869.680 ;
        RECT 1099.500 565.460 1099.760 565.720 ;
        RECT 1099.040 517.860 1099.300 518.120 ;
        RECT 1099.040 517.180 1099.300 517.440 ;
        RECT 1098.580 469.240 1098.840 469.500 ;
        RECT 1097.660 420.960 1097.920 421.220 ;
        RECT 1099.040 420.960 1099.300 421.220 ;
        RECT 1099.040 352.280 1099.300 352.540 ;
        RECT 1098.580 331.200 1098.840 331.460 ;
        RECT 1098.580 282.920 1098.840 283.180 ;
        RECT 1099.040 282.920 1099.300 283.180 ;
        RECT 1099.040 212.200 1099.300 212.460 ;
        RECT 1099.960 179.560 1100.220 179.820 ;
        RECT 1099.040 138.080 1099.300 138.340 ;
        RECT 1099.960 138.080 1100.220 138.340 ;
        RECT 1098.580 90.140 1098.840 90.400 ;
        RECT 1099.040 89.800 1099.300 90.060 ;
        RECT 734.260 28.940 734.520 29.200 ;
        RECT 1099.040 28.940 1099.300 29.200 ;
      LAYER met2 ;
        RECT 1101.710 1100.580 1101.990 1104.000 ;
        RECT 1101.710 1100.000 1102.000 1100.580 ;
        RECT 1101.860 1078.810 1102.000 1100.000 ;
        RECT 1099.040 1078.490 1099.300 1078.810 ;
        RECT 1101.800 1078.490 1102.060 1078.810 ;
        RECT 1099.100 1028.490 1099.240 1078.490 ;
        RECT 1099.040 1028.170 1099.300 1028.490 ;
        RECT 1099.040 1014.230 1099.300 1014.550 ;
        RECT 1099.100 980.210 1099.240 1014.230 ;
        RECT 1099.040 979.890 1099.300 980.210 ;
        RECT 1098.580 979.550 1098.840 979.870 ;
        RECT 1098.640 966.125 1098.780 979.550 ;
        RECT 1098.570 965.755 1098.850 966.125 ;
        RECT 1099.950 965.755 1100.230 966.125 ;
        RECT 1100.020 869.710 1100.160 965.755 ;
        RECT 1099.040 869.390 1099.300 869.710 ;
        RECT 1099.960 869.390 1100.220 869.710 ;
        RECT 1099.100 787.170 1099.240 869.390 ;
        RECT 1098.640 787.030 1099.240 787.170 ;
        RECT 1098.640 786.490 1098.780 787.030 ;
        RECT 1098.640 786.350 1099.240 786.490 ;
        RECT 1099.100 681.770 1099.240 786.350 ;
        RECT 1099.100 681.630 1100.160 681.770 ;
        RECT 1100.020 669.645 1100.160 681.630 ;
        RECT 1099.030 669.275 1099.310 669.645 ;
        RECT 1099.950 669.275 1100.230 669.645 ;
        RECT 1099.100 589.970 1099.240 669.275 ;
        RECT 1099.100 589.830 1099.700 589.970 ;
        RECT 1099.560 565.750 1099.700 589.830 ;
        RECT 1099.500 565.430 1099.760 565.750 ;
        RECT 1099.040 517.830 1099.300 518.150 ;
        RECT 1099.100 517.470 1099.240 517.830 ;
        RECT 1099.040 517.150 1099.300 517.470 ;
        RECT 1098.580 469.210 1098.840 469.530 ;
        RECT 1098.640 469.045 1098.780 469.210 ;
        RECT 1097.650 468.675 1097.930 469.045 ;
        RECT 1098.570 468.675 1098.850 469.045 ;
        RECT 1097.720 421.250 1097.860 468.675 ;
        RECT 1097.660 420.930 1097.920 421.250 ;
        RECT 1099.040 420.930 1099.300 421.250 ;
        RECT 1099.100 352.570 1099.240 420.930 ;
        RECT 1099.040 352.250 1099.300 352.570 ;
        RECT 1098.580 331.170 1098.840 331.490 ;
        RECT 1098.640 283.210 1098.780 331.170 ;
        RECT 1098.580 282.890 1098.840 283.210 ;
        RECT 1099.040 282.890 1099.300 283.210 ;
        RECT 1099.100 256.770 1099.240 282.890 ;
        RECT 1098.640 256.630 1099.240 256.770 ;
        RECT 1098.640 255.410 1098.780 256.630 ;
        RECT 1098.640 255.270 1099.240 255.410 ;
        RECT 1099.100 212.490 1099.240 255.270 ;
        RECT 1099.040 212.170 1099.300 212.490 ;
        RECT 1099.960 179.530 1100.220 179.850 ;
        RECT 1100.020 138.370 1100.160 179.530 ;
        RECT 1099.040 138.050 1099.300 138.370 ;
        RECT 1099.960 138.050 1100.220 138.370 ;
        RECT 1099.100 137.770 1099.240 138.050 ;
        RECT 1098.640 137.630 1099.240 137.770 ;
        RECT 1098.640 90.430 1098.780 137.630 ;
        RECT 1098.580 90.110 1098.840 90.430 ;
        RECT 1099.040 89.770 1099.300 90.090 ;
        RECT 1099.100 29.230 1099.240 89.770 ;
        RECT 734.260 28.910 734.520 29.230 ;
        RECT 1099.040 28.910 1099.300 29.230 ;
        RECT 734.320 2.000 734.460 28.910 ;
        RECT 734.110 -4.000 734.670 2.000 ;
      LAYER via2 ;
        RECT 1098.570 965.800 1098.850 966.080 ;
        RECT 1099.950 965.800 1100.230 966.080 ;
        RECT 1099.030 669.320 1099.310 669.600 ;
        RECT 1099.950 669.320 1100.230 669.600 ;
        RECT 1097.650 468.720 1097.930 469.000 ;
        RECT 1098.570 468.720 1098.850 469.000 ;
      LAYER met3 ;
        RECT 1098.545 966.090 1098.875 966.105 ;
        RECT 1099.925 966.090 1100.255 966.105 ;
        RECT 1098.545 965.790 1100.255 966.090 ;
        RECT 1098.545 965.775 1098.875 965.790 ;
        RECT 1099.925 965.775 1100.255 965.790 ;
        RECT 1099.005 669.610 1099.335 669.625 ;
        RECT 1099.925 669.610 1100.255 669.625 ;
        RECT 1099.005 669.310 1100.255 669.610 ;
        RECT 1099.005 669.295 1099.335 669.310 ;
        RECT 1099.925 669.295 1100.255 669.310 ;
        RECT 1097.625 469.010 1097.955 469.025 ;
        RECT 1098.545 469.010 1098.875 469.025 ;
        RECT 1097.625 468.710 1098.875 469.010 ;
        RECT 1097.625 468.695 1097.955 468.710 ;
        RECT 1098.545 468.695 1098.875 468.710 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1438.490 1089.600 1438.810 1089.660 ;
        RECT 1441.710 1089.600 1442.030 1089.660 ;
        RECT 1438.490 1089.460 1442.030 1089.600 ;
        RECT 1438.490 1089.400 1438.810 1089.460 ;
        RECT 1441.710 1089.400 1442.030 1089.460 ;
        RECT 1441.710 18.260 1442.030 18.320 ;
        RECT 1715.410 18.260 1715.730 18.320 ;
        RECT 1441.710 18.120 1715.730 18.260 ;
        RECT 1441.710 18.060 1442.030 18.120 ;
        RECT 1715.410 18.060 1715.730 18.120 ;
      LAYER via ;
        RECT 1438.520 1089.400 1438.780 1089.660 ;
        RECT 1441.740 1089.400 1442.000 1089.660 ;
        RECT 1441.740 18.060 1442.000 18.320 ;
        RECT 1715.440 18.060 1715.700 18.320 ;
      LAYER met2 ;
        RECT 1438.430 1100.580 1438.710 1104.000 ;
        RECT 1438.430 1100.000 1438.720 1100.580 ;
        RECT 1438.580 1089.690 1438.720 1100.000 ;
        RECT 1438.520 1089.370 1438.780 1089.690 ;
        RECT 1441.740 1089.370 1442.000 1089.690 ;
        RECT 1441.800 18.350 1441.940 1089.370 ;
        RECT 1441.740 18.030 1442.000 18.350 ;
        RECT 1715.440 18.030 1715.700 18.350 ;
        RECT 1715.500 2.000 1715.640 18.030 ;
        RECT 1715.290 -4.000 1715.850 2.000 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1446.845 689.605 1447.015 717.655 ;
        RECT 1446.385 379.525 1446.555 427.635 ;
        RECT 1446.845 282.965 1447.015 331.075 ;
        RECT 1446.385 40.205 1446.555 65.535 ;
      LAYER mcon ;
        RECT 1446.845 717.485 1447.015 717.655 ;
        RECT 1446.385 427.465 1446.555 427.635 ;
        RECT 1446.845 330.905 1447.015 331.075 ;
        RECT 1446.385 65.365 1446.555 65.535 ;
      LAYER met1 ;
        RECT 1444.930 1062.740 1445.250 1062.800 ;
        RECT 1446.770 1062.740 1447.090 1062.800 ;
        RECT 1444.930 1062.600 1447.090 1062.740 ;
        RECT 1444.930 1062.540 1445.250 1062.600 ;
        RECT 1446.770 1062.540 1447.090 1062.600 ;
        RECT 1445.850 1014.460 1446.170 1014.520 ;
        RECT 1447.230 1014.460 1447.550 1014.520 ;
        RECT 1445.850 1014.320 1447.550 1014.460 ;
        RECT 1445.850 1014.260 1446.170 1014.320 ;
        RECT 1447.230 1014.260 1447.550 1014.320 ;
        RECT 1446.310 966.180 1446.630 966.240 ;
        RECT 1447.230 966.180 1447.550 966.240 ;
        RECT 1446.310 966.040 1447.550 966.180 ;
        RECT 1446.310 965.980 1446.630 966.040 ;
        RECT 1447.230 965.980 1447.550 966.040 ;
        RECT 1446.310 917.900 1446.630 917.960 ;
        RECT 1447.230 917.900 1447.550 917.960 ;
        RECT 1446.310 917.760 1447.550 917.900 ;
        RECT 1446.310 917.700 1446.630 917.760 ;
        RECT 1447.230 917.700 1447.550 917.760 ;
        RECT 1446.310 869.620 1446.630 869.680 ;
        RECT 1447.230 869.620 1447.550 869.680 ;
        RECT 1446.310 869.480 1447.550 869.620 ;
        RECT 1446.310 869.420 1446.630 869.480 ;
        RECT 1447.230 869.420 1447.550 869.480 ;
        RECT 1446.770 821.000 1447.090 821.060 ;
        RECT 1447.230 821.000 1447.550 821.060 ;
        RECT 1446.770 820.860 1447.550 821.000 ;
        RECT 1446.770 820.800 1447.090 820.860 ;
        RECT 1447.230 820.800 1447.550 820.860 ;
        RECT 1446.310 814.200 1446.630 814.260 ;
        RECT 1447.230 814.200 1447.550 814.260 ;
        RECT 1446.310 814.060 1447.550 814.200 ;
        RECT 1446.310 814.000 1446.630 814.060 ;
        RECT 1447.230 814.000 1447.550 814.060 ;
        RECT 1446.770 717.640 1447.090 717.700 ;
        RECT 1446.575 717.500 1447.090 717.640 ;
        RECT 1446.770 717.440 1447.090 717.500 ;
        RECT 1446.770 689.760 1447.090 689.820 ;
        RECT 1446.575 689.620 1447.090 689.760 ;
        RECT 1446.770 689.560 1447.090 689.620 ;
        RECT 1446.770 628.220 1447.090 628.280 ;
        RECT 1447.230 628.220 1447.550 628.280 ;
        RECT 1446.770 628.080 1447.550 628.220 ;
        RECT 1446.770 628.020 1447.090 628.080 ;
        RECT 1447.230 628.020 1447.550 628.080 ;
        RECT 1445.850 579.600 1446.170 579.660 ;
        RECT 1447.230 579.600 1447.550 579.660 ;
        RECT 1445.850 579.460 1447.550 579.600 ;
        RECT 1445.850 579.400 1446.170 579.460 ;
        RECT 1447.230 579.400 1447.550 579.460 ;
        RECT 1446.325 427.620 1446.615 427.665 ;
        RECT 1446.770 427.620 1447.090 427.680 ;
        RECT 1446.325 427.480 1447.090 427.620 ;
        RECT 1446.325 427.435 1446.615 427.480 ;
        RECT 1446.770 427.420 1447.090 427.480 ;
        RECT 1446.310 379.680 1446.630 379.740 ;
        RECT 1446.115 379.540 1446.630 379.680 ;
        RECT 1446.310 379.480 1446.630 379.540 ;
        RECT 1446.310 338.200 1446.630 338.260 ;
        RECT 1446.770 338.200 1447.090 338.260 ;
        RECT 1446.310 338.060 1447.090 338.200 ;
        RECT 1446.310 338.000 1446.630 338.060 ;
        RECT 1446.770 338.000 1447.090 338.060 ;
        RECT 1446.770 331.060 1447.090 331.120 ;
        RECT 1446.575 330.920 1447.090 331.060 ;
        RECT 1446.770 330.860 1447.090 330.920 ;
        RECT 1446.785 283.120 1447.075 283.165 ;
        RECT 1447.230 283.120 1447.550 283.180 ;
        RECT 1446.785 282.980 1447.550 283.120 ;
        RECT 1446.785 282.935 1447.075 282.980 ;
        RECT 1447.230 282.920 1447.550 282.980 ;
        RECT 1446.770 241.640 1447.090 241.700 ;
        RECT 1447.230 241.640 1447.550 241.700 ;
        RECT 1446.770 241.500 1447.550 241.640 ;
        RECT 1446.770 241.440 1447.090 241.500 ;
        RECT 1447.230 241.440 1447.550 241.500 ;
        RECT 1446.310 145.080 1446.630 145.140 ;
        RECT 1447.230 145.080 1447.550 145.140 ;
        RECT 1446.310 144.940 1447.550 145.080 ;
        RECT 1446.310 144.880 1446.630 144.940 ;
        RECT 1447.230 144.880 1447.550 144.940 ;
        RECT 1446.310 65.520 1446.630 65.580 ;
        RECT 1446.115 65.380 1446.630 65.520 ;
        RECT 1446.310 65.320 1446.630 65.380 ;
        RECT 1446.325 40.360 1446.615 40.405 ;
        RECT 1733.350 40.360 1733.670 40.420 ;
        RECT 1446.325 40.220 1733.670 40.360 ;
        RECT 1446.325 40.175 1446.615 40.220 ;
        RECT 1733.350 40.160 1733.670 40.220 ;
      LAYER via ;
        RECT 1444.960 1062.540 1445.220 1062.800 ;
        RECT 1446.800 1062.540 1447.060 1062.800 ;
        RECT 1445.880 1014.260 1446.140 1014.520 ;
        RECT 1447.260 1014.260 1447.520 1014.520 ;
        RECT 1446.340 965.980 1446.600 966.240 ;
        RECT 1447.260 965.980 1447.520 966.240 ;
        RECT 1446.340 917.700 1446.600 917.960 ;
        RECT 1447.260 917.700 1447.520 917.960 ;
        RECT 1446.340 869.420 1446.600 869.680 ;
        RECT 1447.260 869.420 1447.520 869.680 ;
        RECT 1446.800 820.800 1447.060 821.060 ;
        RECT 1447.260 820.800 1447.520 821.060 ;
        RECT 1446.340 814.000 1446.600 814.260 ;
        RECT 1447.260 814.000 1447.520 814.260 ;
        RECT 1446.800 717.440 1447.060 717.700 ;
        RECT 1446.800 689.560 1447.060 689.820 ;
        RECT 1446.800 628.020 1447.060 628.280 ;
        RECT 1447.260 628.020 1447.520 628.280 ;
        RECT 1445.880 579.400 1446.140 579.660 ;
        RECT 1447.260 579.400 1447.520 579.660 ;
        RECT 1446.800 427.420 1447.060 427.680 ;
        RECT 1446.340 379.480 1446.600 379.740 ;
        RECT 1446.340 338.000 1446.600 338.260 ;
        RECT 1446.800 338.000 1447.060 338.260 ;
        RECT 1446.800 330.860 1447.060 331.120 ;
        RECT 1447.260 282.920 1447.520 283.180 ;
        RECT 1446.800 241.440 1447.060 241.700 ;
        RECT 1447.260 241.440 1447.520 241.700 ;
        RECT 1446.340 144.880 1446.600 145.140 ;
        RECT 1447.260 144.880 1447.520 145.140 ;
        RECT 1446.340 65.320 1446.600 65.580 ;
        RECT 1733.380 40.160 1733.640 40.420 ;
      LAYER met2 ;
        RECT 1444.870 1100.580 1445.150 1104.000 ;
        RECT 1444.870 1100.000 1445.160 1100.580 ;
        RECT 1445.020 1062.830 1445.160 1100.000 ;
        RECT 1444.960 1062.510 1445.220 1062.830 ;
        RECT 1446.800 1062.685 1447.060 1062.830 ;
        RECT 1445.870 1062.315 1446.150 1062.685 ;
        RECT 1446.790 1062.315 1447.070 1062.685 ;
        RECT 1445.940 1014.550 1446.080 1062.315 ;
        RECT 1445.880 1014.230 1446.140 1014.550 ;
        RECT 1447.260 1014.405 1447.520 1014.550 ;
        RECT 1446.330 1014.035 1446.610 1014.405 ;
        RECT 1447.250 1014.035 1447.530 1014.405 ;
        RECT 1446.400 966.270 1446.540 1014.035 ;
        RECT 1446.340 966.125 1446.600 966.270 ;
        RECT 1447.260 966.125 1447.520 966.270 ;
        RECT 1446.330 965.755 1446.610 966.125 ;
        RECT 1447.250 965.755 1447.530 966.125 ;
        RECT 1446.400 917.990 1446.540 965.755 ;
        RECT 1446.340 917.845 1446.600 917.990 ;
        RECT 1447.260 917.845 1447.520 917.990 ;
        RECT 1446.330 917.475 1446.610 917.845 ;
        RECT 1447.250 917.475 1447.530 917.845 ;
        RECT 1446.400 869.710 1446.540 917.475 ;
        RECT 1446.340 869.390 1446.600 869.710 ;
        RECT 1447.260 869.390 1447.520 869.710 ;
        RECT 1447.320 834.090 1447.460 869.390 ;
        RECT 1446.860 833.950 1447.460 834.090 ;
        RECT 1446.860 821.090 1447.000 833.950 ;
        RECT 1446.800 820.770 1447.060 821.090 ;
        RECT 1447.260 820.770 1447.520 821.090 ;
        RECT 1447.320 814.290 1447.460 820.770 ;
        RECT 1446.340 813.970 1446.600 814.290 ;
        RECT 1447.260 813.970 1447.520 814.290 ;
        RECT 1446.400 766.205 1446.540 813.970 ;
        RECT 1446.330 765.835 1446.610 766.205 ;
        RECT 1447.250 765.835 1447.530 766.205 ;
        RECT 1447.320 724.610 1447.460 765.835 ;
        RECT 1446.860 724.470 1447.460 724.610 ;
        RECT 1446.860 717.730 1447.000 724.470 ;
        RECT 1446.800 717.410 1447.060 717.730 ;
        RECT 1446.800 689.530 1447.060 689.850 ;
        RECT 1446.860 669.530 1447.000 689.530 ;
        RECT 1446.860 669.390 1447.460 669.530 ;
        RECT 1447.320 628.310 1447.460 669.390 ;
        RECT 1446.800 627.990 1447.060 628.310 ;
        RECT 1447.260 627.990 1447.520 628.310 ;
        RECT 1446.860 603.570 1447.000 627.990 ;
        RECT 1446.860 603.430 1447.460 603.570 ;
        RECT 1447.320 579.690 1447.460 603.430 ;
        RECT 1445.880 579.370 1446.140 579.690 ;
        RECT 1447.260 579.370 1447.520 579.690 ;
        RECT 1445.940 531.605 1446.080 579.370 ;
        RECT 1445.870 531.235 1446.150 531.605 ;
        RECT 1446.790 531.235 1447.070 531.605 ;
        RECT 1446.860 507.010 1447.000 531.235 ;
        RECT 1446.860 506.870 1447.460 507.010 ;
        RECT 1447.320 434.930 1447.460 506.870 ;
        RECT 1446.860 434.790 1447.460 434.930 ;
        RECT 1446.860 427.710 1447.000 434.790 ;
        RECT 1446.800 427.390 1447.060 427.710 ;
        RECT 1446.340 379.450 1446.600 379.770 ;
        RECT 1446.400 338.290 1446.540 379.450 ;
        RECT 1446.340 337.970 1446.600 338.290 ;
        RECT 1446.800 337.970 1447.060 338.290 ;
        RECT 1446.860 331.150 1447.000 337.970 ;
        RECT 1446.800 330.830 1447.060 331.150 ;
        RECT 1447.260 282.890 1447.520 283.210 ;
        RECT 1447.320 241.730 1447.460 282.890 ;
        RECT 1446.800 241.410 1447.060 241.730 ;
        RECT 1447.260 241.410 1447.520 241.730 ;
        RECT 1446.860 217.330 1447.000 241.410 ;
        RECT 1446.860 217.190 1447.460 217.330 ;
        RECT 1447.320 145.170 1447.460 217.190 ;
        RECT 1446.340 144.850 1446.600 145.170 ;
        RECT 1447.260 144.850 1447.520 145.170 ;
        RECT 1446.400 90.285 1446.540 144.850 ;
        RECT 1446.330 89.915 1446.610 90.285 ;
        RECT 1446.330 89.235 1446.610 89.605 ;
        RECT 1446.400 65.610 1446.540 89.235 ;
        RECT 1446.340 65.290 1446.600 65.610 ;
        RECT 1733.380 40.130 1733.640 40.450 ;
        RECT 1733.440 2.000 1733.580 40.130 ;
        RECT 1733.230 -4.000 1733.790 2.000 ;
      LAYER via2 ;
        RECT 1445.870 1062.360 1446.150 1062.640 ;
        RECT 1446.790 1062.360 1447.070 1062.640 ;
        RECT 1446.330 1014.080 1446.610 1014.360 ;
        RECT 1447.250 1014.080 1447.530 1014.360 ;
        RECT 1446.330 965.800 1446.610 966.080 ;
        RECT 1447.250 965.800 1447.530 966.080 ;
        RECT 1446.330 917.520 1446.610 917.800 ;
        RECT 1447.250 917.520 1447.530 917.800 ;
        RECT 1446.330 765.880 1446.610 766.160 ;
        RECT 1447.250 765.880 1447.530 766.160 ;
        RECT 1445.870 531.280 1446.150 531.560 ;
        RECT 1446.790 531.280 1447.070 531.560 ;
        RECT 1446.330 89.960 1446.610 90.240 ;
        RECT 1446.330 89.280 1446.610 89.560 ;
      LAYER met3 ;
        RECT 1445.845 1062.650 1446.175 1062.665 ;
        RECT 1446.765 1062.650 1447.095 1062.665 ;
        RECT 1445.845 1062.350 1447.095 1062.650 ;
        RECT 1445.845 1062.335 1446.175 1062.350 ;
        RECT 1446.765 1062.335 1447.095 1062.350 ;
        RECT 1446.305 1014.370 1446.635 1014.385 ;
        RECT 1447.225 1014.370 1447.555 1014.385 ;
        RECT 1446.305 1014.070 1447.555 1014.370 ;
        RECT 1446.305 1014.055 1446.635 1014.070 ;
        RECT 1447.225 1014.055 1447.555 1014.070 ;
        RECT 1446.305 966.090 1446.635 966.105 ;
        RECT 1447.225 966.090 1447.555 966.105 ;
        RECT 1446.305 965.790 1447.555 966.090 ;
        RECT 1446.305 965.775 1446.635 965.790 ;
        RECT 1447.225 965.775 1447.555 965.790 ;
        RECT 1446.305 917.810 1446.635 917.825 ;
        RECT 1447.225 917.810 1447.555 917.825 ;
        RECT 1446.305 917.510 1447.555 917.810 ;
        RECT 1446.305 917.495 1446.635 917.510 ;
        RECT 1447.225 917.495 1447.555 917.510 ;
        RECT 1446.305 766.170 1446.635 766.185 ;
        RECT 1447.225 766.170 1447.555 766.185 ;
        RECT 1446.305 765.870 1447.555 766.170 ;
        RECT 1446.305 765.855 1446.635 765.870 ;
        RECT 1447.225 765.855 1447.555 765.870 ;
        RECT 1445.845 531.570 1446.175 531.585 ;
        RECT 1446.765 531.570 1447.095 531.585 ;
        RECT 1445.845 531.270 1447.095 531.570 ;
        RECT 1445.845 531.255 1446.175 531.270 ;
        RECT 1446.765 531.255 1447.095 531.270 ;
        RECT 1446.305 89.935 1446.635 90.265 ;
        RECT 1446.320 89.585 1446.620 89.935 ;
        RECT 1446.305 89.255 1446.635 89.585 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1450.910 1086.540 1451.230 1086.600 ;
        RECT 1455.510 1086.540 1455.830 1086.600 ;
        RECT 1450.910 1086.400 1455.830 1086.540 ;
        RECT 1450.910 1086.340 1451.230 1086.400 ;
        RECT 1455.510 1086.340 1455.830 1086.400 ;
        RECT 1455.510 17.920 1455.830 17.980 ;
        RECT 1751.290 17.920 1751.610 17.980 ;
        RECT 1455.510 17.780 1751.610 17.920 ;
        RECT 1455.510 17.720 1455.830 17.780 ;
        RECT 1751.290 17.720 1751.610 17.780 ;
      LAYER via ;
        RECT 1450.940 1086.340 1451.200 1086.600 ;
        RECT 1455.540 1086.340 1455.800 1086.600 ;
        RECT 1455.540 17.720 1455.800 17.980 ;
        RECT 1751.320 17.720 1751.580 17.980 ;
      LAYER met2 ;
        RECT 1450.850 1100.580 1451.130 1104.000 ;
        RECT 1450.850 1100.000 1451.140 1100.580 ;
        RECT 1451.000 1086.630 1451.140 1100.000 ;
        RECT 1450.940 1086.310 1451.200 1086.630 ;
        RECT 1455.540 1086.310 1455.800 1086.630 ;
        RECT 1455.600 18.010 1455.740 1086.310 ;
        RECT 1455.540 17.690 1455.800 18.010 ;
        RECT 1751.320 17.690 1751.580 18.010 ;
        RECT 1751.380 2.000 1751.520 17.690 ;
        RECT 1751.170 -4.000 1751.730 2.000 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1456.890 1089.600 1457.210 1089.660 ;
        RECT 1462.410 1089.600 1462.730 1089.660 ;
        RECT 1456.890 1089.460 1462.730 1089.600 ;
        RECT 1456.890 1089.400 1457.210 1089.460 ;
        RECT 1462.410 1089.400 1462.730 1089.460 ;
        RECT 1462.410 17.580 1462.730 17.640 ;
        RECT 1768.770 17.580 1769.090 17.640 ;
        RECT 1462.410 17.440 1769.090 17.580 ;
        RECT 1462.410 17.380 1462.730 17.440 ;
        RECT 1768.770 17.380 1769.090 17.440 ;
      LAYER via ;
        RECT 1456.920 1089.400 1457.180 1089.660 ;
        RECT 1462.440 1089.400 1462.700 1089.660 ;
        RECT 1462.440 17.380 1462.700 17.640 ;
        RECT 1768.800 17.380 1769.060 17.640 ;
      LAYER met2 ;
        RECT 1456.830 1100.580 1457.110 1104.000 ;
        RECT 1456.830 1100.000 1457.120 1100.580 ;
        RECT 1456.980 1089.690 1457.120 1100.000 ;
        RECT 1456.920 1089.370 1457.180 1089.690 ;
        RECT 1462.440 1089.370 1462.700 1089.690 ;
        RECT 1462.500 17.670 1462.640 1089.370 ;
        RECT 1462.440 17.350 1462.700 17.670 ;
        RECT 1768.800 17.350 1769.060 17.670 ;
        RECT 1768.860 2.000 1769.000 17.350 ;
        RECT 1768.650 -4.000 1769.210 2.000 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1486.405 16.235 1486.575 17.255 ;
        RECT 1486.405 16.065 1487.495 16.235 ;
        RECT 1508.025 16.065 1508.195 17.255 ;
      LAYER mcon ;
        RECT 1486.405 17.085 1486.575 17.255 ;
        RECT 1508.025 17.085 1508.195 17.255 ;
        RECT 1487.325 16.065 1487.495 16.235 ;
      LAYER met1 ;
        RECT 1463.330 1088.580 1463.650 1088.640 ;
        RECT 1469.310 1088.580 1469.630 1088.640 ;
        RECT 1463.330 1088.440 1469.630 1088.580 ;
        RECT 1463.330 1088.380 1463.650 1088.440 ;
        RECT 1469.310 1088.380 1469.630 1088.440 ;
        RECT 1469.310 17.240 1469.630 17.300 ;
        RECT 1486.345 17.240 1486.635 17.285 ;
        RECT 1469.310 17.100 1486.635 17.240 ;
        RECT 1469.310 17.040 1469.630 17.100 ;
        RECT 1486.345 17.055 1486.635 17.100 ;
        RECT 1507.965 17.240 1508.255 17.285 ;
        RECT 1786.710 17.240 1787.030 17.300 ;
        RECT 1507.965 17.100 1787.030 17.240 ;
        RECT 1507.965 17.055 1508.255 17.100 ;
        RECT 1786.710 17.040 1787.030 17.100 ;
        RECT 1487.265 16.220 1487.555 16.265 ;
        RECT 1507.965 16.220 1508.255 16.265 ;
        RECT 1487.265 16.080 1508.255 16.220 ;
        RECT 1487.265 16.035 1487.555 16.080 ;
        RECT 1507.965 16.035 1508.255 16.080 ;
      LAYER via ;
        RECT 1463.360 1088.380 1463.620 1088.640 ;
        RECT 1469.340 1088.380 1469.600 1088.640 ;
        RECT 1469.340 17.040 1469.600 17.300 ;
        RECT 1786.740 17.040 1787.000 17.300 ;
      LAYER met2 ;
        RECT 1463.270 1100.580 1463.550 1104.000 ;
        RECT 1463.270 1100.000 1463.560 1100.580 ;
        RECT 1463.420 1088.670 1463.560 1100.000 ;
        RECT 1463.360 1088.350 1463.620 1088.670 ;
        RECT 1469.340 1088.350 1469.600 1088.670 ;
        RECT 1469.400 17.330 1469.540 1088.350 ;
        RECT 1469.340 17.010 1469.600 17.330 ;
        RECT 1786.740 17.010 1787.000 17.330 ;
        RECT 1786.800 2.000 1786.940 17.010 ;
        RECT 1786.590 -4.000 1787.150 2.000 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1469.310 1089.600 1469.630 1089.660 ;
        RECT 1597.190 1089.600 1597.510 1089.660 ;
        RECT 1469.310 1089.460 1597.510 1089.600 ;
        RECT 1469.310 1089.400 1469.630 1089.460 ;
        RECT 1597.190 1089.400 1597.510 1089.460 ;
        RECT 1597.190 15.200 1597.510 15.260 ;
        RECT 1804.650 15.200 1804.970 15.260 ;
        RECT 1597.190 15.060 1804.970 15.200 ;
        RECT 1597.190 15.000 1597.510 15.060 ;
        RECT 1804.650 15.000 1804.970 15.060 ;
      LAYER via ;
        RECT 1469.340 1089.400 1469.600 1089.660 ;
        RECT 1597.220 1089.400 1597.480 1089.660 ;
        RECT 1597.220 15.000 1597.480 15.260 ;
        RECT 1804.680 15.000 1804.940 15.260 ;
      LAYER met2 ;
        RECT 1469.250 1100.580 1469.530 1104.000 ;
        RECT 1469.250 1100.000 1469.540 1100.580 ;
        RECT 1469.400 1089.690 1469.540 1100.000 ;
        RECT 1469.340 1089.370 1469.600 1089.690 ;
        RECT 1597.220 1089.370 1597.480 1089.690 ;
        RECT 1597.280 15.290 1597.420 1089.370 ;
        RECT 1597.220 14.970 1597.480 15.290 ;
        RECT 1804.680 14.970 1804.940 15.290 ;
        RECT 1804.740 2.000 1804.880 14.970 ;
        RECT 1804.530 -4.000 1805.090 2.000 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1475.750 37.980 1476.070 38.040 ;
        RECT 1822.590 37.980 1822.910 38.040 ;
        RECT 1475.750 37.840 1822.910 37.980 ;
        RECT 1475.750 37.780 1476.070 37.840 ;
        RECT 1822.590 37.780 1822.910 37.840 ;
      LAYER via ;
        RECT 1475.780 37.780 1476.040 38.040 ;
        RECT 1822.620 37.780 1822.880 38.040 ;
      LAYER met2 ;
        RECT 1475.230 1100.650 1475.510 1104.000 ;
        RECT 1475.230 1100.510 1475.980 1100.650 ;
        RECT 1475.230 1100.000 1475.510 1100.510 ;
        RECT 1475.840 38.070 1475.980 1100.510 ;
        RECT 1475.780 37.750 1476.040 38.070 ;
        RECT 1822.620 37.750 1822.880 38.070 ;
        RECT 1822.680 2.000 1822.820 37.750 ;
        RECT 1822.470 -4.000 1823.030 2.000 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1482.190 73.680 1482.510 73.740 ;
        RECT 1835.470 73.680 1835.790 73.740 ;
        RECT 1482.190 73.540 1835.790 73.680 ;
        RECT 1482.190 73.480 1482.510 73.540 ;
        RECT 1835.470 73.480 1835.790 73.540 ;
        RECT 1835.470 2.620 1835.790 2.680 ;
        RECT 1840.070 2.620 1840.390 2.680 ;
        RECT 1835.470 2.480 1840.390 2.620 ;
        RECT 1835.470 2.420 1835.790 2.480 ;
        RECT 1840.070 2.420 1840.390 2.480 ;
      LAYER via ;
        RECT 1482.220 73.480 1482.480 73.740 ;
        RECT 1835.500 73.480 1835.760 73.740 ;
        RECT 1835.500 2.420 1835.760 2.680 ;
        RECT 1840.100 2.420 1840.360 2.680 ;
      LAYER met2 ;
        RECT 1481.210 1100.650 1481.490 1104.000 ;
        RECT 1481.210 1100.510 1482.420 1100.650 ;
        RECT 1481.210 1100.000 1481.490 1100.510 ;
        RECT 1482.280 73.770 1482.420 1100.510 ;
        RECT 1482.220 73.450 1482.480 73.770 ;
        RECT 1835.500 73.450 1835.760 73.770 ;
        RECT 1835.560 2.710 1835.700 73.450 ;
        RECT 1835.500 2.390 1835.760 2.710 ;
        RECT 1840.100 2.390 1840.360 2.710 ;
        RECT 1840.160 2.000 1840.300 2.390 ;
        RECT 1839.950 -4.000 1840.510 2.000 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1488.630 73.340 1488.950 73.400 ;
        RECT 1856.170 73.340 1856.490 73.400 ;
        RECT 1488.630 73.200 1856.490 73.340 ;
        RECT 1488.630 73.140 1488.950 73.200 ;
        RECT 1856.170 73.140 1856.490 73.200 ;
      LAYER via ;
        RECT 1488.660 73.140 1488.920 73.400 ;
        RECT 1856.200 73.140 1856.460 73.400 ;
      LAYER met2 ;
        RECT 1487.650 1100.650 1487.930 1104.000 ;
        RECT 1487.650 1100.510 1488.860 1100.650 ;
        RECT 1487.650 1100.000 1487.930 1100.510 ;
        RECT 1488.720 73.430 1488.860 1100.510 ;
        RECT 1488.660 73.110 1488.920 73.430 ;
        RECT 1856.200 73.110 1856.460 73.430 ;
        RECT 1856.260 2.450 1856.400 73.110 ;
        RECT 1856.260 2.310 1858.240 2.450 ;
        RECT 1858.100 2.000 1858.240 2.310 ;
        RECT 1857.890 -4.000 1858.450 2.000 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1496.065 724.625 1496.235 739.075 ;
        RECT 1496.065 620.925 1496.235 642.515 ;
        RECT 1496.065 511.105 1496.235 517.735 ;
      LAYER mcon ;
        RECT 1496.065 738.905 1496.235 739.075 ;
        RECT 1496.065 642.345 1496.235 642.515 ;
        RECT 1496.065 517.565 1496.235 517.735 ;
      LAYER met1 ;
        RECT 1495.990 739.060 1496.310 739.120 ;
        RECT 1495.795 738.920 1496.310 739.060 ;
        RECT 1495.990 738.860 1496.310 738.920 ;
        RECT 1495.990 724.780 1496.310 724.840 ;
        RECT 1495.795 724.640 1496.310 724.780 ;
        RECT 1495.990 724.580 1496.310 724.640 ;
        RECT 1495.990 642.500 1496.310 642.560 ;
        RECT 1495.795 642.360 1496.310 642.500 ;
        RECT 1495.990 642.300 1496.310 642.360 ;
        RECT 1495.990 621.080 1496.310 621.140 ;
        RECT 1495.795 620.940 1496.310 621.080 ;
        RECT 1495.990 620.880 1496.310 620.940 ;
        RECT 1495.990 517.720 1496.310 517.780 ;
        RECT 1495.795 517.580 1496.310 517.720 ;
        RECT 1495.990 517.520 1496.310 517.580 ;
        RECT 1495.990 511.260 1496.310 511.320 ;
        RECT 1495.795 511.120 1496.310 511.260 ;
        RECT 1495.990 511.060 1496.310 511.120 ;
        RECT 1494.610 510.580 1494.930 510.640 ;
        RECT 1495.990 510.580 1496.310 510.640 ;
        RECT 1494.610 510.440 1496.310 510.580 ;
        RECT 1494.610 510.380 1494.930 510.440 ;
        RECT 1495.990 510.380 1496.310 510.440 ;
        RECT 1495.530 73.000 1495.850 73.060 ;
        RECT 1875.950 73.000 1876.270 73.060 ;
        RECT 1495.530 72.860 1876.270 73.000 ;
        RECT 1495.530 72.800 1495.850 72.860 ;
        RECT 1875.950 72.800 1876.270 72.860 ;
      LAYER via ;
        RECT 1496.020 738.860 1496.280 739.120 ;
        RECT 1496.020 724.580 1496.280 724.840 ;
        RECT 1496.020 642.300 1496.280 642.560 ;
        RECT 1496.020 620.880 1496.280 621.140 ;
        RECT 1496.020 517.520 1496.280 517.780 ;
        RECT 1496.020 511.060 1496.280 511.320 ;
        RECT 1494.640 510.380 1494.900 510.640 ;
        RECT 1496.020 510.380 1496.280 510.640 ;
        RECT 1495.560 72.800 1495.820 73.060 ;
        RECT 1875.980 72.800 1876.240 73.060 ;
      LAYER met2 ;
        RECT 1493.630 1100.650 1493.910 1104.000 ;
        RECT 1493.630 1100.510 1495.300 1100.650 ;
        RECT 1493.630 1100.000 1493.910 1100.510 ;
        RECT 1495.160 1088.410 1495.300 1100.510 ;
        RECT 1495.160 1088.270 1496.220 1088.410 ;
        RECT 1496.080 980.290 1496.220 1088.270 ;
        RECT 1495.160 980.150 1496.220 980.290 ;
        RECT 1495.160 979.610 1495.300 980.150 ;
        RECT 1495.160 979.470 1495.760 979.610 ;
        RECT 1495.620 904.130 1495.760 979.470 ;
        RECT 1495.620 903.990 1496.220 904.130 ;
        RECT 1496.080 835.450 1496.220 903.990 ;
        RECT 1495.160 835.310 1496.220 835.450 ;
        RECT 1495.160 834.770 1495.300 835.310 ;
        RECT 1495.160 834.630 1495.760 834.770 ;
        RECT 1495.620 834.090 1495.760 834.630 ;
        RECT 1495.620 833.950 1496.220 834.090 ;
        RECT 1496.080 739.150 1496.220 833.950 ;
        RECT 1496.020 738.830 1496.280 739.150 ;
        RECT 1496.020 724.550 1496.280 724.870 ;
        RECT 1496.080 642.590 1496.220 724.550 ;
        RECT 1496.020 642.270 1496.280 642.590 ;
        RECT 1496.020 620.850 1496.280 621.170 ;
        RECT 1496.080 517.810 1496.220 620.850 ;
        RECT 1496.020 517.490 1496.280 517.810 ;
        RECT 1496.020 511.030 1496.280 511.350 ;
        RECT 1496.080 510.670 1496.220 511.030 ;
        RECT 1494.640 510.350 1494.900 510.670 ;
        RECT 1496.020 510.350 1496.280 510.670 ;
        RECT 1494.700 435.045 1494.840 510.350 ;
        RECT 1494.630 434.675 1494.910 435.045 ;
        RECT 1496.010 434.675 1496.290 435.045 ;
        RECT 1496.080 158.850 1496.220 434.675 ;
        RECT 1495.620 158.710 1496.220 158.850 ;
        RECT 1495.620 73.090 1495.760 158.710 ;
        RECT 1495.560 72.770 1495.820 73.090 ;
        RECT 1875.980 72.770 1876.240 73.090 ;
        RECT 1876.040 2.000 1876.180 72.770 ;
        RECT 1875.830 -4.000 1876.390 2.000 ;
      LAYER via2 ;
        RECT 1494.630 434.720 1494.910 435.000 ;
        RECT 1496.010 434.720 1496.290 435.000 ;
      LAYER met3 ;
        RECT 1494.605 435.010 1494.935 435.025 ;
        RECT 1495.985 435.010 1496.315 435.025 ;
        RECT 1494.605 434.710 1496.315 435.010 ;
        RECT 1494.605 434.695 1494.935 434.710 ;
        RECT 1495.985 434.695 1496.315 434.710 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1104.990 1052.200 1105.310 1052.260 ;
        RECT 1106.830 1052.200 1107.150 1052.260 ;
        RECT 1104.990 1052.060 1107.150 1052.200 ;
        RECT 1104.990 1052.000 1105.310 1052.060 ;
        RECT 1106.830 1052.000 1107.150 1052.060 ;
        RECT 752.170 28.800 752.490 28.860 ;
        RECT 1104.990 28.800 1105.310 28.860 ;
        RECT 752.170 28.660 1105.310 28.800 ;
        RECT 752.170 28.600 752.490 28.660 ;
        RECT 1104.990 28.600 1105.310 28.660 ;
      LAYER via ;
        RECT 1105.020 1052.000 1105.280 1052.260 ;
        RECT 1106.860 1052.000 1107.120 1052.260 ;
        RECT 752.200 28.600 752.460 28.860 ;
        RECT 1105.020 28.600 1105.280 28.860 ;
      LAYER met2 ;
        RECT 1108.150 1100.650 1108.430 1104.000 ;
        RECT 1106.920 1100.510 1108.430 1100.650 ;
        RECT 1106.920 1052.290 1107.060 1100.510 ;
        RECT 1108.150 1100.000 1108.430 1100.510 ;
        RECT 1105.020 1051.970 1105.280 1052.290 ;
        RECT 1106.860 1051.970 1107.120 1052.290 ;
        RECT 1105.080 28.890 1105.220 1051.970 ;
        RECT 752.200 28.570 752.460 28.890 ;
        RECT 1105.020 28.570 1105.280 28.890 ;
        RECT 752.260 2.000 752.400 28.570 ;
        RECT 752.050 -4.000 752.610 2.000 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1502.505 724.625 1502.675 739.075 ;
        RECT 1502.505 620.925 1502.675 642.515 ;
        RECT 1502.505 517.565 1502.675 545.955 ;
      LAYER mcon ;
        RECT 1502.505 738.905 1502.675 739.075 ;
        RECT 1502.505 642.345 1502.675 642.515 ;
        RECT 1502.505 545.785 1502.675 545.955 ;
      LAYER met1 ;
        RECT 1499.670 1062.740 1499.990 1062.800 ;
        RECT 1502.430 1062.740 1502.750 1062.800 ;
        RECT 1499.670 1062.600 1502.750 1062.740 ;
        RECT 1499.670 1062.540 1499.990 1062.600 ;
        RECT 1502.430 1062.540 1502.750 1062.600 ;
        RECT 1502.430 739.060 1502.750 739.120 ;
        RECT 1502.235 738.920 1502.750 739.060 ;
        RECT 1502.430 738.860 1502.750 738.920 ;
        RECT 1502.430 724.780 1502.750 724.840 ;
        RECT 1502.235 724.640 1502.750 724.780 ;
        RECT 1502.430 724.580 1502.750 724.640 ;
        RECT 1502.430 642.500 1502.750 642.560 ;
        RECT 1502.235 642.360 1502.750 642.500 ;
        RECT 1502.430 642.300 1502.750 642.360 ;
        RECT 1502.430 621.080 1502.750 621.140 ;
        RECT 1502.235 620.940 1502.750 621.080 ;
        RECT 1502.430 620.880 1502.750 620.940 ;
        RECT 1502.430 545.940 1502.750 546.000 ;
        RECT 1502.235 545.800 1502.750 545.940 ;
        RECT 1502.430 545.740 1502.750 545.800 ;
        RECT 1502.430 517.720 1502.750 517.780 ;
        RECT 1502.235 517.580 1502.750 517.720 ;
        RECT 1502.430 517.520 1502.750 517.580 ;
        RECT 1501.970 72.660 1502.290 72.720 ;
        RECT 1890.670 72.660 1890.990 72.720 ;
        RECT 1501.970 72.520 1890.990 72.660 ;
        RECT 1501.970 72.460 1502.290 72.520 ;
        RECT 1890.670 72.460 1890.990 72.520 ;
      LAYER via ;
        RECT 1499.700 1062.540 1499.960 1062.800 ;
        RECT 1502.460 1062.540 1502.720 1062.800 ;
        RECT 1502.460 738.860 1502.720 739.120 ;
        RECT 1502.460 724.580 1502.720 724.840 ;
        RECT 1502.460 642.300 1502.720 642.560 ;
        RECT 1502.460 620.880 1502.720 621.140 ;
        RECT 1502.460 545.740 1502.720 546.000 ;
        RECT 1502.460 517.520 1502.720 517.780 ;
        RECT 1502.000 72.460 1502.260 72.720 ;
        RECT 1890.700 72.460 1890.960 72.720 ;
      LAYER met2 ;
        RECT 1499.610 1100.580 1499.890 1104.000 ;
        RECT 1499.610 1100.000 1499.900 1100.580 ;
        RECT 1499.760 1062.830 1499.900 1100.000 ;
        RECT 1499.700 1062.510 1499.960 1062.830 ;
        RECT 1502.460 1062.510 1502.720 1062.830 ;
        RECT 1502.520 980.290 1502.660 1062.510 ;
        RECT 1501.600 980.150 1502.660 980.290 ;
        RECT 1501.600 979.610 1501.740 980.150 ;
        RECT 1501.600 979.470 1502.200 979.610 ;
        RECT 1502.060 904.130 1502.200 979.470 ;
        RECT 1502.060 903.990 1502.660 904.130 ;
        RECT 1502.520 835.450 1502.660 903.990 ;
        RECT 1501.600 835.310 1502.660 835.450 ;
        RECT 1501.600 834.770 1501.740 835.310 ;
        RECT 1501.600 834.630 1502.200 834.770 ;
        RECT 1502.060 834.090 1502.200 834.630 ;
        RECT 1502.060 833.950 1502.660 834.090 ;
        RECT 1502.520 739.150 1502.660 833.950 ;
        RECT 1502.460 738.830 1502.720 739.150 ;
        RECT 1502.460 724.550 1502.720 724.870 ;
        RECT 1502.520 642.590 1502.660 724.550 ;
        RECT 1502.460 642.270 1502.720 642.590 ;
        RECT 1502.460 620.850 1502.720 621.170 ;
        RECT 1502.520 546.030 1502.660 620.850 ;
        RECT 1502.460 545.710 1502.720 546.030 ;
        RECT 1502.460 517.490 1502.720 517.810 ;
        RECT 1502.520 158.850 1502.660 517.490 ;
        RECT 1502.060 158.710 1502.660 158.850 ;
        RECT 1502.060 72.750 1502.200 158.710 ;
        RECT 1502.000 72.430 1502.260 72.750 ;
        RECT 1890.700 72.430 1890.960 72.750 ;
        RECT 1890.760 2.450 1890.900 72.430 ;
        RECT 1890.760 2.310 1894.120 2.450 ;
        RECT 1893.980 2.000 1894.120 2.310 ;
        RECT 1893.770 -4.000 1894.330 2.000 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1661.665 1089.105 1661.835 1090.295 ;
      LAYER mcon ;
        RECT 1661.665 1090.125 1661.835 1090.295 ;
      LAYER met1 ;
        RECT 1661.605 1090.280 1661.895 1090.325 ;
        RECT 1673.090 1090.280 1673.410 1090.340 ;
        RECT 1661.605 1090.140 1673.410 1090.280 ;
        RECT 1661.605 1090.095 1661.895 1090.140 ;
        RECT 1673.090 1090.080 1673.410 1090.140 ;
        RECT 1506.110 1089.260 1506.430 1089.320 ;
        RECT 1661.605 1089.260 1661.895 1089.305 ;
        RECT 1506.110 1089.120 1661.895 1089.260 ;
        RECT 1506.110 1089.060 1506.430 1089.120 ;
        RECT 1661.605 1089.075 1661.895 1089.120 ;
        RECT 1673.090 14.520 1673.410 14.580 ;
        RECT 1911.370 14.520 1911.690 14.580 ;
        RECT 1673.090 14.380 1911.690 14.520 ;
        RECT 1673.090 14.320 1673.410 14.380 ;
        RECT 1911.370 14.320 1911.690 14.380 ;
      LAYER via ;
        RECT 1673.120 1090.080 1673.380 1090.340 ;
        RECT 1506.140 1089.060 1506.400 1089.320 ;
        RECT 1673.120 14.320 1673.380 14.580 ;
        RECT 1911.400 14.320 1911.660 14.580 ;
      LAYER met2 ;
        RECT 1506.050 1100.580 1506.330 1104.000 ;
        RECT 1506.050 1100.000 1506.340 1100.580 ;
        RECT 1506.200 1089.350 1506.340 1100.000 ;
        RECT 1673.120 1090.050 1673.380 1090.370 ;
        RECT 1506.140 1089.030 1506.400 1089.350 ;
        RECT 1673.180 14.610 1673.320 1090.050 ;
        RECT 1673.120 14.290 1673.380 14.610 ;
        RECT 1911.400 14.290 1911.660 14.610 ;
        RECT 1911.460 14.010 1911.600 14.290 ;
        RECT 1911.460 13.870 1912.060 14.010 ;
        RECT 1911.920 2.000 1912.060 13.870 ;
        RECT 1911.710 -4.000 1912.270 2.000 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1536.085 1084.005 1536.255 1085.195 ;
      LAYER mcon ;
        RECT 1536.085 1085.025 1536.255 1085.195 ;
      LAYER met1 ;
        RECT 1512.090 1085.180 1512.410 1085.240 ;
        RECT 1536.025 1085.180 1536.315 1085.225 ;
        RECT 1512.090 1085.040 1536.315 1085.180 ;
        RECT 1512.090 1084.980 1512.410 1085.040 ;
        RECT 1536.025 1084.995 1536.315 1085.040 ;
        RECT 1536.025 1084.160 1536.315 1084.205 ;
        RECT 1925.170 1084.160 1925.490 1084.220 ;
        RECT 1536.025 1084.020 1925.490 1084.160 ;
        RECT 1536.025 1083.975 1536.315 1084.020 ;
        RECT 1925.170 1083.960 1925.490 1084.020 ;
        RECT 1925.170 2.620 1925.490 2.680 ;
        RECT 1929.310 2.620 1929.630 2.680 ;
        RECT 1925.170 2.480 1929.630 2.620 ;
        RECT 1925.170 2.420 1925.490 2.480 ;
        RECT 1929.310 2.420 1929.630 2.480 ;
      LAYER via ;
        RECT 1512.120 1084.980 1512.380 1085.240 ;
        RECT 1925.200 1083.960 1925.460 1084.220 ;
        RECT 1925.200 2.420 1925.460 2.680 ;
        RECT 1929.340 2.420 1929.600 2.680 ;
      LAYER met2 ;
        RECT 1512.030 1100.580 1512.310 1104.000 ;
        RECT 1512.030 1100.000 1512.320 1100.580 ;
        RECT 1512.180 1085.270 1512.320 1100.000 ;
        RECT 1512.120 1084.950 1512.380 1085.270 ;
        RECT 1925.200 1083.930 1925.460 1084.250 ;
        RECT 1925.260 2.710 1925.400 1083.930 ;
        RECT 1925.200 2.390 1925.460 2.710 ;
        RECT 1929.340 2.390 1929.600 2.710 ;
        RECT 1929.400 2.000 1929.540 2.390 ;
        RECT 1929.190 -4.000 1929.750 2.000 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1703.910 1089.260 1704.230 1089.320 ;
        RECT 1727.830 1089.260 1728.150 1089.320 ;
        RECT 1703.910 1089.120 1728.150 1089.260 ;
        RECT 1703.910 1089.060 1704.230 1089.120 ;
        RECT 1727.830 1089.060 1728.150 1089.120 ;
        RECT 1518.070 1088.580 1518.390 1088.640 ;
        RECT 1656.530 1088.580 1656.850 1088.640 ;
        RECT 1518.070 1088.440 1656.850 1088.580 ;
        RECT 1518.070 1088.380 1518.390 1088.440 ;
        RECT 1656.530 1088.380 1656.850 1088.440 ;
        RECT 1728.750 14.180 1729.070 14.240 ;
        RECT 1947.250 14.180 1947.570 14.240 ;
        RECT 1728.750 14.040 1947.570 14.180 ;
        RECT 1728.750 13.980 1729.070 14.040 ;
        RECT 1947.250 13.980 1947.570 14.040 ;
      LAYER via ;
        RECT 1703.940 1089.060 1704.200 1089.320 ;
        RECT 1727.860 1089.060 1728.120 1089.320 ;
        RECT 1518.100 1088.380 1518.360 1088.640 ;
        RECT 1656.560 1088.380 1656.820 1088.640 ;
        RECT 1728.780 13.980 1729.040 14.240 ;
        RECT 1947.280 13.980 1947.540 14.240 ;
      LAYER met2 ;
        RECT 1518.010 1100.580 1518.290 1104.000 ;
        RECT 1518.010 1100.000 1518.300 1100.580 ;
        RECT 1518.160 1088.670 1518.300 1100.000 ;
        RECT 1703.940 1089.205 1704.200 1089.350 ;
        RECT 1656.550 1088.835 1656.830 1089.205 ;
        RECT 1703.930 1088.835 1704.210 1089.205 ;
        RECT 1727.860 1089.030 1728.120 1089.350 ;
        RECT 1656.620 1088.670 1656.760 1088.835 ;
        RECT 1518.100 1088.350 1518.360 1088.670 ;
        RECT 1656.560 1088.350 1656.820 1088.670 ;
        RECT 1727.920 1088.410 1728.060 1089.030 ;
        RECT 1727.920 1088.270 1728.980 1088.410 ;
        RECT 1728.840 14.270 1728.980 1088.270 ;
        RECT 1728.780 13.950 1729.040 14.270 ;
        RECT 1947.280 13.950 1947.540 14.270 ;
        RECT 1947.340 2.000 1947.480 13.950 ;
        RECT 1947.130 -4.000 1947.690 2.000 ;
      LAYER via2 ;
        RECT 1656.550 1088.880 1656.830 1089.160 ;
        RECT 1703.930 1088.880 1704.210 1089.160 ;
      LAYER met3 ;
        RECT 1656.525 1089.170 1656.855 1089.185 ;
        RECT 1703.905 1089.170 1704.235 1089.185 ;
        RECT 1656.525 1088.870 1704.235 1089.170 ;
        RECT 1656.525 1088.855 1656.855 1088.870 ;
        RECT 1703.905 1088.855 1704.235 1088.870 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1542.065 1084.345 1543.615 1084.515 ;
      LAYER mcon ;
        RECT 1543.445 1084.345 1543.615 1084.515 ;
      LAYER met1 ;
        RECT 1524.510 1084.500 1524.830 1084.560 ;
        RECT 1542.005 1084.500 1542.295 1084.545 ;
        RECT 1524.510 1084.360 1542.295 1084.500 ;
        RECT 1524.510 1084.300 1524.830 1084.360 ;
        RECT 1542.005 1084.315 1542.295 1084.360 ;
        RECT 1543.385 1084.500 1543.675 1084.545 ;
        RECT 1959.670 1084.500 1959.990 1084.560 ;
        RECT 1543.385 1084.360 1959.990 1084.500 ;
        RECT 1543.385 1084.315 1543.675 1084.360 ;
        RECT 1959.670 1084.300 1959.990 1084.360 ;
        RECT 1959.670 2.620 1959.990 2.680 ;
        RECT 1965.190 2.620 1965.510 2.680 ;
        RECT 1959.670 2.480 1965.510 2.620 ;
        RECT 1959.670 2.420 1959.990 2.480 ;
        RECT 1965.190 2.420 1965.510 2.480 ;
      LAYER via ;
        RECT 1524.540 1084.300 1524.800 1084.560 ;
        RECT 1959.700 1084.300 1959.960 1084.560 ;
        RECT 1959.700 2.420 1959.960 2.680 ;
        RECT 1965.220 2.420 1965.480 2.680 ;
      LAYER met2 ;
        RECT 1524.450 1100.580 1524.730 1104.000 ;
        RECT 1524.450 1100.000 1524.740 1100.580 ;
        RECT 1524.600 1084.590 1524.740 1100.000 ;
        RECT 1524.540 1084.270 1524.800 1084.590 ;
        RECT 1959.700 1084.270 1959.960 1084.590 ;
        RECT 1959.760 2.710 1959.900 1084.270 ;
        RECT 1959.700 2.390 1959.960 2.710 ;
        RECT 1965.220 2.390 1965.480 2.710 ;
        RECT 1965.280 2.000 1965.420 2.390 ;
        RECT 1965.070 -4.000 1965.630 2.000 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1530.490 1087.220 1530.810 1087.280 ;
        RECT 1610.990 1087.220 1611.310 1087.280 ;
        RECT 1530.490 1087.080 1611.310 1087.220 ;
        RECT 1530.490 1087.020 1530.810 1087.080 ;
        RECT 1610.990 1087.020 1611.310 1087.080 ;
        RECT 1610.990 14.860 1611.310 14.920 ;
        RECT 1983.130 14.860 1983.450 14.920 ;
        RECT 1610.990 14.720 1983.450 14.860 ;
        RECT 1610.990 14.660 1611.310 14.720 ;
        RECT 1983.130 14.660 1983.450 14.720 ;
      LAYER via ;
        RECT 1530.520 1087.020 1530.780 1087.280 ;
        RECT 1611.020 1087.020 1611.280 1087.280 ;
        RECT 1611.020 14.660 1611.280 14.920 ;
        RECT 1983.160 14.660 1983.420 14.920 ;
      LAYER met2 ;
        RECT 1530.430 1100.580 1530.710 1104.000 ;
        RECT 1530.430 1100.000 1530.720 1100.580 ;
        RECT 1530.580 1087.310 1530.720 1100.000 ;
        RECT 1530.520 1086.990 1530.780 1087.310 ;
        RECT 1611.020 1086.990 1611.280 1087.310 ;
        RECT 1611.080 14.950 1611.220 1086.990 ;
        RECT 1611.020 14.630 1611.280 14.950 ;
        RECT 1983.160 14.630 1983.420 14.950 ;
        RECT 1983.220 2.000 1983.360 14.630 ;
        RECT 1983.010 -4.000 1983.570 2.000 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1536.470 1085.180 1536.790 1085.240 ;
        RECT 1536.470 1085.040 1560.160 1085.180 ;
        RECT 1536.470 1084.980 1536.790 1085.040 ;
        RECT 1560.020 1084.840 1560.160 1085.040 ;
        RECT 2001.070 1084.840 2001.390 1084.900 ;
        RECT 1560.020 1084.700 2001.390 1084.840 ;
        RECT 2001.070 1084.640 2001.390 1084.700 ;
      LAYER via ;
        RECT 1536.500 1084.980 1536.760 1085.240 ;
        RECT 2001.100 1084.640 2001.360 1084.900 ;
      LAYER met2 ;
        RECT 1536.410 1100.580 1536.690 1104.000 ;
        RECT 1536.410 1100.000 1536.700 1100.580 ;
        RECT 1536.560 1085.270 1536.700 1100.000 ;
        RECT 1536.500 1084.950 1536.760 1085.270 ;
        RECT 2001.100 1084.610 2001.360 1084.930 ;
        RECT 2001.160 2.000 2001.300 1084.610 ;
        RECT 2000.950 -4.000 2001.510 2.000 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1559.545 1083.665 1559.715 1084.855 ;
      LAYER mcon ;
        RECT 1559.545 1084.685 1559.715 1084.855 ;
      LAYER met1 ;
        RECT 1542.910 1084.840 1543.230 1084.900 ;
        RECT 1559.485 1084.840 1559.775 1084.885 ;
        RECT 1542.910 1084.700 1559.775 1084.840 ;
        RECT 1542.910 1084.640 1543.230 1084.700 ;
        RECT 1559.485 1084.655 1559.775 1084.700 ;
        RECT 1559.485 1083.820 1559.775 1083.865 ;
        RECT 1559.485 1083.680 1607.540 1083.820 ;
        RECT 1559.485 1083.635 1559.775 1083.680 ;
        RECT 1607.400 1083.480 1607.540 1083.680 ;
        RECT 1617.890 1083.480 1618.210 1083.540 ;
        RECT 1607.400 1083.340 1618.210 1083.480 ;
        RECT 1617.890 1083.280 1618.210 1083.340 ;
        RECT 1617.890 15.540 1618.210 15.600 ;
        RECT 2018.550 15.540 2018.870 15.600 ;
        RECT 1617.890 15.400 2018.870 15.540 ;
        RECT 1617.890 15.340 1618.210 15.400 ;
        RECT 2018.550 15.340 2018.870 15.400 ;
      LAYER via ;
        RECT 1542.940 1084.640 1543.200 1084.900 ;
        RECT 1617.920 1083.280 1618.180 1083.540 ;
        RECT 1617.920 15.340 1618.180 15.600 ;
        RECT 2018.580 15.340 2018.840 15.600 ;
      LAYER met2 ;
        RECT 1542.850 1100.580 1543.130 1104.000 ;
        RECT 1542.850 1100.000 1543.140 1100.580 ;
        RECT 1543.000 1084.930 1543.140 1100.000 ;
        RECT 1542.940 1084.610 1543.200 1084.930 ;
        RECT 1617.920 1083.250 1618.180 1083.570 ;
        RECT 1617.980 15.630 1618.120 1083.250 ;
        RECT 1617.920 15.310 1618.180 15.630 ;
        RECT 2018.580 15.310 2018.840 15.630 ;
        RECT 2018.640 2.000 2018.780 15.310 ;
        RECT 2018.430 -4.000 2018.990 2.000 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1599.565 1085.025 1599.735 1086.215 ;
      LAYER mcon ;
        RECT 1599.565 1086.045 1599.735 1086.215 ;
      LAYER met1 ;
        RECT 1599.505 1086.200 1599.795 1086.245 ;
        RECT 1573.360 1086.060 1599.795 1086.200 ;
        RECT 1550.270 1085.860 1550.590 1085.920 ;
        RECT 1573.360 1085.860 1573.500 1086.060 ;
        RECT 1599.505 1086.015 1599.795 1086.060 ;
        RECT 1550.270 1085.720 1573.500 1085.860 ;
        RECT 1550.270 1085.660 1550.590 1085.720 ;
        RECT 1599.505 1085.180 1599.795 1085.225 ;
        RECT 2035.570 1085.180 2035.890 1085.240 ;
        RECT 1599.505 1085.040 2035.890 1085.180 ;
        RECT 1599.505 1084.995 1599.795 1085.040 ;
        RECT 2035.570 1084.980 2035.890 1085.040 ;
      LAYER via ;
        RECT 1550.300 1085.660 1550.560 1085.920 ;
        RECT 2035.600 1084.980 2035.860 1085.240 ;
      LAYER met2 ;
        RECT 1548.830 1100.650 1549.110 1104.000 ;
        RECT 1548.830 1100.510 1550.500 1100.650 ;
        RECT 1548.830 1100.000 1549.110 1100.510 ;
        RECT 1550.360 1085.950 1550.500 1100.510 ;
        RECT 1550.300 1085.630 1550.560 1085.950 ;
        RECT 2035.600 1084.950 2035.860 1085.270 ;
        RECT 2035.660 16.730 2035.800 1084.950 ;
        RECT 2035.660 16.590 2036.720 16.730 ;
        RECT 2036.580 2.000 2036.720 16.590 ;
        RECT 2036.370 -4.000 2036.930 2.000 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1554.870 1086.880 1555.190 1086.940 ;
        RECT 1554.870 1086.740 1563.380 1086.880 ;
        RECT 1554.870 1086.680 1555.190 1086.740 ;
        RECT 1563.240 1086.540 1563.380 1086.740 ;
        RECT 1631.690 1086.540 1632.010 1086.600 ;
        RECT 1563.240 1086.400 1632.010 1086.540 ;
        RECT 1631.690 1086.340 1632.010 1086.400 ;
        RECT 1631.690 15.880 1632.010 15.940 ;
        RECT 2054.430 15.880 2054.750 15.940 ;
        RECT 1631.690 15.740 2054.750 15.880 ;
        RECT 1631.690 15.680 1632.010 15.740 ;
        RECT 2054.430 15.680 2054.750 15.740 ;
      LAYER via ;
        RECT 1554.900 1086.680 1555.160 1086.940 ;
        RECT 1631.720 1086.340 1631.980 1086.600 ;
        RECT 1631.720 15.680 1631.980 15.940 ;
        RECT 2054.460 15.680 2054.720 15.940 ;
      LAYER met2 ;
        RECT 1554.810 1100.580 1555.090 1104.000 ;
        RECT 1554.810 1100.000 1555.100 1100.580 ;
        RECT 1554.960 1086.970 1555.100 1100.000 ;
        RECT 1554.900 1086.650 1555.160 1086.970 ;
        RECT 1631.720 1086.310 1631.980 1086.630 ;
        RECT 1631.780 15.970 1631.920 1086.310 ;
        RECT 1631.720 15.650 1631.980 15.970 ;
        RECT 2054.460 15.650 2054.720 15.970 ;
        RECT 2054.520 2.000 2054.660 15.650 ;
        RECT 2054.310 -4.000 2054.870 2.000 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1111.430 1052.200 1111.750 1052.260 ;
        RECT 1112.350 1052.200 1112.670 1052.260 ;
        RECT 1111.430 1052.060 1112.670 1052.200 ;
        RECT 1111.430 1052.000 1111.750 1052.060 ;
        RECT 1112.350 1052.000 1112.670 1052.060 ;
        RECT 769.650 35.600 769.970 35.660 ;
        RECT 1111.430 35.600 1111.750 35.660 ;
        RECT 769.650 35.460 1111.750 35.600 ;
        RECT 769.650 35.400 769.970 35.460 ;
        RECT 1111.430 35.400 1111.750 35.460 ;
      LAYER via ;
        RECT 1111.460 1052.000 1111.720 1052.260 ;
        RECT 1112.380 1052.000 1112.640 1052.260 ;
        RECT 769.680 35.400 769.940 35.660 ;
        RECT 1111.460 35.400 1111.720 35.660 ;
      LAYER met2 ;
        RECT 1114.130 1100.650 1114.410 1104.000 ;
        RECT 1112.440 1100.510 1114.410 1100.650 ;
        RECT 1112.440 1052.290 1112.580 1100.510 ;
        RECT 1114.130 1100.000 1114.410 1100.510 ;
        RECT 1111.460 1051.970 1111.720 1052.290 ;
        RECT 1112.380 1051.970 1112.640 1052.290 ;
        RECT 1111.520 35.690 1111.660 1051.970 ;
        RECT 769.680 35.370 769.940 35.690 ;
        RECT 1111.460 35.370 1111.720 35.690 ;
        RECT 769.740 2.000 769.880 35.370 ;
        RECT 769.530 -4.000 770.090 2.000 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2070.070 1085.520 2070.390 1085.580 ;
        RECT 1587.160 1085.380 2070.390 1085.520 ;
        RECT 1560.850 1085.180 1561.170 1085.240 ;
        RECT 1587.160 1085.180 1587.300 1085.380 ;
        RECT 2070.070 1085.320 2070.390 1085.380 ;
        RECT 1560.850 1085.040 1587.300 1085.180 ;
        RECT 1560.850 1084.980 1561.170 1085.040 ;
      LAYER via ;
        RECT 1560.880 1084.980 1561.140 1085.240 ;
        RECT 2070.100 1085.320 2070.360 1085.580 ;
      LAYER met2 ;
        RECT 1560.790 1100.580 1561.070 1104.000 ;
        RECT 1560.790 1100.000 1561.080 1100.580 ;
        RECT 1560.940 1085.270 1561.080 1100.000 ;
        RECT 2070.100 1085.290 2070.360 1085.610 ;
        RECT 1560.880 1084.950 1561.140 1085.270 ;
        RECT 2070.160 16.730 2070.300 1085.290 ;
        RECT 2070.160 16.590 2072.600 16.730 ;
        RECT 2072.460 2.000 2072.600 16.590 ;
        RECT 2072.250 -4.000 2072.810 2.000 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1567.290 1086.880 1567.610 1086.940 ;
        RECT 1638.590 1086.880 1638.910 1086.940 ;
        RECT 1567.290 1086.740 1638.910 1086.880 ;
        RECT 1567.290 1086.680 1567.610 1086.740 ;
        RECT 1638.590 1086.680 1638.910 1086.740 ;
        RECT 1638.590 16.560 1638.910 16.620 ;
        RECT 2089.850 16.560 2090.170 16.620 ;
        RECT 1638.590 16.420 2090.170 16.560 ;
        RECT 1638.590 16.360 1638.910 16.420 ;
        RECT 2089.850 16.360 2090.170 16.420 ;
      LAYER via ;
        RECT 1567.320 1086.680 1567.580 1086.940 ;
        RECT 1638.620 1086.680 1638.880 1086.940 ;
        RECT 1638.620 16.360 1638.880 16.620 ;
        RECT 2089.880 16.360 2090.140 16.620 ;
      LAYER met2 ;
        RECT 1567.230 1100.580 1567.510 1104.000 ;
        RECT 1567.230 1100.000 1567.520 1100.580 ;
        RECT 1567.380 1086.970 1567.520 1100.000 ;
        RECT 1567.320 1086.650 1567.580 1086.970 ;
        RECT 1638.620 1086.650 1638.880 1086.970 ;
        RECT 1638.680 16.650 1638.820 1086.650 ;
        RECT 1638.620 16.330 1638.880 16.650 ;
        RECT 2089.880 16.330 2090.140 16.650 ;
        RECT 2089.940 2.000 2090.080 16.330 ;
        RECT 2089.730 -4.000 2090.290 2.000 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1574.190 1085.860 1574.510 1085.920 ;
        RECT 2104.570 1085.860 2104.890 1085.920 ;
        RECT 1574.190 1085.720 2104.890 1085.860 ;
        RECT 1574.190 1085.660 1574.510 1085.720 ;
        RECT 2104.570 1085.660 2104.890 1085.720 ;
      LAYER via ;
        RECT 1574.220 1085.660 1574.480 1085.920 ;
        RECT 2104.600 1085.660 2104.860 1085.920 ;
      LAYER met2 ;
        RECT 1573.210 1100.580 1573.490 1104.000 ;
        RECT 1573.210 1100.000 1573.500 1100.580 ;
        RECT 1573.360 1085.690 1573.500 1100.000 ;
        RECT 1574.220 1085.690 1574.480 1085.950 ;
        RECT 1573.360 1085.630 1574.480 1085.690 ;
        RECT 2104.600 1085.630 2104.860 1085.950 ;
        RECT 1573.360 1085.550 1574.420 1085.630 ;
        RECT 2104.660 16.730 2104.800 1085.630 ;
        RECT 2104.660 16.590 2108.020 16.730 ;
        RECT 2107.880 2.000 2108.020 16.590 ;
        RECT 2107.670 -4.000 2108.230 2.000 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1700.690 1090.620 1701.010 1090.680 ;
        RECT 1657.080 1090.480 1701.010 1090.620 ;
        RECT 1657.080 1090.280 1657.220 1090.480 ;
        RECT 1700.690 1090.420 1701.010 1090.480 ;
        RECT 1656.160 1090.140 1657.220 1090.280 ;
        RECT 1579.250 1089.940 1579.570 1090.000 ;
        RECT 1656.160 1089.940 1656.300 1090.140 ;
        RECT 1579.250 1089.800 1656.300 1089.940 ;
        RECT 1579.250 1089.740 1579.570 1089.800 ;
        RECT 1700.690 16.220 1701.010 16.280 ;
        RECT 2125.730 16.220 2126.050 16.280 ;
        RECT 1700.690 16.080 2126.050 16.220 ;
        RECT 1700.690 16.020 1701.010 16.080 ;
        RECT 2125.730 16.020 2126.050 16.080 ;
      LAYER via ;
        RECT 1700.720 1090.420 1700.980 1090.680 ;
        RECT 1579.280 1089.740 1579.540 1090.000 ;
        RECT 1700.720 16.020 1700.980 16.280 ;
        RECT 2125.760 16.020 2126.020 16.280 ;
      LAYER met2 ;
        RECT 1579.190 1100.580 1579.470 1104.000 ;
        RECT 1579.190 1100.000 1579.480 1100.580 ;
        RECT 1579.340 1090.030 1579.480 1100.000 ;
        RECT 1700.720 1090.390 1700.980 1090.710 ;
        RECT 1579.280 1089.710 1579.540 1090.030 ;
        RECT 1700.780 16.310 1700.920 1090.390 ;
        RECT 1700.720 15.990 1700.980 16.310 ;
        RECT 2125.760 15.990 2126.020 16.310 ;
        RECT 2125.820 2.000 2125.960 15.990 ;
        RECT 2125.610 -4.000 2126.170 2.000 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1600.025 1086.045 1600.195 1087.575 ;
      LAYER mcon ;
        RECT 1600.025 1087.405 1600.195 1087.575 ;
      LAYER met1 ;
        RECT 1585.690 1087.560 1586.010 1087.620 ;
        RECT 1599.965 1087.560 1600.255 1087.605 ;
        RECT 1585.690 1087.420 1600.255 1087.560 ;
        RECT 1585.690 1087.360 1586.010 1087.420 ;
        RECT 1599.965 1087.375 1600.255 1087.420 ;
        RECT 1599.965 1086.200 1600.255 1086.245 ;
        RECT 2139.070 1086.200 2139.390 1086.260 ;
        RECT 1599.965 1086.060 2139.390 1086.200 ;
        RECT 1599.965 1086.015 1600.255 1086.060 ;
        RECT 2139.070 1086.000 2139.390 1086.060 ;
      LAYER via ;
        RECT 1585.720 1087.360 1585.980 1087.620 ;
        RECT 2139.100 1086.000 2139.360 1086.260 ;
      LAYER met2 ;
        RECT 1585.630 1100.580 1585.910 1104.000 ;
        RECT 1585.630 1100.000 1585.920 1100.580 ;
        RECT 1585.780 1087.650 1585.920 1100.000 ;
        RECT 1585.720 1087.330 1585.980 1087.650 ;
        RECT 2139.100 1085.970 2139.360 1086.290 ;
        RECT 2139.160 16.730 2139.300 1085.970 ;
        RECT 2139.160 16.590 2143.900 16.730 ;
        RECT 2143.760 2.000 2143.900 16.590 ;
        RECT 2143.550 -4.000 2144.110 2.000 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1752.745 1088.765 1752.915 1089.615 ;
        RECT 1824.965 15.045 1825.135 17.255 ;
      LAYER mcon ;
        RECT 1752.745 1089.445 1752.915 1089.615 ;
        RECT 1824.965 17.085 1825.135 17.255 ;
      LAYER met1 ;
        RECT 1752.685 1089.600 1752.975 1089.645 ;
        RECT 1790.390 1089.600 1790.710 1089.660 ;
        RECT 1752.685 1089.460 1790.710 1089.600 ;
        RECT 1752.685 1089.415 1752.975 1089.460 ;
        RECT 1790.390 1089.400 1790.710 1089.460 ;
        RECT 1591.670 1088.920 1591.990 1088.980 ;
        RECT 1752.685 1088.920 1752.975 1088.965 ;
        RECT 1591.670 1088.780 1752.975 1088.920 ;
        RECT 1591.670 1088.720 1591.990 1088.780 ;
        RECT 1752.685 1088.735 1752.975 1088.780 ;
        RECT 1790.390 17.240 1790.710 17.300 ;
        RECT 1824.905 17.240 1825.195 17.285 ;
        RECT 1790.390 17.100 1825.195 17.240 ;
        RECT 1790.390 17.040 1790.710 17.100 ;
        RECT 1824.905 17.055 1825.195 17.100 ;
        RECT 1824.905 15.200 1825.195 15.245 ;
        RECT 2161.610 15.200 2161.930 15.260 ;
        RECT 1824.905 15.060 2161.930 15.200 ;
        RECT 1824.905 15.015 1825.195 15.060 ;
        RECT 2161.610 15.000 2161.930 15.060 ;
      LAYER via ;
        RECT 1790.420 1089.400 1790.680 1089.660 ;
        RECT 1591.700 1088.720 1591.960 1088.980 ;
        RECT 1790.420 17.040 1790.680 17.300 ;
        RECT 2161.640 15.000 2161.900 15.260 ;
      LAYER met2 ;
        RECT 1591.610 1100.580 1591.890 1104.000 ;
        RECT 1591.610 1100.000 1591.900 1100.580 ;
        RECT 1591.760 1089.010 1591.900 1100.000 ;
        RECT 1790.420 1089.370 1790.680 1089.690 ;
        RECT 1591.700 1088.690 1591.960 1089.010 ;
        RECT 1790.480 17.330 1790.620 1089.370 ;
        RECT 1790.420 17.010 1790.680 17.330 ;
        RECT 2161.640 14.970 2161.900 15.290 ;
        RECT 2161.700 2.000 2161.840 14.970 ;
        RECT 2161.490 -4.000 2162.050 2.000 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1597.650 1088.240 1597.970 1088.300 ;
        RECT 2173.570 1088.240 2173.890 1088.300 ;
        RECT 1597.650 1088.100 2173.890 1088.240 ;
        RECT 1597.650 1088.040 1597.970 1088.100 ;
        RECT 2173.570 1088.040 2173.890 1088.100 ;
      LAYER via ;
        RECT 1597.680 1088.040 1597.940 1088.300 ;
        RECT 2173.600 1088.040 2173.860 1088.300 ;
      LAYER met2 ;
        RECT 1597.590 1100.580 1597.870 1104.000 ;
        RECT 1597.590 1100.000 1597.880 1100.580 ;
        RECT 1597.740 1088.330 1597.880 1100.000 ;
        RECT 1597.680 1088.010 1597.940 1088.330 ;
        RECT 2173.600 1088.010 2173.860 1088.330 ;
        RECT 2173.660 16.730 2173.800 1088.010 ;
        RECT 2173.660 16.590 2179.320 16.730 ;
        RECT 2179.180 2.000 2179.320 16.590 ;
        RECT 2178.970 -4.000 2179.530 2.000 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1607.845 1087.405 1608.015 1089.615 ;
        RECT 1617.965 1087.405 1618.135 1089.615 ;
        RECT 1646.485 1089.445 1646.655 1090.295 ;
      LAYER mcon ;
        RECT 1646.485 1090.125 1646.655 1090.295 ;
        RECT 1607.845 1089.445 1608.015 1089.615 ;
        RECT 1617.965 1089.445 1618.135 1089.615 ;
      LAYER met1 ;
        RECT 1646.425 1090.280 1646.715 1090.325 ;
        RECT 1652.390 1090.280 1652.710 1090.340 ;
        RECT 1646.425 1090.140 1652.710 1090.280 ;
        RECT 1646.425 1090.095 1646.715 1090.140 ;
        RECT 1652.390 1090.080 1652.710 1090.140 ;
        RECT 1604.090 1089.600 1604.410 1089.660 ;
        RECT 1607.785 1089.600 1608.075 1089.645 ;
        RECT 1604.090 1089.460 1608.075 1089.600 ;
        RECT 1604.090 1089.400 1604.410 1089.460 ;
        RECT 1607.785 1089.415 1608.075 1089.460 ;
        RECT 1617.905 1089.600 1618.195 1089.645 ;
        RECT 1646.425 1089.600 1646.715 1089.645 ;
        RECT 1617.905 1089.460 1646.715 1089.600 ;
        RECT 1617.905 1089.415 1618.195 1089.460 ;
        RECT 1646.425 1089.415 1646.715 1089.460 ;
        RECT 1607.785 1087.560 1608.075 1087.605 ;
        RECT 1617.905 1087.560 1618.195 1087.605 ;
        RECT 1607.785 1087.420 1618.195 1087.560 ;
        RECT 1607.785 1087.375 1608.075 1087.420 ;
        RECT 1617.905 1087.375 1618.195 1087.420 ;
        RECT 1652.390 19.960 1652.710 20.020 ;
        RECT 2197.030 19.960 2197.350 20.020 ;
        RECT 1652.390 19.820 2197.350 19.960 ;
        RECT 1652.390 19.760 1652.710 19.820 ;
        RECT 2197.030 19.760 2197.350 19.820 ;
      LAYER via ;
        RECT 1652.420 1090.080 1652.680 1090.340 ;
        RECT 1604.120 1089.400 1604.380 1089.660 ;
        RECT 1652.420 19.760 1652.680 20.020 ;
        RECT 2197.060 19.760 2197.320 20.020 ;
      LAYER met2 ;
        RECT 1604.030 1100.580 1604.310 1104.000 ;
        RECT 1604.030 1100.000 1604.320 1100.580 ;
        RECT 1604.180 1089.690 1604.320 1100.000 ;
        RECT 1652.420 1090.050 1652.680 1090.370 ;
        RECT 1604.120 1089.370 1604.380 1089.690 ;
        RECT 1652.480 20.050 1652.620 1090.050 ;
        RECT 1652.420 19.730 1652.680 20.050 ;
        RECT 2197.060 19.730 2197.320 20.050 ;
        RECT 2197.120 2.000 2197.260 19.730 ;
        RECT 2196.910 -4.000 2197.470 2.000 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1655.685 1083.325 1655.855 1087.915 ;
      LAYER mcon ;
        RECT 1655.685 1087.745 1655.855 1087.915 ;
      LAYER met1 ;
        RECT 1655.625 1087.900 1655.915 1087.945 ;
        RECT 2214.970 1087.900 2215.290 1087.960 ;
        RECT 1655.625 1087.760 2215.290 1087.900 ;
        RECT 1655.625 1087.715 1655.915 1087.760 ;
        RECT 2214.970 1087.700 2215.290 1087.760 ;
        RECT 1610.070 1083.820 1610.390 1083.880 ;
        RECT 1610.070 1083.680 1652.620 1083.820 ;
        RECT 1610.070 1083.620 1610.390 1083.680 ;
        RECT 1652.480 1083.480 1652.620 1083.680 ;
        RECT 1655.625 1083.480 1655.915 1083.525 ;
        RECT 1652.480 1083.340 1655.915 1083.480 ;
        RECT 1655.625 1083.295 1655.915 1083.340 ;
      LAYER via ;
        RECT 2215.000 1087.700 2215.260 1087.960 ;
        RECT 1610.100 1083.620 1610.360 1083.880 ;
      LAYER met2 ;
        RECT 1610.010 1100.580 1610.290 1104.000 ;
        RECT 1610.010 1100.000 1610.300 1100.580 ;
        RECT 1610.160 1083.910 1610.300 1100.000 ;
        RECT 2215.000 1087.670 2215.260 1087.990 ;
        RECT 1610.100 1083.590 1610.360 1083.910 ;
        RECT 2215.060 2.000 2215.200 1087.670 ;
        RECT 2214.850 -4.000 2215.410 2.000 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1697.545 1087.065 1697.715 1088.595 ;
      LAYER mcon ;
        RECT 1697.545 1088.425 1697.715 1088.595 ;
      LAYER met1 ;
        RECT 1697.485 1088.580 1697.775 1088.625 ;
        RECT 1705.290 1088.580 1705.610 1088.640 ;
        RECT 1697.485 1088.440 1705.610 1088.580 ;
        RECT 1697.485 1088.395 1697.775 1088.440 ;
        RECT 1705.290 1088.380 1705.610 1088.440 ;
        RECT 1616.050 1087.220 1616.370 1087.280 ;
        RECT 1697.485 1087.220 1697.775 1087.265 ;
        RECT 1616.050 1087.080 1662.740 1087.220 ;
        RECT 1616.050 1087.020 1616.370 1087.080 ;
        RECT 1662.600 1086.880 1662.740 1087.080 ;
        RECT 1690.660 1087.080 1697.775 1087.220 ;
        RECT 1690.660 1086.880 1690.800 1087.080 ;
        RECT 1697.485 1087.035 1697.775 1087.080 ;
        RECT 1662.600 1086.740 1690.800 1086.880 ;
        RECT 1705.290 1083.820 1705.610 1083.880 ;
        RECT 1707.590 1083.820 1707.910 1083.880 ;
        RECT 1705.290 1083.680 1707.910 1083.820 ;
        RECT 1705.290 1083.620 1705.610 1083.680 ;
        RECT 1707.590 1083.620 1707.910 1083.680 ;
        RECT 1707.590 16.900 1707.910 16.960 ;
        RECT 2232.910 16.900 2233.230 16.960 ;
        RECT 1707.590 16.760 2233.230 16.900 ;
        RECT 1707.590 16.700 1707.910 16.760 ;
        RECT 2232.910 16.700 2233.230 16.760 ;
      LAYER via ;
        RECT 1705.320 1088.380 1705.580 1088.640 ;
        RECT 1616.080 1087.020 1616.340 1087.280 ;
        RECT 1705.320 1083.620 1705.580 1083.880 ;
        RECT 1707.620 1083.620 1707.880 1083.880 ;
        RECT 1707.620 16.700 1707.880 16.960 ;
        RECT 2232.940 16.700 2233.200 16.960 ;
      LAYER met2 ;
        RECT 1615.990 1100.580 1616.270 1104.000 ;
        RECT 1615.990 1100.000 1616.280 1100.580 ;
        RECT 1616.140 1087.310 1616.280 1100.000 ;
        RECT 1705.320 1088.350 1705.580 1088.670 ;
        RECT 1616.080 1086.990 1616.340 1087.310 ;
        RECT 1705.380 1083.910 1705.520 1088.350 ;
        RECT 1705.320 1083.590 1705.580 1083.910 ;
        RECT 1707.620 1083.590 1707.880 1083.910 ;
        RECT 1707.680 16.990 1707.820 1083.590 ;
        RECT 1707.620 16.670 1707.880 16.990 ;
        RECT 2232.940 16.670 2233.200 16.990 ;
        RECT 2233.000 2.000 2233.140 16.670 ;
        RECT 2232.790 -4.000 2233.350 2.000 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1118.790 1090.620 1119.110 1090.680 ;
        RECT 1119.710 1090.620 1120.030 1090.680 ;
        RECT 1118.790 1090.480 1120.030 1090.620 ;
        RECT 1118.790 1090.420 1119.110 1090.480 ;
        RECT 1119.710 1090.420 1120.030 1090.480 ;
        RECT 787.590 35.260 787.910 35.320 ;
        RECT 1118.790 35.260 1119.110 35.320 ;
        RECT 787.590 35.120 1119.110 35.260 ;
        RECT 787.590 35.060 787.910 35.120 ;
        RECT 1118.790 35.060 1119.110 35.120 ;
      LAYER via ;
        RECT 1118.820 1090.420 1119.080 1090.680 ;
        RECT 1119.740 1090.420 1120.000 1090.680 ;
        RECT 787.620 35.060 787.880 35.320 ;
        RECT 1118.820 35.060 1119.080 35.320 ;
      LAYER met2 ;
        RECT 1120.110 1100.650 1120.390 1104.000 ;
        RECT 1119.800 1100.510 1120.390 1100.650 ;
        RECT 1119.800 1090.710 1119.940 1100.510 ;
        RECT 1120.110 1100.000 1120.390 1100.510 ;
        RECT 1118.820 1090.390 1119.080 1090.710 ;
        RECT 1119.740 1090.390 1120.000 1090.710 ;
        RECT 1118.880 35.350 1119.020 1090.390 ;
        RECT 787.620 35.030 787.880 35.350 ;
        RECT 1118.820 35.030 1119.080 35.350 ;
        RECT 787.680 2.000 787.820 35.030 ;
        RECT 787.470 -4.000 788.030 2.000 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1622.490 1087.560 1622.810 1087.620 ;
        RECT 2249.470 1087.560 2249.790 1087.620 ;
        RECT 1622.490 1087.420 2249.790 1087.560 ;
        RECT 1622.490 1087.360 1622.810 1087.420 ;
        RECT 2249.470 1087.360 2249.790 1087.420 ;
      LAYER via ;
        RECT 1622.520 1087.360 1622.780 1087.620 ;
        RECT 2249.500 1087.360 2249.760 1087.620 ;
      LAYER met2 ;
        RECT 1622.430 1100.580 1622.710 1104.000 ;
        RECT 1622.430 1100.000 1622.720 1100.580 ;
        RECT 1622.580 1087.650 1622.720 1100.000 ;
        RECT 1622.520 1087.330 1622.780 1087.650 ;
        RECT 2249.500 1087.330 2249.760 1087.650 ;
        RECT 2249.560 17.410 2249.700 1087.330 ;
        RECT 2249.560 17.270 2251.080 17.410 ;
        RECT 2250.940 2.000 2251.080 17.270 ;
        RECT 2250.730 -4.000 2251.290 2.000 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1728.365 758.965 1728.535 807.075 ;
        RECT 1727.905 614.125 1728.075 662.235 ;
        RECT 1727.905 372.725 1728.075 420.835 ;
        RECT 1728.365 234.685 1728.535 300.135 ;
        RECT 1728.365 89.845 1728.535 137.955 ;
      LAYER mcon ;
        RECT 1728.365 806.905 1728.535 807.075 ;
        RECT 1727.905 662.065 1728.075 662.235 ;
        RECT 1727.905 420.665 1728.075 420.835 ;
        RECT 1728.365 299.965 1728.535 300.135 ;
        RECT 1728.365 137.785 1728.535 137.955 ;
      LAYER met1 ;
        RECT 1628.470 1083.480 1628.790 1083.540 ;
        RECT 1728.290 1083.480 1728.610 1083.540 ;
        RECT 1628.470 1083.340 1652.160 1083.480 ;
        RECT 1628.470 1083.280 1628.790 1083.340 ;
        RECT 1652.020 1082.800 1652.160 1083.340 ;
        RECT 1656.160 1083.340 1728.610 1083.480 ;
        RECT 1656.160 1082.800 1656.300 1083.340 ;
        RECT 1728.290 1083.280 1728.610 1083.340 ;
        RECT 1652.020 1082.660 1656.300 1082.800 ;
        RECT 1727.370 862.480 1727.690 862.540 ;
        RECT 1728.290 862.480 1728.610 862.540 ;
        RECT 1727.370 862.340 1728.610 862.480 ;
        RECT 1727.370 862.280 1727.690 862.340 ;
        RECT 1728.290 862.280 1728.610 862.340 ;
        RECT 1728.290 807.060 1728.610 807.120 ;
        RECT 1728.095 806.920 1728.610 807.060 ;
        RECT 1728.290 806.860 1728.610 806.920 ;
        RECT 1728.290 759.120 1728.610 759.180 ;
        RECT 1728.095 758.980 1728.610 759.120 ;
        RECT 1728.290 758.920 1728.610 758.980 ;
        RECT 1727.830 690.440 1728.150 690.500 ;
        RECT 1729.210 690.440 1729.530 690.500 ;
        RECT 1727.830 690.300 1729.530 690.440 ;
        RECT 1727.830 690.240 1728.150 690.300 ;
        RECT 1729.210 690.240 1729.530 690.300 ;
        RECT 1727.830 662.220 1728.150 662.280 ;
        RECT 1727.635 662.080 1728.150 662.220 ;
        RECT 1727.830 662.020 1728.150 662.080 ;
        RECT 1727.830 614.280 1728.150 614.340 ;
        RECT 1727.635 614.140 1728.150 614.280 ;
        RECT 1727.830 614.080 1728.150 614.140 ;
        RECT 1727.830 420.820 1728.150 420.880 ;
        RECT 1727.635 420.680 1728.150 420.820 ;
        RECT 1727.830 420.620 1728.150 420.680 ;
        RECT 1727.845 372.880 1728.135 372.925 ;
        RECT 1728.290 372.880 1728.610 372.940 ;
        RECT 1727.845 372.740 1728.610 372.880 ;
        RECT 1727.845 372.695 1728.135 372.740 ;
        RECT 1728.290 372.680 1728.610 372.740 ;
        RECT 1727.830 300.120 1728.150 300.180 ;
        RECT 1728.305 300.120 1728.595 300.165 ;
        RECT 1727.830 299.980 1728.595 300.120 ;
        RECT 1727.830 299.920 1728.150 299.980 ;
        RECT 1728.305 299.935 1728.595 299.980 ;
        RECT 1728.290 234.840 1728.610 234.900 ;
        RECT 1728.290 234.700 1728.805 234.840 ;
        RECT 1728.290 234.640 1728.610 234.700 ;
        RECT 1728.290 137.940 1728.610 138.000 ;
        RECT 1728.095 137.800 1728.610 137.940 ;
        RECT 1728.290 137.740 1728.610 137.800 ;
        RECT 1728.290 90.000 1728.610 90.060 ;
        RECT 1728.095 89.860 1728.610 90.000 ;
        RECT 1728.290 89.800 1728.610 89.860 ;
        RECT 1728.290 20.300 1728.610 20.360 ;
        RECT 2268.330 20.300 2268.650 20.360 ;
        RECT 1728.290 20.160 2268.650 20.300 ;
        RECT 1728.290 20.100 1728.610 20.160 ;
        RECT 2268.330 20.100 2268.650 20.160 ;
      LAYER via ;
        RECT 1628.500 1083.280 1628.760 1083.540 ;
        RECT 1728.320 1083.280 1728.580 1083.540 ;
        RECT 1727.400 862.280 1727.660 862.540 ;
        RECT 1728.320 862.280 1728.580 862.540 ;
        RECT 1728.320 806.860 1728.580 807.120 ;
        RECT 1728.320 758.920 1728.580 759.180 ;
        RECT 1727.860 690.240 1728.120 690.500 ;
        RECT 1729.240 690.240 1729.500 690.500 ;
        RECT 1727.860 662.020 1728.120 662.280 ;
        RECT 1727.860 614.080 1728.120 614.340 ;
        RECT 1727.860 420.620 1728.120 420.880 ;
        RECT 1728.320 372.680 1728.580 372.940 ;
        RECT 1727.860 299.920 1728.120 300.180 ;
        RECT 1728.320 234.640 1728.580 234.900 ;
        RECT 1728.320 137.740 1728.580 138.000 ;
        RECT 1728.320 89.800 1728.580 90.060 ;
        RECT 1728.320 20.100 1728.580 20.360 ;
        RECT 2268.360 20.100 2268.620 20.360 ;
      LAYER met2 ;
        RECT 1628.410 1100.580 1628.690 1104.000 ;
        RECT 1628.410 1100.000 1628.700 1100.580 ;
        RECT 1628.560 1083.570 1628.700 1100.000 ;
        RECT 1628.500 1083.250 1628.760 1083.570 ;
        RECT 1728.320 1083.250 1728.580 1083.570 ;
        RECT 1728.380 980.290 1728.520 1083.250 ;
        RECT 1727.920 980.150 1728.520 980.290 ;
        RECT 1727.920 979.610 1728.060 980.150 ;
        RECT 1727.920 979.470 1728.520 979.610 ;
        RECT 1728.380 862.570 1728.520 979.470 ;
        RECT 1727.400 862.250 1727.660 862.570 ;
        RECT 1728.320 862.250 1728.580 862.570 ;
        RECT 1727.460 814.485 1727.600 862.250 ;
        RECT 1727.390 814.115 1727.670 814.485 ;
        RECT 1728.310 814.115 1728.590 814.485 ;
        RECT 1728.380 807.150 1728.520 814.115 ;
        RECT 1728.320 806.830 1728.580 807.150 ;
        RECT 1728.320 758.890 1728.580 759.210 ;
        RECT 1728.380 741.610 1728.520 758.890 ;
        RECT 1727.920 741.470 1728.520 741.610 ;
        RECT 1727.920 690.530 1728.060 741.470 ;
        RECT 1727.860 690.210 1728.120 690.530 ;
        RECT 1729.240 690.210 1729.500 690.530 ;
        RECT 1729.300 662.845 1729.440 690.210 ;
        RECT 1728.310 662.730 1728.590 662.845 ;
        RECT 1727.920 662.590 1728.590 662.730 ;
        RECT 1727.920 662.310 1728.060 662.590 ;
        RECT 1728.310 662.475 1728.590 662.590 ;
        RECT 1729.230 662.475 1729.510 662.845 ;
        RECT 1727.860 661.990 1728.120 662.310 ;
        RECT 1727.860 614.050 1728.120 614.370 ;
        RECT 1727.920 613.770 1728.060 614.050 ;
        RECT 1727.460 613.630 1728.060 613.770 ;
        RECT 1727.460 572.290 1727.600 613.630 ;
        RECT 1727.460 572.150 1728.060 572.290 ;
        RECT 1727.920 524.010 1728.060 572.150 ;
        RECT 1727.920 523.870 1728.520 524.010 ;
        RECT 1728.380 434.930 1728.520 523.870 ;
        RECT 1727.920 434.790 1728.520 434.930 ;
        RECT 1727.920 420.910 1728.060 434.790 ;
        RECT 1727.860 420.590 1728.120 420.910 ;
        RECT 1728.320 372.650 1728.580 372.970 ;
        RECT 1728.380 324.090 1728.520 372.650 ;
        RECT 1727.920 323.950 1728.520 324.090 ;
        RECT 1727.920 300.210 1728.060 323.950 ;
        RECT 1727.860 299.890 1728.120 300.210 ;
        RECT 1728.320 234.610 1728.580 234.930 ;
        RECT 1728.380 138.030 1728.520 234.610 ;
        RECT 1728.320 137.710 1728.580 138.030 ;
        RECT 1728.320 89.770 1728.580 90.090 ;
        RECT 1728.380 20.390 1728.520 89.770 ;
        RECT 1728.320 20.070 1728.580 20.390 ;
        RECT 2268.360 20.070 2268.620 20.390 ;
        RECT 2268.420 2.000 2268.560 20.070 ;
        RECT 2268.210 -4.000 2268.770 2.000 ;
      LAYER via2 ;
        RECT 1727.390 814.160 1727.670 814.440 ;
        RECT 1728.310 814.160 1728.590 814.440 ;
        RECT 1728.310 662.520 1728.590 662.800 ;
        RECT 1729.230 662.520 1729.510 662.800 ;
      LAYER met3 ;
        RECT 1727.365 814.450 1727.695 814.465 ;
        RECT 1728.285 814.450 1728.615 814.465 ;
        RECT 1727.365 814.150 1728.615 814.450 ;
        RECT 1727.365 814.135 1727.695 814.150 ;
        RECT 1728.285 814.135 1728.615 814.150 ;
        RECT 1728.285 662.810 1728.615 662.825 ;
        RECT 1729.205 662.810 1729.535 662.825 ;
        RECT 1728.285 662.510 1729.535 662.810 ;
        RECT 1728.285 662.495 1728.615 662.510 ;
        RECT 1729.205 662.495 1729.535 662.510 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1702.605 1087.065 1703.695 1087.235 ;
        RECT 1702.605 1086.385 1702.775 1087.065 ;
      LAYER mcon ;
        RECT 1703.525 1087.065 1703.695 1087.235 ;
      LAYER met1 ;
        RECT 1703.465 1087.220 1703.755 1087.265 ;
        RECT 2283.970 1087.220 2284.290 1087.280 ;
        RECT 1703.465 1087.080 2284.290 1087.220 ;
        RECT 1703.465 1087.035 1703.755 1087.080 ;
        RECT 2283.970 1087.020 2284.290 1087.080 ;
        RECT 1634.450 1086.540 1634.770 1086.600 ;
        RECT 1702.545 1086.540 1702.835 1086.585 ;
        RECT 1634.450 1086.400 1702.835 1086.540 ;
        RECT 1634.450 1086.340 1634.770 1086.400 ;
        RECT 1702.545 1086.355 1702.835 1086.400 ;
      LAYER via ;
        RECT 2284.000 1087.020 2284.260 1087.280 ;
        RECT 1634.480 1086.340 1634.740 1086.600 ;
      LAYER met2 ;
        RECT 1634.390 1100.580 1634.670 1104.000 ;
        RECT 1634.390 1100.000 1634.680 1100.580 ;
        RECT 1634.540 1086.630 1634.680 1100.000 ;
        RECT 2284.000 1086.990 2284.260 1087.310 ;
        RECT 1634.480 1086.310 1634.740 1086.630 ;
        RECT 2284.060 16.730 2284.200 1086.990 ;
        RECT 2284.060 16.590 2286.500 16.730 ;
        RECT 2286.360 2.000 2286.500 16.590 ;
        RECT 2286.150 -4.000 2286.710 2.000 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1662.125 1086.725 1662.295 1089.275 ;
        RECT 1676.845 1087.065 1677.015 1089.275 ;
        RECT 1687.425 1089.105 1689.435 1089.275 ;
        RECT 1703.065 1089.105 1703.235 1090.295 ;
        RECT 1683.285 1087.065 1683.455 1088.595 ;
        RECT 1687.425 1088.425 1687.595 1089.105 ;
      LAYER mcon ;
        RECT 1703.065 1090.125 1703.235 1090.295 ;
        RECT 1662.125 1089.105 1662.295 1089.275 ;
        RECT 1676.845 1089.105 1677.015 1089.275 ;
        RECT 1689.265 1089.105 1689.435 1089.275 ;
        RECT 1683.285 1088.425 1683.455 1088.595 ;
      LAYER met1 ;
        RECT 1703.005 1090.280 1703.295 1090.325 ;
        RECT 1703.005 1090.140 1704.140 1090.280 ;
        RECT 1703.005 1090.095 1703.295 1090.140 ;
        RECT 1704.000 1089.940 1704.140 1090.140 ;
        RECT 1704.000 1089.800 1746.000 1089.940 ;
        RECT 1662.065 1089.260 1662.355 1089.305 ;
        RECT 1676.785 1089.260 1677.075 1089.305 ;
        RECT 1662.065 1089.120 1677.075 1089.260 ;
        RECT 1662.065 1089.075 1662.355 1089.120 ;
        RECT 1676.785 1089.075 1677.075 1089.120 ;
        RECT 1689.205 1089.260 1689.495 1089.305 ;
        RECT 1703.005 1089.260 1703.295 1089.305 ;
        RECT 1689.205 1089.120 1703.295 1089.260 ;
        RECT 1745.860 1089.260 1746.000 1089.800 ;
        RECT 1762.790 1089.260 1763.110 1089.320 ;
        RECT 1745.860 1089.120 1763.110 1089.260 ;
        RECT 1689.205 1089.075 1689.495 1089.120 ;
        RECT 1703.005 1089.075 1703.295 1089.120 ;
        RECT 1762.790 1089.060 1763.110 1089.120 ;
        RECT 1683.225 1088.580 1683.515 1088.625 ;
        RECT 1687.365 1088.580 1687.655 1088.625 ;
        RECT 1683.225 1088.440 1687.655 1088.580 ;
        RECT 1683.225 1088.395 1683.515 1088.440 ;
        RECT 1687.365 1088.395 1687.655 1088.440 ;
        RECT 1676.785 1087.220 1677.075 1087.265 ;
        RECT 1683.225 1087.220 1683.515 1087.265 ;
        RECT 1676.785 1087.080 1683.515 1087.220 ;
        RECT 1676.785 1087.035 1677.075 1087.080 ;
        RECT 1683.225 1087.035 1683.515 1087.080 ;
        RECT 1640.890 1086.880 1641.210 1086.940 ;
        RECT 1662.065 1086.880 1662.355 1086.925 ;
        RECT 1640.890 1086.740 1662.355 1086.880 ;
        RECT 1640.890 1086.680 1641.210 1086.740 ;
        RECT 1662.065 1086.695 1662.355 1086.740 ;
        RECT 1762.330 20.640 1762.650 20.700 ;
        RECT 2304.210 20.640 2304.530 20.700 ;
        RECT 1762.330 20.500 2304.530 20.640 ;
        RECT 1762.330 20.440 1762.650 20.500 ;
        RECT 2304.210 20.440 2304.530 20.500 ;
      LAYER via ;
        RECT 1762.820 1089.060 1763.080 1089.320 ;
        RECT 1640.920 1086.680 1641.180 1086.940 ;
        RECT 1762.360 20.440 1762.620 20.700 ;
        RECT 2304.240 20.440 2304.500 20.700 ;
      LAYER met2 ;
        RECT 1640.830 1100.580 1641.110 1104.000 ;
        RECT 1640.830 1100.000 1641.120 1100.580 ;
        RECT 1640.980 1086.970 1641.120 1100.000 ;
        RECT 1762.820 1089.030 1763.080 1089.350 ;
        RECT 1640.920 1086.650 1641.180 1086.970 ;
        RECT 1762.880 41.210 1763.020 1089.030 ;
        RECT 1762.420 41.070 1763.020 41.210 ;
        RECT 1762.420 20.730 1762.560 41.070 ;
        RECT 1762.360 20.410 1762.620 20.730 ;
        RECT 2304.240 20.410 2304.500 20.730 ;
        RECT 2304.300 2.000 2304.440 20.410 ;
        RECT 2304.090 -4.000 2304.650 2.000 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1703.525 1089.785 1704.155 1089.955 ;
        RECT 1703.985 1086.725 1704.155 1089.785 ;
      LAYER met1 ;
        RECT 1703.465 1089.940 1703.755 1089.985 ;
        RECT 1656.620 1089.800 1703.755 1089.940 ;
        RECT 1646.870 1089.600 1647.190 1089.660 ;
        RECT 1656.620 1089.600 1656.760 1089.800 ;
        RECT 1703.465 1089.755 1703.755 1089.800 ;
        RECT 1646.870 1089.460 1656.760 1089.600 ;
        RECT 1646.870 1089.400 1647.190 1089.460 ;
        RECT 1703.925 1086.880 1704.215 1086.925 ;
        RECT 2318.470 1086.880 2318.790 1086.940 ;
        RECT 1703.925 1086.740 2318.790 1086.880 ;
        RECT 1703.925 1086.695 1704.215 1086.740 ;
        RECT 2318.470 1086.680 2318.790 1086.740 ;
        RECT 2318.470 2.620 2318.790 2.680 ;
        RECT 2322.150 2.620 2322.470 2.680 ;
        RECT 2318.470 2.480 2322.470 2.620 ;
        RECT 2318.470 2.420 2318.790 2.480 ;
        RECT 2322.150 2.420 2322.470 2.480 ;
      LAYER via ;
        RECT 1646.900 1089.400 1647.160 1089.660 ;
        RECT 2318.500 1086.680 2318.760 1086.940 ;
        RECT 2318.500 2.420 2318.760 2.680 ;
        RECT 2322.180 2.420 2322.440 2.680 ;
      LAYER met2 ;
        RECT 1646.810 1100.580 1647.090 1104.000 ;
        RECT 1646.810 1100.000 1647.100 1100.580 ;
        RECT 1646.960 1089.690 1647.100 1100.000 ;
        RECT 1646.900 1089.370 1647.160 1089.690 ;
        RECT 2318.500 1086.650 2318.760 1086.970 ;
        RECT 2318.560 2.710 2318.700 1086.650 ;
        RECT 2318.500 2.390 2318.760 2.710 ;
        RECT 2322.180 2.390 2322.440 2.710 ;
        RECT 2322.240 2.000 2322.380 2.390 ;
        RECT 2322.030 -4.000 2322.590 2.000 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1652.850 1083.820 1653.170 1083.880 ;
        RECT 1686.890 1083.820 1687.210 1083.880 ;
        RECT 1652.850 1083.680 1687.210 1083.820 ;
        RECT 1652.850 1083.620 1653.170 1083.680 ;
        RECT 1686.890 1083.620 1687.210 1083.680 ;
        RECT 1686.890 19.620 1687.210 19.680 ;
        RECT 2339.630 19.620 2339.950 19.680 ;
        RECT 1686.890 19.480 2339.950 19.620 ;
        RECT 1686.890 19.420 1687.210 19.480 ;
        RECT 2339.630 19.420 2339.950 19.480 ;
      LAYER via ;
        RECT 1652.880 1083.620 1653.140 1083.880 ;
        RECT 1686.920 1083.620 1687.180 1083.880 ;
        RECT 1686.920 19.420 1687.180 19.680 ;
        RECT 2339.660 19.420 2339.920 19.680 ;
      LAYER met2 ;
        RECT 1652.790 1100.580 1653.070 1104.000 ;
        RECT 1652.790 1100.000 1653.080 1100.580 ;
        RECT 1652.940 1083.910 1653.080 1100.000 ;
        RECT 1652.880 1083.590 1653.140 1083.910 ;
        RECT 1686.920 1083.590 1687.180 1083.910 ;
        RECT 1686.980 19.710 1687.120 1083.590 ;
        RECT 1686.920 19.390 1687.180 19.710 ;
        RECT 2339.660 19.390 2339.920 19.710 ;
        RECT 2339.720 2.000 2339.860 19.390 ;
        RECT 2339.510 -4.000 2340.070 2.000 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1658.770 1100.580 1659.050 1104.000 ;
        RECT 1658.770 1100.000 1659.060 1100.580 ;
        RECT 1658.920 1086.485 1659.060 1100.000 ;
        RECT 1658.850 1086.115 1659.130 1086.485 ;
        RECT 2352.990 1086.115 2353.270 1086.485 ;
        RECT 2353.060 2.450 2353.200 1086.115 ;
        RECT 2353.060 2.310 2357.800 2.450 ;
        RECT 2357.660 2.000 2357.800 2.310 ;
        RECT 2357.450 -4.000 2358.010 2.000 ;
      LAYER via2 ;
        RECT 1658.850 1086.160 1659.130 1086.440 ;
        RECT 2352.990 1086.160 2353.270 1086.440 ;
      LAYER met3 ;
        RECT 1658.825 1086.450 1659.155 1086.465 ;
        RECT 2352.965 1086.450 2353.295 1086.465 ;
        RECT 1658.825 1086.150 2353.295 1086.450 ;
        RECT 1658.825 1086.135 1659.155 1086.150 ;
        RECT 2352.965 1086.135 2353.295 1086.150 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1666.650 1072.940 1666.970 1073.000 ;
        RECT 1669.410 1072.940 1669.730 1073.000 ;
        RECT 1666.650 1072.800 1669.730 1072.940 ;
        RECT 1666.650 1072.740 1666.970 1072.800 ;
        RECT 1669.410 1072.740 1669.730 1072.800 ;
        RECT 1669.410 19.280 1669.730 19.340 ;
        RECT 2375.510 19.280 2375.830 19.340 ;
        RECT 1669.410 19.140 2375.830 19.280 ;
        RECT 1669.410 19.080 1669.730 19.140 ;
        RECT 2375.510 19.080 2375.830 19.140 ;
      LAYER via ;
        RECT 1666.680 1072.740 1666.940 1073.000 ;
        RECT 1669.440 1072.740 1669.700 1073.000 ;
        RECT 1669.440 19.080 1669.700 19.340 ;
        RECT 2375.540 19.080 2375.800 19.340 ;
      LAYER met2 ;
        RECT 1665.210 1100.650 1665.490 1104.000 ;
        RECT 1665.210 1100.510 1666.880 1100.650 ;
        RECT 1665.210 1100.000 1665.490 1100.510 ;
        RECT 1666.740 1073.030 1666.880 1100.510 ;
        RECT 1666.680 1072.710 1666.940 1073.030 ;
        RECT 1669.440 1072.710 1669.700 1073.030 ;
        RECT 1669.500 19.370 1669.640 1072.710 ;
        RECT 1669.440 19.050 1669.700 19.370 ;
        RECT 2375.540 19.050 2375.800 19.370 ;
        RECT 2375.600 2.000 2375.740 19.050 ;
        RECT 2375.390 -4.000 2375.950 2.000 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1697.085 1086.725 1697.255 1090.975 ;
      LAYER mcon ;
        RECT 1697.085 1090.805 1697.255 1090.975 ;
      LAYER met1 ;
        RECT 1673.090 1090.960 1673.410 1091.020 ;
        RECT 1697.025 1090.960 1697.315 1091.005 ;
        RECT 1673.090 1090.820 1697.315 1090.960 ;
        RECT 1673.090 1090.760 1673.410 1090.820 ;
        RECT 1697.025 1090.775 1697.315 1090.820 ;
        RECT 1697.025 1086.880 1697.315 1086.925 ;
        RECT 1697.025 1086.740 1703.220 1086.880 ;
        RECT 1697.025 1086.695 1697.315 1086.740 ;
        RECT 1703.080 1086.540 1703.220 1086.740 ;
        RECT 2387.470 1086.540 2387.790 1086.600 ;
        RECT 1703.080 1086.400 2387.790 1086.540 ;
        RECT 2387.470 1086.340 2387.790 1086.400 ;
        RECT 2387.470 19.280 2387.790 19.340 ;
        RECT 2393.450 19.280 2393.770 19.340 ;
        RECT 2387.470 19.140 2393.770 19.280 ;
        RECT 2387.470 19.080 2387.790 19.140 ;
        RECT 2393.450 19.080 2393.770 19.140 ;
      LAYER via ;
        RECT 1673.120 1090.760 1673.380 1091.020 ;
        RECT 2387.500 1086.340 2387.760 1086.600 ;
        RECT 2387.500 19.080 2387.760 19.340 ;
        RECT 2393.480 19.080 2393.740 19.340 ;
      LAYER met2 ;
        RECT 1671.190 1100.650 1671.470 1104.000 ;
        RECT 1671.190 1100.510 1673.320 1100.650 ;
        RECT 1671.190 1100.000 1671.470 1100.510 ;
        RECT 1673.180 1091.050 1673.320 1100.510 ;
        RECT 1673.120 1090.730 1673.380 1091.050 ;
        RECT 2387.500 1086.310 2387.760 1086.630 ;
        RECT 2387.560 19.370 2387.700 1086.310 ;
        RECT 2387.500 19.050 2387.760 19.370 ;
        RECT 2393.480 19.050 2393.740 19.370 ;
        RECT 2393.540 2.000 2393.680 19.050 ;
        RECT 2393.330 -4.000 2393.890 2.000 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1677.230 1089.260 1677.550 1089.320 ;
        RECT 1683.210 1089.260 1683.530 1089.320 ;
        RECT 1677.230 1089.120 1683.530 1089.260 ;
        RECT 1677.230 1089.060 1677.550 1089.120 ;
        RECT 1683.210 1089.060 1683.530 1089.120 ;
        RECT 1683.210 18.940 1683.530 19.000 ;
        RECT 2411.390 18.940 2411.710 19.000 ;
        RECT 1683.210 18.800 2411.710 18.940 ;
        RECT 1683.210 18.740 1683.530 18.800 ;
        RECT 2411.390 18.740 2411.710 18.800 ;
      LAYER via ;
        RECT 1677.260 1089.060 1677.520 1089.320 ;
        RECT 1683.240 1089.060 1683.500 1089.320 ;
        RECT 1683.240 18.740 1683.500 19.000 ;
        RECT 2411.420 18.740 2411.680 19.000 ;
      LAYER met2 ;
        RECT 1677.170 1100.580 1677.450 1104.000 ;
        RECT 1677.170 1100.000 1677.460 1100.580 ;
        RECT 1677.320 1089.350 1677.460 1100.000 ;
        RECT 1677.260 1089.030 1677.520 1089.350 ;
        RECT 1683.240 1089.030 1683.500 1089.350 ;
        RECT 1683.300 19.030 1683.440 1089.030 ;
        RECT 1683.240 18.710 1683.500 19.030 ;
        RECT 2411.420 18.710 2411.680 19.030 ;
        RECT 2411.480 2.000 2411.620 18.710 ;
        RECT 2411.270 -4.000 2411.830 2.000 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 805.530 34.920 805.850 34.980 ;
        RECT 1125.230 34.920 1125.550 34.980 ;
        RECT 805.530 34.780 1125.550 34.920 ;
        RECT 805.530 34.720 805.850 34.780 ;
        RECT 1125.230 34.720 1125.550 34.780 ;
      LAYER via ;
        RECT 805.560 34.720 805.820 34.980 ;
        RECT 1125.260 34.720 1125.520 34.980 ;
      LAYER met2 ;
        RECT 1126.090 1100.650 1126.370 1104.000 ;
        RECT 1125.320 1100.510 1126.370 1100.650 ;
        RECT 1125.320 35.010 1125.460 1100.510 ;
        RECT 1126.090 1100.000 1126.370 1100.510 ;
        RECT 805.560 34.690 805.820 35.010 ;
        RECT 1125.260 34.690 1125.520 35.010 ;
        RECT 805.620 2.000 805.760 34.690 ;
        RECT 805.410 -4.000 805.970 2.000 ;
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.000 2917.370 2.000 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 851.010 1100.650 851.290 1104.000 ;
        RECT 850.240 1100.510 851.290 1100.650 ;
        RECT 850.240 24.325 850.380 1100.510 ;
        RECT 851.010 1100.000 851.290 1100.510 ;
        RECT 2.850 23.955 3.130 24.325 ;
        RECT 850.170 23.955 850.450 24.325 ;
        RECT 2.920 2.000 3.060 23.955 ;
        RECT 2.710 -4.000 3.270 2.000 ;
      LAYER via2 ;
        RECT 2.850 24.000 3.130 24.280 ;
        RECT 850.170 24.000 850.450 24.280 ;
      LAYER met3 ;
        RECT 2.825 24.290 3.155 24.305 ;
        RECT 850.145 24.290 850.475 24.305 ;
        RECT 2.825 23.990 850.475 24.290 ;
        RECT 2.825 23.975 3.155 23.990 ;
        RECT 850.145 23.975 850.475 23.990 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 849.230 1052.200 849.550 1052.260 ;
        RECT 851.530 1052.200 851.850 1052.260 ;
        RECT 849.230 1052.060 851.850 1052.200 ;
        RECT 849.230 1052.000 849.550 1052.060 ;
        RECT 851.530 1052.000 851.850 1052.060 ;
        RECT 8.350 24.040 8.670 24.100 ;
        RECT 849.230 24.040 849.550 24.100 ;
        RECT 8.350 23.900 849.550 24.040 ;
        RECT 8.350 23.840 8.670 23.900 ;
        RECT 849.230 23.840 849.550 23.900 ;
      LAYER via ;
        RECT 849.260 1052.000 849.520 1052.260 ;
        RECT 851.560 1052.000 851.820 1052.260 ;
        RECT 8.380 23.840 8.640 24.100 ;
        RECT 849.260 23.840 849.520 24.100 ;
      LAYER met2 ;
        RECT 852.850 1100.650 853.130 1104.000 ;
        RECT 851.620 1100.510 853.130 1100.650 ;
        RECT 851.620 1052.290 851.760 1100.510 ;
        RECT 852.850 1100.000 853.130 1100.510 ;
        RECT 849.260 1051.970 849.520 1052.290 ;
        RECT 851.560 1051.970 851.820 1052.290 ;
        RECT 849.320 24.130 849.460 1051.970 ;
        RECT 8.380 23.810 8.640 24.130 ;
        RECT 849.260 23.810 849.520 24.130 ;
        RECT 8.440 2.000 8.580 23.810 ;
        RECT 8.230 -4.000 8.790 2.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 849.690 1052.540 850.010 1052.600 ;
        RECT 853.370 1052.540 853.690 1052.600 ;
        RECT 849.690 1052.400 853.690 1052.540 ;
        RECT 849.690 1052.340 850.010 1052.400 ;
        RECT 853.370 1052.340 853.690 1052.400 ;
        RECT 14.330 24.380 14.650 24.440 ;
        RECT 849.690 24.380 850.010 24.440 ;
        RECT 14.330 24.240 850.010 24.380 ;
        RECT 14.330 24.180 14.650 24.240 ;
        RECT 849.690 24.180 850.010 24.240 ;
      LAYER via ;
        RECT 849.720 1052.340 849.980 1052.600 ;
        RECT 853.400 1052.340 853.660 1052.600 ;
        RECT 14.360 24.180 14.620 24.440 ;
        RECT 849.720 24.180 849.980 24.440 ;
      LAYER met2 ;
        RECT 854.690 1100.650 854.970 1104.000 ;
        RECT 853.460 1100.510 854.970 1100.650 ;
        RECT 853.460 1052.630 853.600 1100.510 ;
        RECT 854.690 1100.000 854.970 1100.510 ;
        RECT 849.720 1052.310 849.980 1052.630 ;
        RECT 853.400 1052.310 853.660 1052.630 ;
        RECT 849.780 24.470 849.920 1052.310 ;
        RECT 14.360 24.150 14.620 24.470 ;
        RECT 849.720 24.150 849.980 24.470 ;
        RECT 14.420 2.000 14.560 24.150 ;
        RECT 14.210 -4.000 14.770 2.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 38.250 24.720 38.570 24.780 ;
        RECT 863.490 24.720 863.810 24.780 ;
        RECT 38.250 24.580 863.810 24.720 ;
        RECT 38.250 24.520 38.570 24.580 ;
        RECT 863.490 24.520 863.810 24.580 ;
      LAYER via ;
        RECT 38.280 24.520 38.540 24.780 ;
        RECT 863.520 24.520 863.780 24.780 ;
      LAYER met2 ;
        RECT 862.970 1100.650 863.250 1104.000 ;
        RECT 862.970 1100.510 863.720 1100.650 ;
        RECT 862.970 1100.000 863.250 1100.510 ;
        RECT 863.580 24.810 863.720 1100.510 ;
        RECT 38.280 24.490 38.540 24.810 ;
        RECT 863.520 24.490 863.780 24.810 ;
        RECT 38.340 2.000 38.480 24.490 ;
        RECT 38.130 -4.000 38.690 2.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 240.650 25.740 240.970 25.800 ;
        RECT 932.490 25.740 932.810 25.800 ;
        RECT 240.650 25.600 932.810 25.740 ;
        RECT 240.650 25.540 240.970 25.600 ;
        RECT 932.490 25.540 932.810 25.600 ;
      LAYER via ;
        RECT 240.680 25.540 240.940 25.800 ;
        RECT 932.520 25.540 932.780 25.800 ;
      LAYER met2 ;
        RECT 932.430 1100.580 932.710 1104.000 ;
        RECT 932.430 1100.000 932.720 1100.580 ;
        RECT 932.580 25.830 932.720 1100.000 ;
        RECT 240.680 25.510 240.940 25.830 ;
        RECT 932.520 25.510 932.780 25.830 ;
        RECT 240.740 2.000 240.880 25.510 ;
        RECT 240.530 -4.000 241.090 2.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 258.130 26.080 258.450 26.140 ;
        RECT 938.930 26.080 939.250 26.140 ;
        RECT 258.130 25.940 939.250 26.080 ;
        RECT 258.130 25.880 258.450 25.940 ;
        RECT 938.930 25.880 939.250 25.940 ;
      LAYER via ;
        RECT 258.160 25.880 258.420 26.140 ;
        RECT 938.960 25.880 939.220 26.140 ;
      LAYER met2 ;
        RECT 938.410 1100.650 938.690 1104.000 ;
        RECT 938.410 1100.510 939.160 1100.650 ;
        RECT 938.410 1100.000 938.690 1100.510 ;
        RECT 939.020 26.170 939.160 1100.510 ;
        RECT 258.160 25.850 258.420 26.170 ;
        RECT 938.960 25.850 939.220 26.170 ;
        RECT 258.220 2.000 258.360 25.850 ;
        RECT 258.010 -4.000 258.570 2.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 939.850 1052.200 940.170 1052.260 ;
        RECT 943.070 1052.200 943.390 1052.260 ;
        RECT 939.850 1052.060 943.390 1052.200 ;
        RECT 939.850 1052.000 940.170 1052.060 ;
        RECT 943.070 1052.000 943.390 1052.060 ;
        RECT 276.070 26.420 276.390 26.480 ;
        RECT 939.850 26.420 940.170 26.480 ;
        RECT 276.070 26.280 940.170 26.420 ;
        RECT 276.070 26.220 276.390 26.280 ;
        RECT 939.850 26.220 940.170 26.280 ;
      LAYER via ;
        RECT 939.880 1052.000 940.140 1052.260 ;
        RECT 943.100 1052.000 943.360 1052.260 ;
        RECT 276.100 26.220 276.360 26.480 ;
        RECT 939.880 26.220 940.140 26.480 ;
      LAYER met2 ;
        RECT 944.850 1100.650 945.130 1104.000 ;
        RECT 943.160 1100.510 945.130 1100.650 ;
        RECT 943.160 1052.290 943.300 1100.510 ;
        RECT 944.850 1100.000 945.130 1100.510 ;
        RECT 939.880 1051.970 940.140 1052.290 ;
        RECT 943.100 1051.970 943.360 1052.290 ;
        RECT 939.940 26.510 940.080 1051.970 ;
        RECT 276.100 26.190 276.360 26.510 ;
        RECT 939.880 26.190 940.140 26.510 ;
        RECT 276.160 2.000 276.300 26.190 ;
        RECT 275.950 -4.000 276.510 2.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 947.745 138.125 947.915 203.575 ;
      LAYER mcon ;
        RECT 947.745 203.405 947.915 203.575 ;
      LAYER met1 ;
        RECT 946.750 1062.740 947.070 1062.800 ;
        RECT 950.890 1062.740 951.210 1062.800 ;
        RECT 946.750 1062.600 951.210 1062.740 ;
        RECT 946.750 1062.540 947.070 1062.600 ;
        RECT 950.890 1062.540 951.210 1062.600 ;
        RECT 947.210 931.640 947.530 931.900 ;
        RECT 947.300 931.160 947.440 931.640 ;
        RECT 947.670 931.160 947.990 931.220 ;
        RECT 947.300 931.020 947.990 931.160 ;
        RECT 947.670 930.960 947.990 931.020 ;
        RECT 947.210 862.820 947.530 862.880 ;
        RECT 947.670 862.820 947.990 862.880 ;
        RECT 947.210 862.680 947.990 862.820 ;
        RECT 947.210 862.620 947.530 862.680 ;
        RECT 947.670 862.620 947.990 862.680 ;
        RECT 946.750 821.000 947.070 821.060 ;
        RECT 947.210 821.000 947.530 821.060 ;
        RECT 946.750 820.860 947.530 821.000 ;
        RECT 946.750 820.800 947.070 820.860 ;
        RECT 947.210 820.800 947.530 820.860 ;
        RECT 946.750 738.520 947.070 738.780 ;
        RECT 946.840 738.100 946.980 738.520 ;
        RECT 946.750 737.840 947.070 738.100 ;
        RECT 946.750 641.620 947.070 641.880 ;
        RECT 946.840 641.480 946.980 641.620 ;
        RECT 947.210 641.480 947.530 641.540 ;
        RECT 946.840 641.340 947.530 641.480 ;
        RECT 947.210 641.280 947.530 641.340 ;
        RECT 946.750 579.600 947.070 579.660 ;
        RECT 947.210 579.600 947.530 579.660 ;
        RECT 946.750 579.460 947.530 579.600 ;
        RECT 946.750 579.400 947.070 579.460 ;
        RECT 947.210 579.400 947.530 579.460 ;
        RECT 946.750 379.680 947.070 379.740 ;
        RECT 947.210 379.680 947.530 379.740 ;
        RECT 946.750 379.540 947.530 379.680 ;
        RECT 946.750 379.480 947.070 379.540 ;
        RECT 947.210 379.480 947.530 379.540 ;
        RECT 947.210 241.300 947.530 241.360 ;
        RECT 947.670 241.300 947.990 241.360 ;
        RECT 947.210 241.160 947.990 241.300 ;
        RECT 947.210 241.100 947.530 241.160 ;
        RECT 947.670 241.100 947.990 241.160 ;
        RECT 947.670 203.560 947.990 203.620 ;
        RECT 947.475 203.420 947.990 203.560 ;
        RECT 947.670 203.360 947.990 203.420 ;
        RECT 947.670 138.280 947.990 138.340 ;
        RECT 947.475 138.140 947.990 138.280 ;
        RECT 947.670 138.080 947.990 138.140 ;
        RECT 946.290 48.520 946.610 48.580 ;
        RECT 947.670 48.520 947.990 48.580 ;
        RECT 946.290 48.380 947.990 48.520 ;
        RECT 946.290 48.320 946.610 48.380 ;
        RECT 947.670 48.320 947.990 48.380 ;
        RECT 294.010 26.760 294.330 26.820 ;
        RECT 946.750 26.760 947.070 26.820 ;
        RECT 294.010 26.620 947.070 26.760 ;
        RECT 294.010 26.560 294.330 26.620 ;
        RECT 946.750 26.560 947.070 26.620 ;
      LAYER via ;
        RECT 946.780 1062.540 947.040 1062.800 ;
        RECT 950.920 1062.540 951.180 1062.800 ;
        RECT 947.240 931.640 947.500 931.900 ;
        RECT 947.700 930.960 947.960 931.220 ;
        RECT 947.240 862.620 947.500 862.880 ;
        RECT 947.700 862.620 947.960 862.880 ;
        RECT 946.780 820.800 947.040 821.060 ;
        RECT 947.240 820.800 947.500 821.060 ;
        RECT 946.780 738.520 947.040 738.780 ;
        RECT 946.780 737.840 947.040 738.100 ;
        RECT 946.780 641.620 947.040 641.880 ;
        RECT 947.240 641.280 947.500 641.540 ;
        RECT 946.780 579.400 947.040 579.660 ;
        RECT 947.240 579.400 947.500 579.660 ;
        RECT 946.780 379.480 947.040 379.740 ;
        RECT 947.240 379.480 947.500 379.740 ;
        RECT 947.240 241.100 947.500 241.360 ;
        RECT 947.700 241.100 947.960 241.360 ;
        RECT 947.700 203.360 947.960 203.620 ;
        RECT 947.700 138.080 947.960 138.340 ;
        RECT 946.320 48.320 946.580 48.580 ;
        RECT 947.700 48.320 947.960 48.580 ;
        RECT 294.040 26.560 294.300 26.820 ;
        RECT 946.780 26.560 947.040 26.820 ;
      LAYER met2 ;
        RECT 950.830 1100.580 951.110 1104.000 ;
        RECT 950.830 1100.000 951.120 1100.580 ;
        RECT 950.980 1062.830 951.120 1100.000 ;
        RECT 946.780 1062.510 947.040 1062.830 ;
        RECT 950.920 1062.510 951.180 1062.830 ;
        RECT 946.840 1027.890 946.980 1062.510 ;
        RECT 946.840 1027.750 947.440 1027.890 ;
        RECT 947.300 931.930 947.440 1027.750 ;
        RECT 947.240 931.610 947.500 931.930 ;
        RECT 947.700 930.930 947.960 931.250 ;
        RECT 947.760 862.910 947.900 930.930 ;
        RECT 947.240 862.590 947.500 862.910 ;
        RECT 947.700 862.590 947.960 862.910 ;
        RECT 947.300 821.090 947.440 862.590 ;
        RECT 946.780 820.770 947.040 821.090 ;
        RECT 947.240 820.770 947.500 821.090 ;
        RECT 946.840 738.810 946.980 820.770 ;
        RECT 946.780 738.490 947.040 738.810 ;
        RECT 946.780 737.810 947.040 738.130 ;
        RECT 946.840 641.910 946.980 737.810 ;
        RECT 946.780 641.590 947.040 641.910 ;
        RECT 947.240 641.250 947.500 641.570 ;
        RECT 947.300 580.565 947.440 641.250 ;
        RECT 947.230 580.195 947.510 580.565 ;
        RECT 946.770 579.515 947.050 579.885 ;
        RECT 946.780 579.370 947.040 579.515 ;
        RECT 947.240 579.370 947.500 579.690 ;
        RECT 947.300 497.490 947.440 579.370 ;
        RECT 947.300 497.350 947.900 497.490 ;
        RECT 947.760 496.810 947.900 497.350 ;
        RECT 947.300 496.670 947.900 496.810 ;
        RECT 947.300 379.770 947.440 496.670 ;
        RECT 946.780 379.450 947.040 379.770 ;
        RECT 947.240 379.450 947.500 379.770 ;
        RECT 946.840 265.610 946.980 379.450 ;
        RECT 946.840 265.470 947.440 265.610 ;
        RECT 947.300 241.390 947.440 265.470 ;
        RECT 947.240 241.070 947.500 241.390 ;
        RECT 947.700 241.070 947.960 241.390 ;
        RECT 947.760 203.650 947.900 241.070 ;
        RECT 947.700 203.330 947.960 203.650 ;
        RECT 947.700 138.050 947.960 138.370 ;
        RECT 947.760 48.610 947.900 138.050 ;
        RECT 946.320 48.290 946.580 48.610 ;
        RECT 947.700 48.290 947.960 48.610 ;
        RECT 946.380 48.010 946.520 48.290 ;
        RECT 946.380 47.870 946.980 48.010 ;
        RECT 946.840 26.850 946.980 47.870 ;
        RECT 294.040 26.530 294.300 26.850 ;
        RECT 946.780 26.530 947.040 26.850 ;
        RECT 294.100 2.000 294.240 26.530 ;
        RECT 293.890 -4.000 294.450 2.000 ;
      LAYER via2 ;
        RECT 947.230 580.240 947.510 580.520 ;
        RECT 946.770 579.560 947.050 579.840 ;
      LAYER met3 ;
        RECT 947.205 580.530 947.535 580.545 ;
        RECT 946.990 580.215 947.535 580.530 ;
        RECT 946.990 579.865 947.290 580.215 ;
        RECT 946.745 579.550 947.290 579.865 ;
        RECT 946.745 579.535 947.075 579.550 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 311.950 27.100 312.270 27.160 ;
        RECT 953.190 27.100 953.510 27.160 ;
        RECT 311.950 26.960 953.510 27.100 ;
        RECT 311.950 26.900 312.270 26.960 ;
        RECT 953.190 26.900 953.510 26.960 ;
      LAYER via ;
        RECT 311.980 26.900 312.240 27.160 ;
        RECT 953.220 26.900 953.480 27.160 ;
      LAYER met2 ;
        RECT 956.810 1100.650 957.090 1104.000 ;
        RECT 955.580 1100.510 957.090 1100.650 ;
        RECT 955.580 1052.370 955.720 1100.510 ;
        RECT 956.810 1100.000 957.090 1100.510 ;
        RECT 953.280 1052.230 955.720 1052.370 ;
        RECT 953.280 27.190 953.420 1052.230 ;
        RECT 311.980 26.870 312.240 27.190 ;
        RECT 953.220 26.870 953.480 27.190 ;
        RECT 312.040 2.000 312.180 26.870 ;
        RECT 311.830 -4.000 312.390 2.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 960.625 965.685 960.795 1007.335 ;
        RECT 961.085 880.345 961.255 910.775 ;
        RECT 961.085 766.105 961.255 783.955 ;
        RECT 961.545 551.905 961.715 613.955 ;
        RECT 961.545 331.245 961.715 420.835 ;
        RECT 960.625 48.365 960.795 96.475 ;
      LAYER mcon ;
        RECT 960.625 1007.165 960.795 1007.335 ;
        RECT 961.085 910.605 961.255 910.775 ;
        RECT 961.085 783.785 961.255 783.955 ;
        RECT 961.545 613.785 961.715 613.955 ;
        RECT 961.545 420.665 961.715 420.835 ;
        RECT 960.625 96.305 960.795 96.475 ;
      LAYER met1 ;
        RECT 961.930 1062.740 962.250 1062.800 ;
        RECT 963.310 1062.740 963.630 1062.800 ;
        RECT 961.930 1062.600 963.630 1062.740 ;
        RECT 961.930 1062.540 962.250 1062.600 ;
        RECT 963.310 1062.540 963.630 1062.600 ;
        RECT 960.565 1007.320 960.855 1007.365 ;
        RECT 961.930 1007.320 962.250 1007.380 ;
        RECT 960.565 1007.180 962.250 1007.320 ;
        RECT 960.565 1007.135 960.855 1007.180 ;
        RECT 961.930 1007.120 962.250 1007.180 ;
        RECT 960.550 965.840 960.870 965.900 ;
        RECT 960.355 965.700 960.870 965.840 ;
        RECT 960.550 965.640 960.870 965.700 ;
        RECT 960.550 917.900 960.870 917.960 ;
        RECT 961.010 917.900 961.330 917.960 ;
        RECT 960.550 917.760 961.330 917.900 ;
        RECT 960.550 917.700 960.870 917.760 ;
        RECT 961.010 917.700 961.330 917.760 ;
        RECT 961.010 910.760 961.330 910.820 ;
        RECT 960.815 910.620 961.330 910.760 ;
        RECT 961.010 910.560 961.330 910.620 ;
        RECT 961.010 880.500 961.330 880.560 ;
        RECT 960.815 880.360 961.330 880.500 ;
        RECT 961.010 880.300 961.330 880.360 ;
        RECT 961.010 783.940 961.330 784.000 ;
        RECT 960.815 783.800 961.330 783.940 ;
        RECT 961.010 783.740 961.330 783.800 ;
        RECT 960.550 766.260 960.870 766.320 ;
        RECT 961.025 766.260 961.315 766.305 ;
        RECT 960.550 766.120 961.315 766.260 ;
        RECT 960.550 766.060 960.870 766.120 ;
        RECT 961.025 766.075 961.315 766.120 ;
        RECT 961.010 620.740 961.330 620.800 ;
        RECT 961.470 620.740 961.790 620.800 ;
        RECT 961.010 620.600 961.790 620.740 ;
        RECT 961.010 620.540 961.330 620.600 ;
        RECT 961.470 620.540 961.790 620.600 ;
        RECT 961.470 613.940 961.790 614.000 ;
        RECT 961.275 613.800 961.790 613.940 ;
        RECT 961.470 613.740 961.790 613.800 ;
        RECT 961.485 552.060 961.775 552.105 ;
        RECT 961.930 552.060 962.250 552.120 ;
        RECT 961.485 551.920 962.250 552.060 ;
        RECT 961.485 551.875 961.775 551.920 ;
        RECT 961.930 551.860 962.250 551.920 ;
        RECT 961.930 476.040 962.250 476.300 ;
        RECT 962.020 475.620 962.160 476.040 ;
        RECT 961.930 475.360 962.250 475.620 ;
        RECT 960.550 452.100 960.870 452.160 ;
        RECT 961.930 452.100 962.250 452.160 ;
        RECT 960.550 451.960 962.250 452.100 ;
        RECT 960.550 451.900 960.870 451.960 ;
        RECT 961.930 451.900 962.250 451.960 ;
        RECT 961.010 420.820 961.330 420.880 ;
        RECT 961.485 420.820 961.775 420.865 ;
        RECT 961.010 420.680 961.775 420.820 ;
        RECT 961.010 420.620 961.330 420.680 ;
        RECT 961.485 420.635 961.775 420.680 ;
        RECT 961.010 331.400 961.330 331.460 ;
        RECT 961.485 331.400 961.775 331.445 ;
        RECT 961.010 331.260 961.775 331.400 ;
        RECT 961.010 331.200 961.330 331.260 ;
        RECT 961.485 331.215 961.775 331.260 ;
        RECT 961.010 255.580 961.330 255.640 ;
        RECT 960.640 255.440 961.330 255.580 ;
        RECT 960.640 255.300 960.780 255.440 ;
        RECT 961.010 255.380 961.330 255.440 ;
        RECT 960.550 255.040 960.870 255.300 ;
        RECT 960.565 96.460 960.855 96.505 ;
        RECT 961.010 96.460 961.330 96.520 ;
        RECT 960.565 96.320 961.330 96.460 ;
        RECT 960.565 96.275 960.855 96.320 ;
        RECT 961.010 96.260 961.330 96.320 ;
        RECT 960.550 48.520 960.870 48.580 ;
        RECT 960.355 48.380 960.870 48.520 ;
        RECT 960.550 48.320 960.870 48.380 ;
        RECT 329.890 27.440 330.210 27.500 ;
        RECT 960.550 27.440 960.870 27.500 ;
        RECT 329.890 27.300 960.870 27.440 ;
        RECT 329.890 27.240 330.210 27.300 ;
        RECT 960.550 27.240 960.870 27.300 ;
      LAYER via ;
        RECT 961.960 1062.540 962.220 1062.800 ;
        RECT 963.340 1062.540 963.600 1062.800 ;
        RECT 961.960 1007.120 962.220 1007.380 ;
        RECT 960.580 965.640 960.840 965.900 ;
        RECT 960.580 917.700 960.840 917.960 ;
        RECT 961.040 917.700 961.300 917.960 ;
        RECT 961.040 910.560 961.300 910.820 ;
        RECT 961.040 880.300 961.300 880.560 ;
        RECT 961.040 783.740 961.300 784.000 ;
        RECT 960.580 766.060 960.840 766.320 ;
        RECT 961.040 620.540 961.300 620.800 ;
        RECT 961.500 620.540 961.760 620.800 ;
        RECT 961.500 613.740 961.760 614.000 ;
        RECT 961.960 551.860 962.220 552.120 ;
        RECT 961.960 476.040 962.220 476.300 ;
        RECT 961.960 475.360 962.220 475.620 ;
        RECT 960.580 451.900 960.840 452.160 ;
        RECT 961.960 451.900 962.220 452.160 ;
        RECT 961.040 420.620 961.300 420.880 ;
        RECT 961.040 331.200 961.300 331.460 ;
        RECT 961.040 255.380 961.300 255.640 ;
        RECT 960.580 255.040 960.840 255.300 ;
        RECT 961.040 96.260 961.300 96.520 ;
        RECT 960.580 48.320 960.840 48.580 ;
        RECT 329.920 27.240 330.180 27.500 ;
        RECT 960.580 27.240 960.840 27.500 ;
      LAYER met2 ;
        RECT 963.250 1100.580 963.530 1104.000 ;
        RECT 963.250 1100.000 963.540 1100.580 ;
        RECT 963.400 1062.830 963.540 1100.000 ;
        RECT 961.960 1062.510 962.220 1062.830 ;
        RECT 963.340 1062.510 963.600 1062.830 ;
        RECT 962.020 1007.410 962.160 1062.510 ;
        RECT 961.960 1007.090 962.220 1007.410 ;
        RECT 960.580 965.610 960.840 965.930 ;
        RECT 960.640 917.990 960.780 965.610 ;
        RECT 960.580 917.670 960.840 917.990 ;
        RECT 961.040 917.670 961.300 917.990 ;
        RECT 961.100 910.850 961.240 917.670 ;
        RECT 961.040 910.530 961.300 910.850 ;
        RECT 961.040 880.270 961.300 880.590 ;
        RECT 961.100 784.030 961.240 880.270 ;
        RECT 961.040 783.710 961.300 784.030 ;
        RECT 960.580 766.090 960.840 766.350 ;
        RECT 960.580 766.030 961.240 766.090 ;
        RECT 960.640 765.950 961.240 766.030 ;
        RECT 961.100 620.830 961.240 765.950 ;
        RECT 961.040 620.510 961.300 620.830 ;
        RECT 961.500 620.510 961.760 620.830 ;
        RECT 961.560 614.030 961.700 620.510 ;
        RECT 961.500 613.710 961.760 614.030 ;
        RECT 961.960 551.830 962.220 552.150 ;
        RECT 962.020 476.330 962.160 551.830 ;
        RECT 961.960 476.010 962.220 476.330 ;
        RECT 961.960 475.330 962.220 475.650 ;
        RECT 962.020 452.190 962.160 475.330 ;
        RECT 960.580 451.870 960.840 452.190 ;
        RECT 961.960 451.870 962.220 452.190 ;
        RECT 960.640 428.130 960.780 451.870 ;
        RECT 960.640 427.990 961.240 428.130 ;
        RECT 961.100 420.910 961.240 427.990 ;
        RECT 961.040 420.590 961.300 420.910 ;
        RECT 961.040 331.170 961.300 331.490 ;
        RECT 961.100 255.670 961.240 331.170 ;
        RECT 961.040 255.350 961.300 255.670 ;
        RECT 960.580 255.010 960.840 255.330 ;
        RECT 960.640 210.530 960.780 255.010 ;
        RECT 960.640 210.390 961.700 210.530 ;
        RECT 961.560 130.290 961.700 210.390 ;
        RECT 961.100 130.150 961.700 130.290 ;
        RECT 961.100 96.550 961.240 130.150 ;
        RECT 961.040 96.230 961.300 96.550 ;
        RECT 960.580 48.290 960.840 48.610 ;
        RECT 960.640 27.530 960.780 48.290 ;
        RECT 329.920 27.210 330.180 27.530 ;
        RECT 960.580 27.210 960.840 27.530 ;
        RECT 329.980 2.000 330.120 27.210 ;
        RECT 329.770 -4.000 330.330 2.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 347.370 23.700 347.690 23.760 ;
        RECT 967.450 23.700 967.770 23.760 ;
        RECT 347.370 23.560 967.770 23.700 ;
        RECT 347.370 23.500 347.690 23.560 ;
        RECT 967.450 23.500 967.770 23.560 ;
      LAYER via ;
        RECT 347.400 23.500 347.660 23.760 ;
        RECT 967.480 23.500 967.740 23.760 ;
      LAYER met2 ;
        RECT 969.230 1100.650 969.510 1104.000 ;
        RECT 967.540 1100.510 969.510 1100.650 ;
        RECT 967.540 23.790 967.680 1100.510 ;
        RECT 969.230 1100.000 969.510 1100.510 ;
        RECT 347.400 23.470 347.660 23.790 ;
        RECT 967.480 23.470 967.740 23.790 ;
        RECT 347.460 2.000 347.600 23.470 ;
        RECT 347.250 -4.000 347.810 2.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 365.310 33.900 365.630 33.960 ;
        RECT 973.890 33.900 974.210 33.960 ;
        RECT 365.310 33.760 974.210 33.900 ;
        RECT 365.310 33.700 365.630 33.760 ;
        RECT 973.890 33.700 974.210 33.760 ;
      LAYER via ;
        RECT 365.340 33.700 365.600 33.960 ;
        RECT 973.920 33.700 974.180 33.960 ;
      LAYER met2 ;
        RECT 975.210 1100.650 975.490 1104.000 ;
        RECT 973.980 1100.510 975.490 1100.650 ;
        RECT 973.980 33.990 974.120 1100.510 ;
        RECT 975.210 1100.000 975.490 1100.510 ;
        RECT 365.340 33.670 365.600 33.990 ;
        RECT 973.920 33.670 974.180 33.990 ;
        RECT 365.400 2.000 365.540 33.670 ;
        RECT 365.190 -4.000 365.750 2.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 383.250 39.000 383.570 39.060 ;
        RECT 980.790 39.000 981.110 39.060 ;
        RECT 383.250 38.860 981.110 39.000 ;
        RECT 383.250 38.800 383.570 38.860 ;
        RECT 980.790 38.800 981.110 38.860 ;
      LAYER via ;
        RECT 383.280 38.800 383.540 39.060 ;
        RECT 980.820 38.800 981.080 39.060 ;
      LAYER met2 ;
        RECT 981.190 1100.650 981.470 1104.000 ;
        RECT 980.880 1100.510 981.470 1100.650 ;
        RECT 980.880 39.090 981.020 1100.510 ;
        RECT 981.190 1100.000 981.470 1100.510 ;
        RECT 383.280 38.770 383.540 39.090 ;
        RECT 980.820 38.770 981.080 39.090 ;
        RECT 383.340 2.000 383.480 38.770 ;
        RECT 383.130 -4.000 383.690 2.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 401.190 39.340 401.510 39.400 ;
        RECT 987.690 39.340 988.010 39.400 ;
        RECT 401.190 39.200 988.010 39.340 ;
        RECT 401.190 39.140 401.510 39.200 ;
        RECT 987.690 39.140 988.010 39.200 ;
      LAYER via ;
        RECT 401.220 39.140 401.480 39.400 ;
        RECT 987.720 39.140 987.980 39.400 ;
      LAYER met2 ;
        RECT 987.630 1100.580 987.910 1104.000 ;
        RECT 987.630 1100.000 987.920 1100.580 ;
        RECT 987.780 39.430 987.920 1100.000 ;
        RECT 401.220 39.110 401.480 39.430 ;
        RECT 987.720 39.110 987.980 39.430 ;
        RECT 401.280 2.000 401.420 39.110 ;
        RECT 401.070 -4.000 401.630 2.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 62.170 25.060 62.490 25.120 ;
        RECT 870.390 25.060 870.710 25.120 ;
        RECT 62.170 24.920 870.710 25.060 ;
        RECT 62.170 24.860 62.490 24.920 ;
        RECT 870.390 24.860 870.710 24.920 ;
      LAYER via ;
        RECT 62.200 24.860 62.460 25.120 ;
        RECT 870.420 24.860 870.680 25.120 ;
      LAYER met2 ;
        RECT 871.250 1100.650 871.530 1104.000 ;
        RECT 870.480 1100.510 871.530 1100.650 ;
        RECT 870.480 25.150 870.620 1100.510 ;
        RECT 871.250 1100.000 871.530 1100.510 ;
        RECT 62.200 24.830 62.460 25.150 ;
        RECT 870.420 24.830 870.680 25.150 ;
        RECT 62.260 2.000 62.400 24.830 ;
        RECT 62.050 -4.000 62.610 2.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 419.130 39.680 419.450 39.740 ;
        RECT 993.670 39.680 993.990 39.740 ;
        RECT 419.130 39.540 993.990 39.680 ;
        RECT 419.130 39.480 419.450 39.540 ;
        RECT 993.670 39.480 993.990 39.540 ;
      LAYER via ;
        RECT 419.160 39.480 419.420 39.740 ;
        RECT 993.700 39.480 993.960 39.740 ;
      LAYER met2 ;
        RECT 993.610 1100.580 993.890 1104.000 ;
        RECT 993.610 1100.000 993.900 1100.580 ;
        RECT 993.760 39.770 993.900 1100.000 ;
        RECT 419.160 39.450 419.420 39.770 ;
        RECT 993.700 39.450 993.960 39.770 ;
        RECT 419.220 2.000 419.360 39.450 ;
        RECT 419.010 -4.000 419.570 2.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 994.130 1041.660 994.450 1041.720 ;
        RECT 998.270 1041.660 998.590 1041.720 ;
        RECT 994.130 1041.520 998.590 1041.660 ;
        RECT 994.130 1041.460 994.450 1041.520 ;
        RECT 998.270 1041.460 998.590 1041.520 ;
        RECT 436.610 40.020 436.930 40.080 ;
        RECT 994.130 40.020 994.450 40.080 ;
        RECT 436.610 39.880 994.450 40.020 ;
        RECT 436.610 39.820 436.930 39.880 ;
        RECT 994.130 39.820 994.450 39.880 ;
      LAYER via ;
        RECT 994.160 1041.460 994.420 1041.720 ;
        RECT 998.300 1041.460 998.560 1041.720 ;
        RECT 436.640 39.820 436.900 40.080 ;
        RECT 994.160 39.820 994.420 40.080 ;
      LAYER met2 ;
        RECT 999.590 1100.650 999.870 1104.000 ;
        RECT 998.360 1100.510 999.870 1100.650 ;
        RECT 998.360 1041.750 998.500 1100.510 ;
        RECT 999.590 1100.000 999.870 1100.510 ;
        RECT 994.160 1041.430 994.420 1041.750 ;
        RECT 998.300 1041.430 998.560 1041.750 ;
        RECT 994.220 40.110 994.360 1041.430 ;
        RECT 436.640 39.790 436.900 40.110 ;
        RECT 994.160 39.790 994.420 40.110 ;
        RECT 436.700 2.000 436.840 39.790 ;
        RECT 436.490 -4.000 437.050 2.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1001.565 579.105 1001.735 620.755 ;
        RECT 1002.025 241.485 1002.195 307.275 ;
        RECT 1002.025 131.325 1002.195 138.295 ;
      LAYER mcon ;
        RECT 1001.565 620.585 1001.735 620.755 ;
        RECT 1002.025 307.105 1002.195 307.275 ;
        RECT 1002.025 138.125 1002.195 138.295 ;
      LAYER met1 ;
        RECT 1004.250 1062.740 1004.570 1062.800 ;
        RECT 1006.090 1062.740 1006.410 1062.800 ;
        RECT 1004.250 1062.600 1006.410 1062.740 ;
        RECT 1004.250 1062.540 1004.570 1062.600 ;
        RECT 1006.090 1062.540 1006.410 1062.600 ;
        RECT 1001.950 738.520 1002.270 738.780 ;
        RECT 1002.040 738.100 1002.180 738.520 ;
        RECT 1001.950 737.840 1002.270 738.100 ;
        RECT 1001.490 620.740 1001.810 620.800 ;
        RECT 1001.295 620.600 1001.810 620.740 ;
        RECT 1001.490 620.540 1001.810 620.600 ;
        RECT 1001.505 579.260 1001.795 579.305 ;
        RECT 1002.870 579.260 1003.190 579.320 ;
        RECT 1001.505 579.120 1003.190 579.260 ;
        RECT 1001.505 579.075 1001.795 579.120 ;
        RECT 1002.870 579.060 1003.190 579.120 ;
        RECT 1001.950 428.300 1002.270 428.360 ;
        RECT 1001.580 428.160 1002.270 428.300 ;
        RECT 1001.580 428.020 1001.720 428.160 ;
        RECT 1001.950 428.100 1002.270 428.160 ;
        RECT 1001.490 427.760 1001.810 428.020 ;
        RECT 1001.490 386.480 1001.810 386.540 ;
        RECT 1001.950 386.480 1002.270 386.540 ;
        RECT 1001.490 386.340 1002.270 386.480 ;
        RECT 1001.490 386.280 1001.810 386.340 ;
        RECT 1001.950 386.280 1002.270 386.340 ;
        RECT 1001.950 307.260 1002.270 307.320 ;
        RECT 1001.755 307.120 1002.270 307.260 ;
        RECT 1001.950 307.060 1002.270 307.120 ;
        RECT 1001.965 241.640 1002.255 241.685 ;
        RECT 1002.410 241.640 1002.730 241.700 ;
        RECT 1001.965 241.500 1002.730 241.640 ;
        RECT 1001.965 241.455 1002.255 241.500 ;
        RECT 1002.410 241.440 1002.730 241.500 ;
        RECT 1001.950 186.560 1002.270 186.620 ;
        RECT 1002.410 186.560 1002.730 186.620 ;
        RECT 1001.950 186.420 1002.730 186.560 ;
        RECT 1001.950 186.360 1002.270 186.420 ;
        RECT 1002.410 186.360 1002.730 186.420 ;
        RECT 1001.950 138.280 1002.270 138.340 ;
        RECT 1001.755 138.140 1002.270 138.280 ;
        RECT 1001.950 138.080 1002.270 138.140 ;
        RECT 1001.950 131.480 1002.270 131.540 ;
        RECT 1001.755 131.340 1002.270 131.480 ;
        RECT 1001.950 131.280 1002.270 131.340 ;
        RECT 1001.950 110.540 1002.270 110.800 ;
        RECT 1002.040 110.120 1002.180 110.540 ;
        RECT 1001.950 109.860 1002.270 110.120 ;
        RECT 454.550 40.360 454.870 40.420 ;
        RECT 1001.950 40.360 1002.270 40.420 ;
        RECT 454.550 40.220 1002.270 40.360 ;
        RECT 454.550 40.160 454.870 40.220 ;
        RECT 1001.950 40.160 1002.270 40.220 ;
      LAYER via ;
        RECT 1004.280 1062.540 1004.540 1062.800 ;
        RECT 1006.120 1062.540 1006.380 1062.800 ;
        RECT 1001.980 738.520 1002.240 738.780 ;
        RECT 1001.980 737.840 1002.240 738.100 ;
        RECT 1001.520 620.540 1001.780 620.800 ;
        RECT 1002.900 579.060 1003.160 579.320 ;
        RECT 1001.980 428.100 1002.240 428.360 ;
        RECT 1001.520 427.760 1001.780 428.020 ;
        RECT 1001.520 386.280 1001.780 386.540 ;
        RECT 1001.980 386.280 1002.240 386.540 ;
        RECT 1001.980 307.060 1002.240 307.320 ;
        RECT 1002.440 241.440 1002.700 241.700 ;
        RECT 1001.980 186.360 1002.240 186.620 ;
        RECT 1002.440 186.360 1002.700 186.620 ;
        RECT 1001.980 138.080 1002.240 138.340 ;
        RECT 1001.980 131.280 1002.240 131.540 ;
        RECT 1001.980 110.540 1002.240 110.800 ;
        RECT 1001.980 109.860 1002.240 110.120 ;
        RECT 454.580 40.160 454.840 40.420 ;
        RECT 1001.980 40.160 1002.240 40.420 ;
      LAYER met2 ;
        RECT 1006.030 1100.580 1006.310 1104.000 ;
        RECT 1006.030 1100.000 1006.320 1100.580 ;
        RECT 1006.180 1062.830 1006.320 1100.000 ;
        RECT 1004.280 1062.510 1004.540 1062.830 ;
        RECT 1006.120 1062.510 1006.380 1062.830 ;
        RECT 1004.340 990.490 1004.480 1062.510 ;
        RECT 1002.500 990.350 1004.480 990.490 ;
        RECT 1002.500 883.730 1002.640 990.350 ;
        RECT 1002.040 883.590 1002.640 883.730 ;
        RECT 1002.040 773.685 1002.180 883.590 ;
        RECT 1001.970 773.315 1002.250 773.685 ;
        RECT 1001.970 772.635 1002.250 773.005 ;
        RECT 1002.040 738.810 1002.180 772.635 ;
        RECT 1001.980 738.490 1002.240 738.810 ;
        RECT 1001.980 737.810 1002.240 738.130 ;
        RECT 1002.040 677.125 1002.180 737.810 ;
        RECT 1001.970 676.755 1002.250 677.125 ;
        RECT 1001.970 676.075 1002.250 676.445 ;
        RECT 1002.040 645.050 1002.180 676.075 ;
        RECT 1001.580 644.910 1002.180 645.050 ;
        RECT 1001.580 620.830 1001.720 644.910 ;
        RECT 1001.520 620.510 1001.780 620.830 ;
        RECT 1002.900 579.030 1003.160 579.350 ;
        RECT 1002.960 483.325 1003.100 579.030 ;
        RECT 1001.970 482.955 1002.250 483.325 ;
        RECT 1002.890 482.955 1003.170 483.325 ;
        RECT 1002.040 428.390 1002.180 482.955 ;
        RECT 1001.980 428.070 1002.240 428.390 ;
        RECT 1001.520 427.730 1001.780 428.050 ;
        RECT 1001.580 386.570 1001.720 427.730 ;
        RECT 1001.520 386.250 1001.780 386.570 ;
        RECT 1001.980 386.250 1002.240 386.570 ;
        RECT 1002.040 307.350 1002.180 386.250 ;
        RECT 1001.980 307.030 1002.240 307.350 ;
        RECT 1002.440 241.410 1002.700 241.730 ;
        RECT 1002.500 186.650 1002.640 241.410 ;
        RECT 1001.980 186.330 1002.240 186.650 ;
        RECT 1002.440 186.330 1002.700 186.650 ;
        RECT 1002.040 138.370 1002.180 186.330 ;
        RECT 1001.980 138.050 1002.240 138.370 ;
        RECT 1001.980 131.250 1002.240 131.570 ;
        RECT 1002.040 110.830 1002.180 131.250 ;
        RECT 1001.980 110.510 1002.240 110.830 ;
        RECT 1001.980 109.830 1002.240 110.150 ;
        RECT 1002.040 40.450 1002.180 109.830 ;
        RECT 454.580 40.130 454.840 40.450 ;
        RECT 1001.980 40.130 1002.240 40.450 ;
        RECT 454.640 2.000 454.780 40.130 ;
        RECT 454.430 -4.000 454.990 2.000 ;
      LAYER via2 ;
        RECT 1001.970 773.360 1002.250 773.640 ;
        RECT 1001.970 772.680 1002.250 772.960 ;
        RECT 1001.970 676.800 1002.250 677.080 ;
        RECT 1001.970 676.120 1002.250 676.400 ;
        RECT 1001.970 483.000 1002.250 483.280 ;
        RECT 1002.890 483.000 1003.170 483.280 ;
      LAYER met3 ;
        RECT 1001.945 773.650 1002.275 773.665 ;
        RECT 1001.270 773.350 1002.275 773.650 ;
        RECT 1001.270 772.970 1001.570 773.350 ;
        RECT 1001.945 773.335 1002.275 773.350 ;
        RECT 1001.945 772.970 1002.275 772.985 ;
        RECT 1001.270 772.670 1002.275 772.970 ;
        RECT 1001.945 772.655 1002.275 772.670 ;
        RECT 1001.945 677.090 1002.275 677.105 ;
        RECT 1001.945 676.775 1002.490 677.090 ;
        RECT 1002.190 676.425 1002.490 676.775 ;
        RECT 1001.945 676.110 1002.490 676.425 ;
        RECT 1001.945 676.095 1002.275 676.110 ;
        RECT 1001.945 483.290 1002.275 483.305 ;
        RECT 1002.865 483.290 1003.195 483.305 ;
        RECT 1001.945 482.990 1003.195 483.290 ;
        RECT 1001.945 482.975 1002.275 482.990 ;
        RECT 1002.865 482.975 1003.195 482.990 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1008.925 620.925 1009.095 669.375 ;
        RECT 1009.385 524.365 1009.555 572.475 ;
        RECT 1009.385 386.325 1009.555 434.775 ;
        RECT 1009.385 269.705 1009.555 307.275 ;
        RECT 1009.385 138.125 1009.555 227.715 ;
      LAYER mcon ;
        RECT 1008.925 669.205 1009.095 669.375 ;
        RECT 1009.385 572.305 1009.555 572.475 ;
        RECT 1009.385 434.605 1009.555 434.775 ;
        RECT 1009.385 307.105 1009.555 307.275 ;
        RECT 1009.385 227.545 1009.555 227.715 ;
      LAYER met1 ;
        RECT 1009.310 1062.740 1009.630 1062.800 ;
        RECT 1012.070 1062.740 1012.390 1062.800 ;
        RECT 1009.310 1062.600 1012.390 1062.740 ;
        RECT 1009.310 1062.540 1009.630 1062.600 ;
        RECT 1012.070 1062.540 1012.390 1062.600 ;
        RECT 1009.310 738.520 1009.630 738.780 ;
        RECT 1009.400 738.100 1009.540 738.520 ;
        RECT 1009.310 737.840 1009.630 738.100 ;
        RECT 1008.865 669.360 1009.155 669.405 ;
        RECT 1009.310 669.360 1009.630 669.420 ;
        RECT 1008.865 669.220 1009.630 669.360 ;
        RECT 1008.865 669.175 1009.155 669.220 ;
        RECT 1009.310 669.160 1009.630 669.220 ;
        RECT 1008.850 621.080 1009.170 621.140 ;
        RECT 1008.655 620.940 1009.170 621.080 ;
        RECT 1008.850 620.880 1009.170 620.940 ;
        RECT 1008.850 579.940 1009.170 580.000 ;
        RECT 1009.310 579.940 1009.630 580.000 ;
        RECT 1008.850 579.800 1009.630 579.940 ;
        RECT 1008.850 579.740 1009.170 579.800 ;
        RECT 1009.310 579.740 1009.630 579.800 ;
        RECT 1009.310 572.460 1009.630 572.520 ;
        RECT 1009.115 572.320 1009.630 572.460 ;
        RECT 1009.310 572.260 1009.630 572.320 ;
        RECT 1009.325 524.520 1009.615 524.565 ;
        RECT 1010.230 524.520 1010.550 524.580 ;
        RECT 1009.325 524.380 1010.550 524.520 ;
        RECT 1009.325 524.335 1009.615 524.380 ;
        RECT 1010.230 524.320 1010.550 524.380 ;
        RECT 1009.310 434.760 1009.630 434.820 ;
        RECT 1009.115 434.620 1009.630 434.760 ;
        RECT 1009.310 434.560 1009.630 434.620 ;
        RECT 1009.310 386.480 1009.630 386.540 ;
        RECT 1009.115 386.340 1009.630 386.480 ;
        RECT 1009.310 386.280 1009.630 386.340 ;
        RECT 1009.310 307.260 1009.630 307.320 ;
        RECT 1009.115 307.120 1009.630 307.260 ;
        RECT 1009.310 307.060 1009.630 307.120 ;
        RECT 1009.325 269.860 1009.615 269.905 ;
        RECT 1010.230 269.860 1010.550 269.920 ;
        RECT 1009.325 269.720 1010.550 269.860 ;
        RECT 1009.325 269.675 1009.615 269.720 ;
        RECT 1010.230 269.660 1010.550 269.720 ;
        RECT 1009.325 227.700 1009.615 227.745 ;
        RECT 1009.770 227.700 1010.090 227.760 ;
        RECT 1009.325 227.560 1010.090 227.700 ;
        RECT 1009.325 227.515 1009.615 227.560 ;
        RECT 1009.770 227.500 1010.090 227.560 ;
        RECT 1009.310 138.280 1009.630 138.340 ;
        RECT 1009.115 138.140 1009.630 138.280 ;
        RECT 1009.310 138.080 1009.630 138.140 ;
        RECT 472.490 40.700 472.810 40.760 ;
        RECT 1009.310 40.700 1009.630 40.760 ;
        RECT 472.490 40.560 1009.630 40.700 ;
        RECT 472.490 40.500 472.810 40.560 ;
        RECT 1009.310 40.500 1009.630 40.560 ;
      LAYER via ;
        RECT 1009.340 1062.540 1009.600 1062.800 ;
        RECT 1012.100 1062.540 1012.360 1062.800 ;
        RECT 1009.340 738.520 1009.600 738.780 ;
        RECT 1009.340 737.840 1009.600 738.100 ;
        RECT 1009.340 669.160 1009.600 669.420 ;
        RECT 1008.880 620.880 1009.140 621.140 ;
        RECT 1008.880 579.740 1009.140 580.000 ;
        RECT 1009.340 579.740 1009.600 580.000 ;
        RECT 1009.340 572.260 1009.600 572.520 ;
        RECT 1010.260 524.320 1010.520 524.580 ;
        RECT 1009.340 434.560 1009.600 434.820 ;
        RECT 1009.340 386.280 1009.600 386.540 ;
        RECT 1009.340 307.060 1009.600 307.320 ;
        RECT 1010.260 269.660 1010.520 269.920 ;
        RECT 1009.800 227.500 1010.060 227.760 ;
        RECT 1009.340 138.080 1009.600 138.340 ;
        RECT 472.520 40.500 472.780 40.760 ;
        RECT 1009.340 40.500 1009.600 40.760 ;
      LAYER met2 ;
        RECT 1012.010 1100.580 1012.290 1104.000 ;
        RECT 1012.010 1100.000 1012.300 1100.580 ;
        RECT 1012.160 1062.830 1012.300 1100.000 ;
        RECT 1009.340 1062.510 1009.600 1062.830 ;
        RECT 1012.100 1062.510 1012.360 1062.830 ;
        RECT 1009.400 1027.890 1009.540 1062.510 ;
        RECT 1009.400 1027.750 1010.000 1027.890 ;
        RECT 1009.860 883.730 1010.000 1027.750 ;
        RECT 1009.400 883.590 1010.000 883.730 ;
        RECT 1009.400 773.685 1009.540 883.590 ;
        RECT 1009.330 773.315 1009.610 773.685 ;
        RECT 1009.330 772.635 1009.610 773.005 ;
        RECT 1009.400 738.810 1009.540 772.635 ;
        RECT 1009.340 738.490 1009.600 738.810 ;
        RECT 1009.340 737.810 1009.600 738.130 ;
        RECT 1009.400 677.125 1009.540 737.810 ;
        RECT 1009.330 676.755 1009.610 677.125 ;
        RECT 1009.330 676.075 1009.610 676.445 ;
        RECT 1009.400 669.450 1009.540 676.075 ;
        RECT 1009.340 669.130 1009.600 669.450 ;
        RECT 1008.880 620.850 1009.140 621.170 ;
        RECT 1008.940 580.030 1009.080 620.850 ;
        RECT 1008.880 579.710 1009.140 580.030 ;
        RECT 1009.340 579.710 1009.600 580.030 ;
        RECT 1009.400 572.550 1009.540 579.710 ;
        RECT 1009.340 572.230 1009.600 572.550 ;
        RECT 1010.260 524.290 1010.520 524.610 ;
        RECT 1010.320 483.325 1010.460 524.290 ;
        RECT 1009.330 482.955 1009.610 483.325 ;
        RECT 1010.250 482.955 1010.530 483.325 ;
        RECT 1009.400 434.850 1009.540 482.955 ;
        RECT 1009.340 434.530 1009.600 434.850 ;
        RECT 1009.340 386.250 1009.600 386.570 ;
        RECT 1009.400 307.350 1009.540 386.250 ;
        RECT 1009.340 307.030 1009.600 307.350 ;
        RECT 1010.260 269.630 1010.520 269.950 ;
        RECT 1010.320 235.010 1010.460 269.630 ;
        RECT 1009.860 234.870 1010.460 235.010 ;
        RECT 1009.860 227.790 1010.000 234.870 ;
        RECT 1009.800 227.470 1010.060 227.790 ;
        RECT 1009.340 138.050 1009.600 138.370 ;
        RECT 1009.400 40.790 1009.540 138.050 ;
        RECT 472.520 40.470 472.780 40.790 ;
        RECT 1009.340 40.470 1009.600 40.790 ;
        RECT 472.580 2.000 472.720 40.470 ;
        RECT 472.370 -4.000 472.930 2.000 ;
      LAYER via2 ;
        RECT 1009.330 773.360 1009.610 773.640 ;
        RECT 1009.330 772.680 1009.610 772.960 ;
        RECT 1009.330 676.800 1009.610 677.080 ;
        RECT 1009.330 676.120 1009.610 676.400 ;
        RECT 1009.330 483.000 1009.610 483.280 ;
        RECT 1010.250 483.000 1010.530 483.280 ;
      LAYER met3 ;
        RECT 1009.305 773.650 1009.635 773.665 ;
        RECT 1008.630 773.350 1009.635 773.650 ;
        RECT 1008.630 772.970 1008.930 773.350 ;
        RECT 1009.305 773.335 1009.635 773.350 ;
        RECT 1009.305 772.970 1009.635 772.985 ;
        RECT 1008.630 772.670 1009.635 772.970 ;
        RECT 1009.305 772.655 1009.635 772.670 ;
        RECT 1009.305 677.090 1009.635 677.105 ;
        RECT 1009.305 676.775 1009.850 677.090 ;
        RECT 1009.550 676.425 1009.850 676.775 ;
        RECT 1009.305 676.110 1009.850 676.425 ;
        RECT 1009.305 676.095 1009.635 676.110 ;
        RECT 1009.305 483.290 1009.635 483.305 ;
        RECT 1010.225 483.290 1010.555 483.305 ;
        RECT 1009.305 482.990 1010.555 483.290 ;
        RECT 1009.305 482.975 1009.635 482.990 ;
        RECT 1010.225 482.975 1010.555 482.990 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1015.825 724.285 1015.995 807.075 ;
        RECT 1015.365 662.405 1015.535 670.055 ;
        RECT 1015.365 572.645 1015.535 620.755 ;
        RECT 1015.365 355.385 1015.535 403.495 ;
        RECT 1015.365 276.165 1015.535 324.275 ;
      LAYER mcon ;
        RECT 1015.825 806.905 1015.995 807.075 ;
        RECT 1015.365 669.885 1015.535 670.055 ;
        RECT 1015.365 620.585 1015.535 620.755 ;
        RECT 1015.365 403.325 1015.535 403.495 ;
        RECT 1015.365 324.105 1015.535 324.275 ;
      LAYER met1 ;
        RECT 1017.130 1062.740 1017.450 1062.800 ;
        RECT 1018.050 1062.740 1018.370 1062.800 ;
        RECT 1017.130 1062.600 1018.370 1062.740 ;
        RECT 1017.130 1062.540 1017.450 1062.600 ;
        RECT 1018.050 1062.540 1018.370 1062.600 ;
        RECT 1016.210 966.180 1016.530 966.240 ;
        RECT 1016.670 966.180 1016.990 966.240 ;
        RECT 1016.210 966.040 1016.990 966.180 ;
        RECT 1016.210 965.980 1016.530 966.040 ;
        RECT 1016.670 965.980 1016.990 966.040 ;
        RECT 1015.750 855.680 1016.070 855.740 ;
        RECT 1016.210 855.680 1016.530 855.740 ;
        RECT 1015.750 855.540 1016.530 855.680 ;
        RECT 1015.750 855.480 1016.070 855.540 ;
        RECT 1016.210 855.480 1016.530 855.540 ;
        RECT 1015.750 807.060 1016.070 807.120 ;
        RECT 1015.555 806.920 1016.070 807.060 ;
        RECT 1015.750 806.860 1016.070 806.920 ;
        RECT 1015.750 724.440 1016.070 724.500 ;
        RECT 1015.555 724.300 1016.070 724.440 ;
        RECT 1015.750 724.240 1016.070 724.300 ;
        RECT 1015.305 670.040 1015.595 670.085 ;
        RECT 1016.210 670.040 1016.530 670.100 ;
        RECT 1015.305 669.900 1016.530 670.040 ;
        RECT 1015.305 669.855 1015.595 669.900 ;
        RECT 1016.210 669.840 1016.530 669.900 ;
        RECT 1015.290 662.560 1015.610 662.620 ;
        RECT 1015.095 662.420 1015.610 662.560 ;
        RECT 1015.290 662.360 1015.610 662.420 ;
        RECT 1015.290 620.740 1015.610 620.800 ;
        RECT 1015.095 620.600 1015.610 620.740 ;
        RECT 1015.290 620.540 1015.610 620.600 ;
        RECT 1015.305 572.800 1015.595 572.845 ;
        RECT 1016.210 572.800 1016.530 572.860 ;
        RECT 1015.305 572.660 1016.530 572.800 ;
        RECT 1015.305 572.615 1015.595 572.660 ;
        RECT 1016.210 572.600 1016.530 572.660 ;
        RECT 1015.290 403.480 1015.610 403.540 ;
        RECT 1015.095 403.340 1015.610 403.480 ;
        RECT 1015.290 403.280 1015.610 403.340 ;
        RECT 1015.290 355.540 1015.610 355.600 ;
        RECT 1015.095 355.400 1015.610 355.540 ;
        RECT 1015.290 355.340 1015.610 355.400 ;
        RECT 1015.290 331.060 1015.610 331.120 ;
        RECT 1016.670 331.060 1016.990 331.120 ;
        RECT 1015.290 330.920 1016.990 331.060 ;
        RECT 1015.290 330.860 1015.610 330.920 ;
        RECT 1016.670 330.860 1016.990 330.920 ;
        RECT 1015.305 324.260 1015.595 324.305 ;
        RECT 1016.670 324.260 1016.990 324.320 ;
        RECT 1015.305 324.120 1016.990 324.260 ;
        RECT 1015.305 324.075 1015.595 324.120 ;
        RECT 1016.670 324.060 1016.990 324.120 ;
        RECT 1015.290 276.320 1015.610 276.380 ;
        RECT 1015.095 276.180 1015.610 276.320 ;
        RECT 1015.290 276.120 1015.610 276.180 ;
        RECT 1015.750 144.740 1016.070 144.800 ;
        RECT 1016.210 144.740 1016.530 144.800 ;
        RECT 1015.750 144.600 1016.530 144.740 ;
        RECT 1015.750 144.540 1016.070 144.600 ;
        RECT 1016.210 144.540 1016.530 144.600 ;
        RECT 490.430 41.040 490.750 41.100 ;
        RECT 1015.750 41.040 1016.070 41.100 ;
        RECT 490.430 40.900 1016.070 41.040 ;
        RECT 490.430 40.840 490.750 40.900 ;
        RECT 1015.750 40.840 1016.070 40.900 ;
      LAYER via ;
        RECT 1017.160 1062.540 1017.420 1062.800 ;
        RECT 1018.080 1062.540 1018.340 1062.800 ;
        RECT 1016.240 965.980 1016.500 966.240 ;
        RECT 1016.700 965.980 1016.960 966.240 ;
        RECT 1015.780 855.480 1016.040 855.740 ;
        RECT 1016.240 855.480 1016.500 855.740 ;
        RECT 1015.780 806.860 1016.040 807.120 ;
        RECT 1015.780 724.240 1016.040 724.500 ;
        RECT 1016.240 669.840 1016.500 670.100 ;
        RECT 1015.320 662.360 1015.580 662.620 ;
        RECT 1015.320 620.540 1015.580 620.800 ;
        RECT 1016.240 572.600 1016.500 572.860 ;
        RECT 1015.320 403.280 1015.580 403.540 ;
        RECT 1015.320 355.340 1015.580 355.600 ;
        RECT 1015.320 330.860 1015.580 331.120 ;
        RECT 1016.700 330.860 1016.960 331.120 ;
        RECT 1016.700 324.060 1016.960 324.320 ;
        RECT 1015.320 276.120 1015.580 276.380 ;
        RECT 1015.780 144.540 1016.040 144.800 ;
        RECT 1016.240 144.540 1016.500 144.800 ;
        RECT 490.460 40.840 490.720 41.100 ;
        RECT 1015.780 40.840 1016.040 41.100 ;
      LAYER met2 ;
        RECT 1017.990 1100.580 1018.270 1104.000 ;
        RECT 1017.990 1100.000 1018.280 1100.580 ;
        RECT 1018.140 1062.830 1018.280 1100.000 ;
        RECT 1017.160 1062.510 1017.420 1062.830 ;
        RECT 1018.080 1062.510 1018.340 1062.830 ;
        RECT 1017.220 1014.290 1017.360 1062.510 ;
        RECT 1016.760 1014.150 1017.360 1014.290 ;
        RECT 1016.760 966.270 1016.900 1014.150 ;
        RECT 1016.240 965.950 1016.500 966.270 ;
        RECT 1016.700 965.950 1016.960 966.270 ;
        RECT 1016.300 855.770 1016.440 965.950 ;
        RECT 1015.780 855.450 1016.040 855.770 ;
        RECT 1016.240 855.450 1016.500 855.770 ;
        RECT 1015.840 807.150 1015.980 855.450 ;
        RECT 1015.780 806.830 1016.040 807.150 ;
        RECT 1015.780 724.210 1016.040 724.530 ;
        RECT 1015.840 717.810 1015.980 724.210 ;
        RECT 1015.840 717.670 1016.440 717.810 ;
        RECT 1016.300 670.130 1016.440 717.670 ;
        RECT 1016.240 669.810 1016.500 670.130 ;
        RECT 1015.320 662.330 1015.580 662.650 ;
        RECT 1015.380 620.830 1015.520 662.330 ;
        RECT 1015.320 620.510 1015.580 620.830 ;
        RECT 1016.240 572.570 1016.500 572.890 ;
        RECT 1016.300 483.210 1016.440 572.570 ;
        RECT 1015.840 483.070 1016.440 483.210 ;
        RECT 1015.840 435.725 1015.980 483.070 ;
        RECT 1015.770 435.355 1016.050 435.725 ;
        RECT 1015.310 434.675 1015.590 435.045 ;
        RECT 1015.380 403.570 1015.520 434.675 ;
        RECT 1015.320 403.250 1015.580 403.570 ;
        RECT 1015.320 355.310 1015.580 355.630 ;
        RECT 1015.380 331.150 1015.520 355.310 ;
        RECT 1015.320 330.830 1015.580 331.150 ;
        RECT 1016.700 330.830 1016.960 331.150 ;
        RECT 1016.760 324.350 1016.900 330.830 ;
        RECT 1016.700 324.030 1016.960 324.350 ;
        RECT 1015.320 276.090 1015.580 276.410 ;
        RECT 1015.380 193.530 1015.520 276.090 ;
        RECT 1015.380 193.390 1015.980 193.530 ;
        RECT 1015.840 144.830 1015.980 193.390 ;
        RECT 1015.780 144.510 1016.040 144.830 ;
        RECT 1016.240 144.510 1016.500 144.830 ;
        RECT 1016.300 110.060 1016.440 144.510 ;
        RECT 1015.840 109.920 1016.440 110.060 ;
        RECT 1015.840 41.130 1015.980 109.920 ;
        RECT 490.460 40.810 490.720 41.130 ;
        RECT 1015.780 40.810 1016.040 41.130 ;
        RECT 490.520 2.000 490.660 40.810 ;
        RECT 490.310 -4.000 490.870 2.000 ;
      LAYER via2 ;
        RECT 1015.770 435.400 1016.050 435.680 ;
        RECT 1015.310 434.720 1015.590 435.000 ;
      LAYER met3 ;
        RECT 1015.745 435.690 1016.075 435.705 ;
        RECT 1015.070 435.390 1016.075 435.690 ;
        RECT 1015.070 435.025 1015.370 435.390 ;
        RECT 1015.745 435.375 1016.075 435.390 ;
        RECT 1015.070 434.710 1015.615 435.025 ;
        RECT 1015.285 434.695 1015.615 434.710 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 507.910 41.380 508.230 41.440 ;
        RECT 1022.650 41.380 1022.970 41.440 ;
        RECT 507.910 41.240 1022.970 41.380 ;
        RECT 507.910 41.180 508.230 41.240 ;
        RECT 1022.650 41.180 1022.970 41.240 ;
      LAYER via ;
        RECT 507.940 41.180 508.200 41.440 ;
        RECT 1022.680 41.180 1022.940 41.440 ;
      LAYER met2 ;
        RECT 1024.430 1100.650 1024.710 1104.000 ;
        RECT 1022.740 1100.510 1024.710 1100.650 ;
        RECT 1022.740 41.470 1022.880 1100.510 ;
        RECT 1024.430 1100.000 1024.710 1100.510 ;
        RECT 507.940 41.150 508.200 41.470 ;
        RECT 1022.680 41.150 1022.940 41.470 ;
        RECT 508.000 2.000 508.140 41.150 ;
        RECT 507.790 -4.000 508.350 2.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 525.850 37.640 526.170 37.700 ;
        RECT 1029.090 37.640 1029.410 37.700 ;
        RECT 525.850 37.500 1029.410 37.640 ;
        RECT 525.850 37.440 526.170 37.500 ;
        RECT 1029.090 37.440 1029.410 37.500 ;
      LAYER via ;
        RECT 525.880 37.440 526.140 37.700 ;
        RECT 1029.120 37.440 1029.380 37.700 ;
      LAYER met2 ;
        RECT 1030.410 1100.650 1030.690 1104.000 ;
        RECT 1029.180 1100.510 1030.690 1100.650 ;
        RECT 1029.180 37.730 1029.320 1100.510 ;
        RECT 1030.410 1100.000 1030.690 1100.510 ;
        RECT 525.880 37.410 526.140 37.730 ;
        RECT 1029.120 37.410 1029.380 37.730 ;
        RECT 525.940 2.000 526.080 37.410 ;
        RECT 525.730 -4.000 526.290 2.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 543.790 37.300 544.110 37.360 ;
        RECT 1035.990 37.300 1036.310 37.360 ;
        RECT 543.790 37.160 1036.310 37.300 ;
        RECT 543.790 37.100 544.110 37.160 ;
        RECT 1035.990 37.100 1036.310 37.160 ;
      LAYER via ;
        RECT 543.820 37.100 544.080 37.360 ;
        RECT 1036.020 37.100 1036.280 37.360 ;
      LAYER met2 ;
        RECT 1036.390 1100.650 1036.670 1104.000 ;
        RECT 1036.080 1100.510 1036.670 1100.650 ;
        RECT 1036.080 37.390 1036.220 1100.510 ;
        RECT 1036.390 1100.000 1036.670 1100.510 ;
        RECT 543.820 37.070 544.080 37.390 ;
        RECT 1036.020 37.070 1036.280 37.390 ;
        RECT 543.880 2.000 544.020 37.070 ;
        RECT 543.670 -4.000 544.230 2.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 561.730 36.960 562.050 37.020 ;
        RECT 1042.890 36.960 1043.210 37.020 ;
        RECT 561.730 36.820 1043.210 36.960 ;
        RECT 561.730 36.760 562.050 36.820 ;
        RECT 1042.890 36.760 1043.210 36.820 ;
      LAYER via ;
        RECT 561.760 36.760 562.020 37.020 ;
        RECT 1042.920 36.760 1043.180 37.020 ;
      LAYER met2 ;
        RECT 1042.830 1100.580 1043.110 1104.000 ;
        RECT 1042.830 1100.000 1043.120 1100.580 ;
        RECT 1042.980 37.050 1043.120 1100.000 ;
        RECT 561.760 36.730 562.020 37.050 ;
        RECT 1042.920 36.730 1043.180 37.050 ;
        RECT 561.820 2.000 561.960 36.730 ;
        RECT 561.610 -4.000 562.170 2.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 579.670 36.620 579.990 36.680 ;
        RECT 1048.870 36.620 1049.190 36.680 ;
        RECT 579.670 36.480 1049.190 36.620 ;
        RECT 579.670 36.420 579.990 36.480 ;
        RECT 1048.870 36.420 1049.190 36.480 ;
      LAYER via ;
        RECT 579.700 36.420 579.960 36.680 ;
        RECT 1048.900 36.420 1049.160 36.680 ;
      LAYER met2 ;
        RECT 1048.810 1100.580 1049.090 1104.000 ;
        RECT 1048.810 1100.000 1049.100 1100.580 ;
        RECT 1048.960 36.710 1049.100 1100.000 ;
        RECT 579.700 36.390 579.960 36.710 ;
        RECT 1048.900 36.390 1049.160 36.710 ;
        RECT 579.760 2.000 579.900 36.390 ;
        RECT 579.550 -4.000 580.110 2.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 86.550 25.400 86.870 25.460 ;
        RECT 877.750 25.400 878.070 25.460 ;
        RECT 86.550 25.260 878.070 25.400 ;
        RECT 86.550 25.200 86.870 25.260 ;
        RECT 877.750 25.200 878.070 25.260 ;
      LAYER via ;
        RECT 86.580 25.200 86.840 25.460 ;
        RECT 877.780 25.200 878.040 25.460 ;
      LAYER met2 ;
        RECT 879.530 1100.650 879.810 1104.000 ;
        RECT 877.840 1100.510 879.810 1100.650 ;
        RECT 877.840 25.490 877.980 1100.510 ;
        RECT 879.530 1100.000 879.810 1100.510 ;
        RECT 86.580 25.170 86.840 25.490 ;
        RECT 877.780 25.170 878.040 25.490 ;
        RECT 86.640 12.650 86.780 25.170 ;
        RECT 86.180 12.510 86.780 12.650 ;
        RECT 86.180 2.000 86.320 12.510 ;
        RECT 85.970 -4.000 86.530 2.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1049.330 1076.680 1049.650 1076.740 ;
        RECT 1053.930 1076.680 1054.250 1076.740 ;
        RECT 1049.330 1076.540 1054.250 1076.680 ;
        RECT 1049.330 1076.480 1049.650 1076.540 ;
        RECT 1053.930 1076.480 1054.250 1076.540 ;
        RECT 597.150 36.280 597.470 36.340 ;
        RECT 1049.330 36.280 1049.650 36.340 ;
        RECT 597.150 36.140 1049.650 36.280 ;
        RECT 597.150 36.080 597.470 36.140 ;
        RECT 1049.330 36.080 1049.650 36.140 ;
      LAYER via ;
        RECT 1049.360 1076.480 1049.620 1076.740 ;
        RECT 1053.960 1076.480 1054.220 1076.740 ;
        RECT 597.180 36.080 597.440 36.340 ;
        RECT 1049.360 36.080 1049.620 36.340 ;
      LAYER met2 ;
        RECT 1054.790 1100.650 1055.070 1104.000 ;
        RECT 1054.020 1100.510 1055.070 1100.650 ;
        RECT 1054.020 1076.770 1054.160 1100.510 ;
        RECT 1054.790 1100.000 1055.070 1100.510 ;
        RECT 1049.360 1076.450 1049.620 1076.770 ;
        RECT 1053.960 1076.450 1054.220 1076.770 ;
        RECT 1049.420 36.370 1049.560 1076.450 ;
        RECT 597.180 36.050 597.440 36.370 ;
        RECT 1049.360 36.050 1049.620 36.370 ;
        RECT 597.240 2.000 597.380 36.050 ;
        RECT 597.030 -4.000 597.590 2.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 615.090 35.940 615.410 36.000 ;
        RECT 1056.690 35.940 1057.010 36.000 ;
        RECT 615.090 35.800 1057.010 35.940 ;
        RECT 615.090 35.740 615.410 35.800 ;
        RECT 1056.690 35.740 1057.010 35.800 ;
      LAYER via ;
        RECT 615.120 35.740 615.380 36.000 ;
        RECT 1056.720 35.740 1056.980 36.000 ;
      LAYER met2 ;
        RECT 1060.770 1100.650 1061.050 1104.000 ;
        RECT 1059.540 1100.510 1061.050 1100.650 ;
        RECT 1059.540 1088.410 1059.680 1100.510 ;
        RECT 1060.770 1100.000 1061.050 1100.510 ;
        RECT 1058.620 1088.270 1059.680 1088.410 ;
        RECT 1058.620 1072.770 1058.760 1088.270 ;
        RECT 1056.780 1072.630 1058.760 1072.770 ;
        RECT 1056.780 36.030 1056.920 1072.630 ;
        RECT 615.120 35.710 615.380 36.030 ;
        RECT 1056.720 35.710 1056.980 36.030 ;
        RECT 615.180 2.000 615.320 35.710 ;
        RECT 614.970 -4.000 615.530 2.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 887.350 1100.650 887.630 1104.000 ;
        RECT 886.120 1100.510 887.630 1100.650 ;
        RECT 886.120 1052.200 886.260 1100.510 ;
        RECT 887.350 1100.000 887.630 1100.510 ;
        RECT 884.280 1052.060 886.260 1052.200 ;
        RECT 884.280 31.125 884.420 1052.060 ;
        RECT 109.570 30.755 109.850 31.125 ;
        RECT 884.210 30.755 884.490 31.125 ;
        RECT 109.640 2.000 109.780 30.755 ;
        RECT 109.430 -4.000 109.990 2.000 ;
      LAYER via2 ;
        RECT 109.570 30.800 109.850 31.080 ;
        RECT 884.210 30.800 884.490 31.080 ;
      LAYER met3 ;
        RECT 109.545 31.090 109.875 31.105 ;
        RECT 884.185 31.090 884.515 31.105 ;
        RECT 109.545 30.790 884.515 31.090 ;
        RECT 109.545 30.775 109.875 30.790 ;
        RECT 884.185 30.775 884.515 30.790 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 890.705 697.425 890.875 745.195 ;
        RECT 890.705 648.805 890.875 696.915 ;
        RECT 891.625 552.245 891.795 600.355 ;
        RECT 890.245 455.345 890.415 475.575 ;
        RECT 890.705 317.645 890.875 406.895 ;
        RECT 890.705 83.045 890.875 131.155 ;
      LAYER mcon ;
        RECT 890.705 745.025 890.875 745.195 ;
        RECT 890.705 696.745 890.875 696.915 ;
        RECT 891.625 600.185 891.795 600.355 ;
        RECT 890.245 475.405 890.415 475.575 ;
        RECT 890.705 406.725 890.875 406.895 ;
        RECT 890.705 130.985 890.875 131.155 ;
      LAYER met1 ;
        RECT 894.310 1062.740 894.630 1062.800 ;
        RECT 895.690 1062.740 896.010 1062.800 ;
        RECT 894.310 1062.600 896.010 1062.740 ;
        RECT 894.310 1062.540 894.630 1062.600 ;
        RECT 895.690 1062.540 896.010 1062.600 ;
        RECT 894.310 938.980 894.630 939.040 ;
        RECT 891.180 938.840 894.630 938.980 ;
        RECT 891.180 938.700 891.320 938.840 ;
        RECT 894.310 938.780 894.630 938.840 ;
        RECT 891.090 938.440 891.410 938.700 ;
        RECT 891.090 932.180 891.410 932.240 ;
        RECT 890.720 932.040 891.410 932.180 ;
        RECT 890.720 931.560 890.860 932.040 ;
        RECT 891.090 931.980 891.410 932.040 ;
        RECT 890.630 931.300 890.950 931.560 ;
        RECT 890.170 793.460 890.490 793.520 ;
        RECT 890.630 793.460 890.950 793.520 ;
        RECT 890.170 793.320 890.950 793.460 ;
        RECT 890.170 793.260 890.490 793.320 ;
        RECT 890.630 793.260 890.950 793.320 ;
        RECT 890.630 745.180 890.950 745.240 ;
        RECT 890.435 745.040 890.950 745.180 ;
        RECT 890.630 744.980 890.950 745.040 ;
        RECT 890.630 697.580 890.950 697.640 ;
        RECT 890.435 697.440 890.950 697.580 ;
        RECT 890.630 697.380 890.950 697.440 ;
        RECT 890.630 696.900 890.950 696.960 ;
        RECT 890.435 696.760 890.950 696.900 ;
        RECT 890.630 696.700 890.950 696.760 ;
        RECT 890.645 648.960 890.935 649.005 ;
        RECT 892.010 648.960 892.330 649.020 ;
        RECT 890.645 648.820 892.330 648.960 ;
        RECT 890.645 648.775 890.935 648.820 ;
        RECT 892.010 648.760 892.330 648.820 ;
        RECT 891.550 600.340 891.870 600.400 ;
        RECT 891.355 600.200 891.870 600.340 ;
        RECT 891.550 600.140 891.870 600.200 ;
        RECT 891.565 552.400 891.855 552.445 ;
        RECT 892.470 552.400 892.790 552.460 ;
        RECT 891.565 552.260 892.790 552.400 ;
        RECT 891.565 552.215 891.855 552.260 ;
        RECT 892.470 552.200 892.790 552.260 ;
        RECT 890.630 534.720 890.950 534.780 ;
        RECT 892.470 534.720 892.790 534.780 ;
        RECT 890.630 534.580 892.790 534.720 ;
        RECT 890.630 534.520 890.950 534.580 ;
        RECT 892.470 534.520 892.790 534.580 ;
        RECT 889.710 510.240 890.030 510.300 ;
        RECT 890.630 510.240 890.950 510.300 ;
        RECT 889.710 510.100 890.950 510.240 ;
        RECT 889.710 510.040 890.030 510.100 ;
        RECT 890.630 510.040 890.950 510.100 ;
        RECT 890.170 475.560 890.490 475.620 ;
        RECT 890.170 475.420 890.685 475.560 ;
        RECT 890.170 475.360 890.490 475.420 ;
        RECT 890.185 455.500 890.475 455.545 ;
        RECT 890.630 455.500 890.950 455.560 ;
        RECT 890.185 455.360 890.950 455.500 ;
        RECT 890.185 455.315 890.475 455.360 ;
        RECT 890.630 455.300 890.950 455.360 ;
        RECT 890.630 406.880 890.950 406.940 ;
        RECT 890.435 406.740 890.950 406.880 ;
        RECT 890.630 406.680 890.950 406.740 ;
        RECT 890.645 317.800 890.935 317.845 ;
        RECT 891.550 317.800 891.870 317.860 ;
        RECT 890.645 317.660 891.870 317.800 ;
        RECT 890.645 317.615 890.935 317.660 ;
        RECT 891.550 317.600 891.870 317.660 ;
        RECT 890.170 269.180 890.490 269.240 ;
        RECT 890.630 269.180 890.950 269.240 ;
        RECT 890.170 269.040 890.950 269.180 ;
        RECT 890.170 268.980 890.490 269.040 ;
        RECT 890.630 268.980 890.950 269.040 ;
        RECT 890.630 179.760 890.950 179.820 ;
        RECT 891.090 179.760 891.410 179.820 ;
        RECT 890.630 179.620 891.410 179.760 ;
        RECT 890.630 179.560 890.950 179.620 ;
        RECT 891.090 179.560 891.410 179.620 ;
        RECT 891.090 159.020 891.410 159.080 ;
        RECT 890.720 158.880 891.410 159.020 ;
        RECT 890.720 158.740 890.860 158.880 ;
        RECT 891.090 158.820 891.410 158.880 ;
        RECT 890.630 158.480 890.950 158.740 ;
        RECT 890.630 131.140 890.950 131.200 ;
        RECT 890.435 131.000 890.950 131.140 ;
        RECT 890.630 130.940 890.950 131.000 ;
        RECT 890.630 83.200 890.950 83.260 ;
        RECT 890.435 83.060 890.950 83.200 ;
        RECT 890.630 83.000 890.950 83.060 ;
        RECT 133.470 31.520 133.790 31.580 ;
        RECT 890.630 31.520 890.950 31.580 ;
        RECT 133.470 31.380 890.950 31.520 ;
        RECT 133.470 31.320 133.790 31.380 ;
        RECT 890.630 31.320 890.950 31.380 ;
      LAYER via ;
        RECT 894.340 1062.540 894.600 1062.800 ;
        RECT 895.720 1062.540 895.980 1062.800 ;
        RECT 894.340 938.780 894.600 939.040 ;
        RECT 891.120 938.440 891.380 938.700 ;
        RECT 891.120 931.980 891.380 932.240 ;
        RECT 890.660 931.300 890.920 931.560 ;
        RECT 890.200 793.260 890.460 793.520 ;
        RECT 890.660 793.260 890.920 793.520 ;
        RECT 890.660 744.980 890.920 745.240 ;
        RECT 890.660 697.380 890.920 697.640 ;
        RECT 890.660 696.700 890.920 696.960 ;
        RECT 892.040 648.760 892.300 649.020 ;
        RECT 891.580 600.140 891.840 600.400 ;
        RECT 892.500 552.200 892.760 552.460 ;
        RECT 890.660 534.520 890.920 534.780 ;
        RECT 892.500 534.520 892.760 534.780 ;
        RECT 889.740 510.040 890.000 510.300 ;
        RECT 890.660 510.040 890.920 510.300 ;
        RECT 890.200 475.360 890.460 475.620 ;
        RECT 890.660 455.300 890.920 455.560 ;
        RECT 890.660 406.680 890.920 406.940 ;
        RECT 891.580 317.600 891.840 317.860 ;
        RECT 890.200 268.980 890.460 269.240 ;
        RECT 890.660 268.980 890.920 269.240 ;
        RECT 890.660 179.560 890.920 179.820 ;
        RECT 891.120 179.560 891.380 179.820 ;
        RECT 891.120 158.820 891.380 159.080 ;
        RECT 890.660 158.480 890.920 158.740 ;
        RECT 890.660 130.940 890.920 131.200 ;
        RECT 890.660 83.000 890.920 83.260 ;
        RECT 133.500 31.320 133.760 31.580 ;
        RECT 890.660 31.320 890.920 31.580 ;
      LAYER met2 ;
        RECT 895.630 1100.580 895.910 1104.000 ;
        RECT 895.630 1100.000 895.920 1100.580 ;
        RECT 895.780 1062.830 895.920 1100.000 ;
        RECT 894.340 1062.510 894.600 1062.830 ;
        RECT 895.720 1062.510 895.980 1062.830 ;
        RECT 894.400 939.070 894.540 1062.510 ;
        RECT 894.340 938.750 894.600 939.070 ;
        RECT 891.120 938.410 891.380 938.730 ;
        RECT 891.180 932.270 891.320 938.410 ;
        RECT 891.120 931.950 891.380 932.270 ;
        RECT 890.660 931.270 890.920 931.590 ;
        RECT 890.720 896.650 890.860 931.270 ;
        RECT 890.720 896.510 891.320 896.650 ;
        RECT 891.180 883.730 891.320 896.510 ;
        RECT 890.260 883.590 891.320 883.730 ;
        RECT 890.260 793.550 890.400 883.590 ;
        RECT 890.200 793.230 890.460 793.550 ;
        RECT 890.660 793.230 890.920 793.550 ;
        RECT 890.720 745.270 890.860 793.230 ;
        RECT 890.660 744.950 890.920 745.270 ;
        RECT 890.660 697.350 890.920 697.670 ;
        RECT 890.720 696.990 890.860 697.350 ;
        RECT 890.660 696.670 890.920 696.990 ;
        RECT 892.040 648.730 892.300 649.050 ;
        RECT 892.100 613.770 892.240 648.730 ;
        RECT 891.640 613.630 892.240 613.770 ;
        RECT 891.640 600.430 891.780 613.630 ;
        RECT 891.580 600.110 891.840 600.430 ;
        RECT 892.500 552.170 892.760 552.490 ;
        RECT 892.560 534.810 892.700 552.170 ;
        RECT 890.660 534.490 890.920 534.810 ;
        RECT 892.500 534.490 892.760 534.810 ;
        RECT 890.720 510.330 890.860 534.490 ;
        RECT 889.740 510.010 890.000 510.330 ;
        RECT 890.660 510.010 890.920 510.330 ;
        RECT 889.800 475.730 889.940 510.010 ;
        RECT 889.800 475.650 890.400 475.730 ;
        RECT 889.800 475.590 890.460 475.650 ;
        RECT 890.200 475.330 890.460 475.590 ;
        RECT 890.660 455.270 890.920 455.590 ;
        RECT 890.720 406.970 890.860 455.270 ;
        RECT 890.660 406.650 890.920 406.970 ;
        RECT 891.580 317.570 891.840 317.890 ;
        RECT 891.640 317.405 891.780 317.570 ;
        RECT 890.190 317.035 890.470 317.405 ;
        RECT 891.570 317.035 891.850 317.405 ;
        RECT 890.260 269.270 890.400 317.035 ;
        RECT 890.200 268.950 890.460 269.270 ;
        RECT 890.660 268.950 890.920 269.270 ;
        RECT 890.720 179.850 890.860 268.950 ;
        RECT 890.660 179.530 890.920 179.850 ;
        RECT 891.120 179.530 891.380 179.850 ;
        RECT 891.180 159.110 891.320 179.530 ;
        RECT 891.120 158.790 891.380 159.110 ;
        RECT 890.660 158.450 890.920 158.770 ;
        RECT 890.720 131.230 890.860 158.450 ;
        RECT 890.660 130.910 890.920 131.230 ;
        RECT 890.660 82.970 890.920 83.290 ;
        RECT 890.720 31.610 890.860 82.970 ;
        RECT 133.500 31.290 133.760 31.610 ;
        RECT 890.660 31.290 890.920 31.610 ;
        RECT 133.560 2.000 133.700 31.290 ;
        RECT 133.350 -4.000 133.910 2.000 ;
      LAYER via2 ;
        RECT 890.190 317.080 890.470 317.360 ;
        RECT 891.570 317.080 891.850 317.360 ;
      LAYER met3 ;
        RECT 890.165 317.370 890.495 317.385 ;
        RECT 891.545 317.370 891.875 317.385 ;
        RECT 890.165 317.070 891.875 317.370 ;
        RECT 890.165 317.055 890.495 317.070 ;
        RECT 891.545 317.055 891.875 317.070 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 897.530 1052.200 897.850 1052.260 ;
        RECT 900.290 1052.200 900.610 1052.260 ;
        RECT 897.530 1052.060 900.610 1052.200 ;
        RECT 897.530 1052.000 897.850 1052.060 ;
        RECT 900.290 1052.000 900.610 1052.060 ;
        RECT 151.410 31.860 151.730 31.920 ;
        RECT 897.530 31.860 897.850 31.920 ;
        RECT 151.410 31.720 897.850 31.860 ;
        RECT 151.410 31.660 151.730 31.720 ;
        RECT 897.530 31.660 897.850 31.720 ;
      LAYER via ;
        RECT 897.560 1052.000 897.820 1052.260 ;
        RECT 900.320 1052.000 900.580 1052.260 ;
        RECT 151.440 31.660 151.700 31.920 ;
        RECT 897.560 31.660 897.820 31.920 ;
      LAYER met2 ;
        RECT 901.610 1100.650 901.890 1104.000 ;
        RECT 900.380 1100.510 901.890 1100.650 ;
        RECT 900.380 1052.290 900.520 1100.510 ;
        RECT 901.610 1100.000 901.890 1100.510 ;
        RECT 897.560 1051.970 897.820 1052.290 ;
        RECT 900.320 1051.970 900.580 1052.290 ;
        RECT 897.620 31.950 897.760 1051.970 ;
        RECT 151.440 31.630 151.700 31.950 ;
        RECT 897.560 31.630 897.820 31.950 ;
        RECT 151.500 2.000 151.640 31.630 ;
        RECT 151.290 -4.000 151.850 2.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 904.430 1052.200 904.750 1052.260 ;
        RECT 906.270 1052.200 906.590 1052.260 ;
        RECT 904.430 1052.060 906.590 1052.200 ;
        RECT 904.430 1052.000 904.750 1052.060 ;
        RECT 906.270 1052.000 906.590 1052.060 ;
        RECT 169.350 32.200 169.670 32.260 ;
        RECT 904.430 32.200 904.750 32.260 ;
        RECT 169.350 32.060 904.750 32.200 ;
        RECT 169.350 32.000 169.670 32.060 ;
        RECT 904.430 32.000 904.750 32.060 ;
      LAYER via ;
        RECT 904.460 1052.000 904.720 1052.260 ;
        RECT 906.300 1052.000 906.560 1052.260 ;
        RECT 169.380 32.000 169.640 32.260 ;
        RECT 904.460 32.000 904.720 32.260 ;
      LAYER met2 ;
        RECT 908.050 1100.650 908.330 1104.000 ;
        RECT 906.360 1100.510 908.330 1100.650 ;
        RECT 906.360 1052.290 906.500 1100.510 ;
        RECT 908.050 1100.000 908.330 1100.510 ;
        RECT 904.460 1051.970 904.720 1052.290 ;
        RECT 906.300 1051.970 906.560 1052.290 ;
        RECT 904.520 32.290 904.660 1051.970 ;
        RECT 169.380 31.970 169.640 32.290 ;
        RECT 904.460 31.970 904.720 32.290 ;
        RECT 169.440 2.000 169.580 31.970 ;
        RECT 169.230 -4.000 169.790 2.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 910.945 910.945 911.115 931.855 ;
        RECT 910.945 882.725 911.115 910.095 ;
        RECT 910.945 807.245 911.115 855.355 ;
        RECT 910.945 783.445 911.115 806.735 ;
        RECT 910.945 620.925 911.115 710.515 ;
        RECT 910.945 589.985 911.115 613.955 ;
        RECT 910.945 496.485 911.115 523.855 ;
        RECT 910.945 421.005 911.115 469.115 ;
        RECT 910.945 138.125 911.115 207.315 ;
      LAYER mcon ;
        RECT 910.945 931.685 911.115 931.855 ;
        RECT 910.945 909.925 911.115 910.095 ;
        RECT 910.945 855.185 911.115 855.355 ;
        RECT 910.945 806.565 911.115 806.735 ;
        RECT 910.945 710.345 911.115 710.515 ;
        RECT 910.945 613.785 911.115 613.955 ;
        RECT 910.945 523.685 911.115 523.855 ;
        RECT 910.945 468.945 911.115 469.115 ;
        RECT 910.945 207.145 911.115 207.315 ;
      LAYER met1 ;
        RECT 911.330 1028.400 911.650 1028.460 ;
        RECT 912.710 1028.400 913.030 1028.460 ;
        RECT 911.330 1028.260 913.030 1028.400 ;
        RECT 911.330 1028.200 911.650 1028.260 ;
        RECT 912.710 1028.200 913.030 1028.260 ;
        RECT 910.870 931.840 911.190 931.900 ;
        RECT 910.870 931.700 911.385 931.840 ;
        RECT 910.870 931.640 911.190 931.700 ;
        RECT 910.870 911.100 911.190 911.160 ;
        RECT 910.870 910.960 911.385 911.100 ;
        RECT 910.870 910.900 911.190 910.960 ;
        RECT 910.870 910.080 911.190 910.140 ;
        RECT 910.870 909.940 911.385 910.080 ;
        RECT 910.870 909.880 911.190 909.940 ;
        RECT 910.885 882.880 911.175 882.925 ;
        RECT 911.330 882.880 911.650 882.940 ;
        RECT 910.885 882.740 911.650 882.880 ;
        RECT 910.885 882.695 911.175 882.740 ;
        RECT 911.330 882.680 911.650 882.740 ;
        RECT 910.885 855.340 911.175 855.385 ;
        RECT 911.330 855.340 911.650 855.400 ;
        RECT 910.885 855.200 911.650 855.340 ;
        RECT 910.885 855.155 911.175 855.200 ;
        RECT 911.330 855.140 911.650 855.200 ;
        RECT 910.870 807.400 911.190 807.460 ;
        RECT 910.675 807.260 911.190 807.400 ;
        RECT 910.870 807.200 911.190 807.260 ;
        RECT 910.870 806.720 911.190 806.780 ;
        RECT 910.675 806.580 911.190 806.720 ;
        RECT 910.870 806.520 911.190 806.580 ;
        RECT 910.870 783.600 911.190 783.660 ;
        RECT 910.675 783.460 911.190 783.600 ;
        RECT 910.870 783.400 911.190 783.460 ;
        RECT 910.870 710.500 911.190 710.560 ;
        RECT 910.675 710.360 911.190 710.500 ;
        RECT 910.870 710.300 911.190 710.360 ;
        RECT 910.870 621.080 911.190 621.140 ;
        RECT 910.870 620.940 911.385 621.080 ;
        RECT 910.870 620.880 911.190 620.940 ;
        RECT 910.870 613.940 911.190 614.000 ;
        RECT 910.675 613.800 911.190 613.940 ;
        RECT 910.870 613.740 911.190 613.800 ;
        RECT 910.870 590.140 911.190 590.200 ;
        RECT 910.675 590.000 911.190 590.140 ;
        RECT 910.870 589.940 911.190 590.000 ;
        RECT 910.870 545.060 911.190 545.320 ;
        RECT 910.960 544.640 911.100 545.060 ;
        RECT 910.870 544.380 911.190 544.640 ;
        RECT 910.870 523.840 911.190 523.900 ;
        RECT 910.870 523.700 911.385 523.840 ;
        RECT 910.870 523.640 911.190 523.700 ;
        RECT 910.885 496.640 911.175 496.685 ;
        RECT 911.330 496.640 911.650 496.700 ;
        RECT 910.885 496.500 911.650 496.640 ;
        RECT 910.885 496.455 911.175 496.500 ;
        RECT 911.330 496.440 911.650 496.500 ;
        RECT 910.885 469.100 911.175 469.145 ;
        RECT 911.330 469.100 911.650 469.160 ;
        RECT 910.885 468.960 911.650 469.100 ;
        RECT 910.885 468.915 911.175 468.960 ;
        RECT 911.330 468.900 911.650 468.960 ;
        RECT 910.870 421.160 911.190 421.220 ;
        RECT 910.675 421.020 911.190 421.160 ;
        RECT 910.870 420.960 911.190 421.020 ;
        RECT 910.870 207.300 911.190 207.360 ;
        RECT 910.675 207.160 911.190 207.300 ;
        RECT 910.870 207.100 911.190 207.160 ;
        RECT 910.870 138.280 911.190 138.340 ;
        RECT 910.870 138.140 911.385 138.280 ;
        RECT 910.870 138.080 911.190 138.140 ;
        RECT 910.870 131.140 911.190 131.200 ;
        RECT 912.250 131.140 912.570 131.200 ;
        RECT 910.870 131.000 912.570 131.140 ;
        RECT 910.870 130.940 911.190 131.000 ;
        RECT 912.250 130.940 912.570 131.000 ;
        RECT 910.870 41.720 911.190 41.780 ;
        RECT 912.250 41.720 912.570 41.780 ;
        RECT 910.870 41.580 912.570 41.720 ;
        RECT 910.870 41.520 911.190 41.580 ;
        RECT 912.250 41.520 912.570 41.580 ;
        RECT 186.830 32.540 187.150 32.600 ;
        RECT 911.330 32.540 911.650 32.600 ;
        RECT 186.830 32.400 911.650 32.540 ;
        RECT 186.830 32.340 187.150 32.400 ;
        RECT 911.330 32.340 911.650 32.400 ;
      LAYER via ;
        RECT 911.360 1028.200 911.620 1028.460 ;
        RECT 912.740 1028.200 913.000 1028.460 ;
        RECT 910.900 931.640 911.160 931.900 ;
        RECT 910.900 910.900 911.160 911.160 ;
        RECT 910.900 909.880 911.160 910.140 ;
        RECT 911.360 882.680 911.620 882.940 ;
        RECT 911.360 855.140 911.620 855.400 ;
        RECT 910.900 807.200 911.160 807.460 ;
        RECT 910.900 806.520 911.160 806.780 ;
        RECT 910.900 783.400 911.160 783.660 ;
        RECT 910.900 710.300 911.160 710.560 ;
        RECT 910.900 620.880 911.160 621.140 ;
        RECT 910.900 613.740 911.160 614.000 ;
        RECT 910.900 589.940 911.160 590.200 ;
        RECT 910.900 545.060 911.160 545.320 ;
        RECT 910.900 544.380 911.160 544.640 ;
        RECT 910.900 523.640 911.160 523.900 ;
        RECT 911.360 496.440 911.620 496.700 ;
        RECT 911.360 468.900 911.620 469.160 ;
        RECT 910.900 420.960 911.160 421.220 ;
        RECT 910.900 207.100 911.160 207.360 ;
        RECT 910.900 138.080 911.160 138.340 ;
        RECT 910.900 130.940 911.160 131.200 ;
        RECT 912.280 130.940 912.540 131.200 ;
        RECT 910.900 41.520 911.160 41.780 ;
        RECT 912.280 41.520 912.540 41.780 ;
        RECT 186.860 32.340 187.120 32.600 ;
        RECT 911.360 32.340 911.620 32.600 ;
      LAYER met2 ;
        RECT 914.030 1100.650 914.310 1104.000 ;
        RECT 912.800 1100.510 914.310 1100.650 ;
        RECT 912.800 1028.490 912.940 1100.510 ;
        RECT 914.030 1100.000 914.310 1100.510 ;
        RECT 911.360 1028.170 911.620 1028.490 ;
        RECT 912.740 1028.170 913.000 1028.490 ;
        RECT 911.420 979.610 911.560 1028.170 ;
        RECT 910.960 979.470 911.560 979.610 ;
        RECT 910.960 931.930 911.100 979.470 ;
        RECT 910.900 931.610 911.160 931.930 ;
        RECT 910.900 910.870 911.160 911.190 ;
        RECT 910.960 910.170 911.100 910.870 ;
        RECT 910.900 909.850 911.160 910.170 ;
        RECT 911.360 882.650 911.620 882.970 ;
        RECT 911.420 855.430 911.560 882.650 ;
        RECT 911.360 855.110 911.620 855.430 ;
        RECT 910.900 807.170 911.160 807.490 ;
        RECT 910.960 806.810 911.100 807.170 ;
        RECT 910.900 806.490 911.160 806.810 ;
        RECT 910.900 783.370 911.160 783.690 ;
        RECT 910.960 710.590 911.100 783.370 ;
        RECT 910.900 710.270 911.160 710.590 ;
        RECT 910.900 620.850 911.160 621.170 ;
        RECT 910.960 614.030 911.100 620.850 ;
        RECT 910.900 613.710 911.160 614.030 ;
        RECT 910.900 589.910 911.160 590.230 ;
        RECT 910.960 545.350 911.100 589.910 ;
        RECT 910.900 545.030 911.160 545.350 ;
        RECT 910.900 544.350 911.160 544.670 ;
        RECT 910.960 523.930 911.100 544.350 ;
        RECT 910.900 523.610 911.160 523.930 ;
        RECT 911.360 496.410 911.620 496.730 ;
        RECT 911.420 469.190 911.560 496.410 ;
        RECT 911.360 468.870 911.620 469.190 ;
        RECT 910.900 420.930 911.160 421.250 ;
        RECT 910.960 207.390 911.100 420.930 ;
        RECT 910.900 207.070 911.160 207.390 ;
        RECT 910.900 138.050 911.160 138.370 ;
        RECT 910.960 131.230 911.100 138.050 ;
        RECT 910.900 130.910 911.160 131.230 ;
        RECT 912.280 130.910 912.540 131.230 ;
        RECT 912.340 41.810 912.480 130.910 ;
        RECT 910.900 41.490 911.160 41.810 ;
        RECT 912.280 41.490 912.540 41.810 ;
        RECT 910.960 41.210 911.100 41.490 ;
        RECT 910.960 41.070 911.560 41.210 ;
        RECT 911.420 32.630 911.560 41.070 ;
        RECT 186.860 32.310 187.120 32.630 ;
        RECT 911.360 32.310 911.620 32.630 ;
        RECT 186.920 2.000 187.060 32.310 ;
        RECT 186.710 -4.000 187.270 2.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 204.770 32.880 205.090 32.940 ;
        RECT 918.690 32.880 919.010 32.940 ;
        RECT 204.770 32.740 919.010 32.880 ;
        RECT 204.770 32.680 205.090 32.740 ;
        RECT 918.690 32.680 919.010 32.740 ;
      LAYER via ;
        RECT 204.800 32.680 205.060 32.940 ;
        RECT 918.720 32.680 918.980 32.940 ;
      LAYER met2 ;
        RECT 920.010 1100.650 920.290 1104.000 ;
        RECT 918.780 1100.510 920.290 1100.650 ;
        RECT 918.780 32.970 918.920 1100.510 ;
        RECT 920.010 1100.000 920.290 1100.510 ;
        RECT 204.800 32.650 205.060 32.970 ;
        RECT 918.720 32.650 918.980 32.970 ;
        RECT 204.860 2.000 205.000 32.650 ;
        RECT 204.650 -4.000 205.210 2.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 222.710 33.220 223.030 33.280 ;
        RECT 925.590 33.220 925.910 33.280 ;
        RECT 222.710 33.080 925.910 33.220 ;
        RECT 222.710 33.020 223.030 33.080 ;
        RECT 925.590 33.020 925.910 33.080 ;
      LAYER via ;
        RECT 222.740 33.020 223.000 33.280 ;
        RECT 925.620 33.020 925.880 33.280 ;
      LAYER met2 ;
        RECT 926.450 1100.650 926.730 1104.000 ;
        RECT 925.680 1100.510 926.730 1100.650 ;
        RECT 925.680 33.310 925.820 1100.510 ;
        RECT 926.450 1100.000 926.730 1100.510 ;
        RECT 222.740 32.990 223.000 33.310 ;
        RECT 925.620 32.990 925.880 33.310 ;
        RECT 222.800 2.000 222.940 32.990 ;
        RECT 222.590 -4.000 223.150 2.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 20.310 30.840 20.630 30.900 ;
        RECT 856.130 30.840 856.450 30.900 ;
        RECT 20.310 30.700 856.450 30.840 ;
        RECT 20.310 30.640 20.630 30.700 ;
        RECT 856.130 30.640 856.450 30.700 ;
      LAYER via ;
        RECT 20.340 30.640 20.600 30.900 ;
        RECT 856.160 30.640 856.420 30.900 ;
      LAYER met2 ;
        RECT 856.990 1100.650 857.270 1104.000 ;
        RECT 856.220 1100.510 857.270 1100.650 ;
        RECT 856.220 30.930 856.360 1100.510 ;
        RECT 856.990 1100.000 857.270 1100.510 ;
        RECT 20.340 30.610 20.600 30.930 ;
        RECT 856.160 30.610 856.420 30.930 ;
        RECT 20.400 2.000 20.540 30.610 ;
        RECT 20.190 -4.000 20.750 2.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 44.230 31.180 44.550 31.240 ;
        RECT 863.950 31.180 864.270 31.240 ;
        RECT 44.230 31.040 864.270 31.180 ;
        RECT 44.230 30.980 44.550 31.040 ;
        RECT 863.950 30.980 864.270 31.040 ;
      LAYER via ;
        RECT 44.260 30.980 44.520 31.240 ;
        RECT 863.980 30.980 864.240 31.240 ;
      LAYER met2 ;
        RECT 865.270 1100.650 865.550 1104.000 ;
        RECT 864.040 1100.510 865.550 1100.650 ;
        RECT 864.040 31.270 864.180 1100.510 ;
        RECT 865.270 1100.000 865.550 1100.510 ;
        RECT 44.260 30.950 44.520 31.270 ;
        RECT 863.980 30.950 864.240 31.270 ;
        RECT 44.320 2.000 44.460 30.950 ;
        RECT 44.110 -4.000 44.670 2.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 932.030 1052.200 932.350 1052.260 ;
        RECT 932.950 1052.200 933.270 1052.260 ;
        RECT 932.030 1052.060 933.270 1052.200 ;
        RECT 932.030 1052.000 932.350 1052.060 ;
        RECT 932.950 1052.000 933.270 1052.060 ;
        RECT 246.630 33.560 246.950 33.620 ;
        RECT 932.030 33.560 932.350 33.620 ;
        RECT 246.630 33.420 932.350 33.560 ;
        RECT 246.630 33.360 246.950 33.420 ;
        RECT 932.030 33.360 932.350 33.420 ;
      LAYER via ;
        RECT 932.060 1052.000 932.320 1052.260 ;
        RECT 932.980 1052.000 933.240 1052.260 ;
        RECT 246.660 33.360 246.920 33.620 ;
        RECT 932.060 33.360 932.320 33.620 ;
      LAYER met2 ;
        RECT 934.270 1100.650 934.550 1104.000 ;
        RECT 933.040 1100.510 934.550 1100.650 ;
        RECT 933.040 1052.290 933.180 1100.510 ;
        RECT 934.270 1100.000 934.550 1100.510 ;
        RECT 932.060 1051.970 932.320 1052.290 ;
        RECT 932.980 1051.970 933.240 1052.290 ;
        RECT 932.120 33.650 932.260 1051.970 ;
        RECT 246.660 33.330 246.920 33.650 ;
        RECT 932.060 33.330 932.320 33.650 ;
        RECT 246.720 2.000 246.860 33.330 ;
        RECT 246.510 -4.000 247.070 2.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 940.710 1100.650 940.990 1104.000 ;
        RECT 939.480 1100.510 940.990 1100.650 ;
        RECT 939.480 37.925 939.620 1100.510 ;
        RECT 940.710 1100.000 940.990 1100.510 ;
        RECT 264.130 37.555 264.410 37.925 ;
        RECT 939.410 37.555 939.690 37.925 ;
        RECT 264.200 2.000 264.340 37.555 ;
        RECT 263.990 -4.000 264.550 2.000 ;
      LAYER via2 ;
        RECT 264.130 37.600 264.410 37.880 ;
        RECT 939.410 37.600 939.690 37.880 ;
      LAYER met3 ;
        RECT 264.105 37.890 264.435 37.905 ;
        RECT 939.385 37.890 939.715 37.905 ;
        RECT 264.105 37.590 939.715 37.890 ;
        RECT 264.105 37.575 264.435 37.590 ;
        RECT 939.385 37.575 939.715 37.590 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 282.050 37.980 282.370 38.040 ;
        RECT 945.830 37.980 946.150 38.040 ;
        RECT 282.050 37.840 946.150 37.980 ;
        RECT 282.050 37.780 282.370 37.840 ;
        RECT 945.830 37.780 946.150 37.840 ;
      LAYER via ;
        RECT 282.080 37.780 282.340 38.040 ;
        RECT 945.860 37.780 946.120 38.040 ;
      LAYER met2 ;
        RECT 946.690 1100.650 946.970 1104.000 ;
        RECT 945.920 1100.510 946.970 1100.650 ;
        RECT 945.920 38.070 946.060 1100.510 ;
        RECT 946.690 1100.000 946.970 1100.510 ;
        RECT 282.080 37.750 282.340 38.070 ;
        RECT 945.860 37.750 946.120 38.070 ;
        RECT 282.140 2.000 282.280 37.750 ;
        RECT 281.930 -4.000 282.490 2.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 299.990 38.320 300.310 38.380 ;
        RECT 952.730 38.320 953.050 38.380 ;
        RECT 299.990 38.180 953.050 38.320 ;
        RECT 299.990 38.120 300.310 38.180 ;
        RECT 952.730 38.120 953.050 38.180 ;
      LAYER via ;
        RECT 300.020 38.120 300.280 38.380 ;
        RECT 952.760 38.120 953.020 38.380 ;
      LAYER met2 ;
        RECT 952.670 1100.580 952.950 1104.000 ;
        RECT 952.670 1100.000 952.960 1100.580 ;
        RECT 952.820 38.410 952.960 1100.000 ;
        RECT 300.020 38.090 300.280 38.410 ;
        RECT 952.760 38.090 953.020 38.410 ;
        RECT 300.080 2.000 300.220 38.090 ;
        RECT 299.870 -4.000 300.430 2.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 317.930 38.660 318.250 38.720 ;
        RECT 959.630 38.660 959.950 38.720 ;
        RECT 317.930 38.520 959.950 38.660 ;
        RECT 317.930 38.460 318.250 38.520 ;
        RECT 959.630 38.460 959.950 38.520 ;
      LAYER via ;
        RECT 317.960 38.460 318.220 38.720 ;
        RECT 959.660 38.460 959.920 38.720 ;
      LAYER met2 ;
        RECT 959.110 1100.650 959.390 1104.000 ;
        RECT 959.110 1100.510 959.860 1100.650 ;
        RECT 959.110 1100.000 959.390 1100.510 ;
        RECT 959.720 38.750 959.860 1100.510 ;
        RECT 317.960 38.430 318.220 38.750 ;
        RECT 959.660 38.430 959.920 38.750 ;
        RECT 318.020 2.000 318.160 38.430 ;
        RECT 317.810 -4.000 318.370 2.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 960.090 1052.200 960.410 1052.260 ;
        RECT 963.770 1052.200 964.090 1052.260 ;
        RECT 960.090 1052.060 964.090 1052.200 ;
        RECT 960.090 1052.000 960.410 1052.060 ;
        RECT 963.770 1052.000 964.090 1052.060 ;
        RECT 335.870 45.800 336.190 45.860 ;
        RECT 960.090 45.800 960.410 45.860 ;
        RECT 335.870 45.660 960.410 45.800 ;
        RECT 335.870 45.600 336.190 45.660 ;
        RECT 960.090 45.600 960.410 45.660 ;
      LAYER via ;
        RECT 960.120 1052.000 960.380 1052.260 ;
        RECT 963.800 1052.000 964.060 1052.260 ;
        RECT 335.900 45.600 336.160 45.860 ;
        RECT 960.120 45.600 960.380 45.860 ;
      LAYER met2 ;
        RECT 965.090 1100.650 965.370 1104.000 ;
        RECT 963.860 1100.510 965.370 1100.650 ;
        RECT 963.860 1052.290 964.000 1100.510 ;
        RECT 965.090 1100.000 965.370 1100.510 ;
        RECT 960.120 1051.970 960.380 1052.290 ;
        RECT 963.800 1051.970 964.060 1052.290 ;
        RECT 960.180 45.890 960.320 1051.970 ;
        RECT 335.900 45.570 336.160 45.890 ;
        RECT 960.120 45.570 960.380 45.890 ;
        RECT 335.960 2.000 336.100 45.570 ;
        RECT 335.750 -4.000 336.310 2.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 966.530 1052.200 966.850 1052.260 ;
        RECT 969.750 1052.200 970.070 1052.260 ;
        RECT 966.530 1052.060 970.070 1052.200 ;
        RECT 966.530 1052.000 966.850 1052.060 ;
        RECT 969.750 1052.000 970.070 1052.060 ;
        RECT 358.410 51.920 358.730 51.980 ;
        RECT 966.530 51.920 966.850 51.980 ;
        RECT 358.410 51.780 966.850 51.920 ;
        RECT 358.410 51.720 358.730 51.780 ;
        RECT 966.530 51.720 966.850 51.780 ;
        RECT 353.350 16.900 353.670 16.960 ;
        RECT 358.410 16.900 358.730 16.960 ;
        RECT 353.350 16.760 358.730 16.900 ;
        RECT 353.350 16.700 353.670 16.760 ;
        RECT 358.410 16.700 358.730 16.760 ;
      LAYER via ;
        RECT 966.560 1052.000 966.820 1052.260 ;
        RECT 969.780 1052.000 970.040 1052.260 ;
        RECT 358.440 51.720 358.700 51.980 ;
        RECT 966.560 51.720 966.820 51.980 ;
        RECT 353.380 16.700 353.640 16.960 ;
        RECT 358.440 16.700 358.700 16.960 ;
      LAYER met2 ;
        RECT 971.070 1100.650 971.350 1104.000 ;
        RECT 969.840 1100.510 971.350 1100.650 ;
        RECT 969.840 1052.290 969.980 1100.510 ;
        RECT 971.070 1100.000 971.350 1100.510 ;
        RECT 966.560 1051.970 966.820 1052.290 ;
        RECT 969.780 1051.970 970.040 1052.290 ;
        RECT 966.620 52.010 966.760 1051.970 ;
        RECT 358.440 51.690 358.700 52.010 ;
        RECT 966.560 51.690 966.820 52.010 ;
        RECT 358.500 16.990 358.640 51.690 ;
        RECT 353.380 16.670 353.640 16.990 ;
        RECT 358.440 16.670 358.700 16.990 ;
        RECT 353.440 2.000 353.580 16.670 ;
        RECT 353.230 -4.000 353.790 2.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 974.425 655.605 974.595 703.715 ;
        RECT 974.425 524.365 974.595 572.475 ;
        RECT 974.425 427.805 974.595 475.915 ;
        RECT 974.425 331.245 974.595 386.155 ;
        RECT 974.425 83.045 974.595 131.155 ;
      LAYER mcon ;
        RECT 974.425 703.545 974.595 703.715 ;
        RECT 974.425 572.305 974.595 572.475 ;
        RECT 974.425 475.745 974.595 475.915 ;
        RECT 974.425 385.985 974.595 386.155 ;
        RECT 974.425 130.985 974.595 131.155 ;
      LAYER met1 ;
        RECT 973.430 1081.780 973.750 1081.840 ;
        RECT 977.570 1081.780 977.890 1081.840 ;
        RECT 973.430 1081.640 977.890 1081.780 ;
        RECT 973.430 1081.580 973.750 1081.640 ;
        RECT 977.570 1081.580 977.890 1081.640 ;
        RECT 973.430 1054.580 973.750 1054.640 ;
        RECT 975.730 1054.580 976.050 1054.640 ;
        RECT 973.430 1054.440 976.050 1054.580 ;
        RECT 973.430 1054.380 973.750 1054.440 ;
        RECT 975.730 1054.380 976.050 1054.440 ;
        RECT 974.810 862.820 975.130 862.880 ;
        RECT 975.270 862.820 975.590 862.880 ;
        RECT 974.810 862.680 975.590 862.820 ;
        RECT 974.810 862.620 975.130 862.680 ;
        RECT 975.270 862.620 975.590 862.680 ;
        RECT 974.365 703.700 974.655 703.745 ;
        RECT 974.810 703.700 975.130 703.760 ;
        RECT 974.365 703.560 975.130 703.700 ;
        RECT 974.365 703.515 974.655 703.560 ;
        RECT 974.810 703.500 975.130 703.560 ;
        RECT 974.350 655.760 974.670 655.820 ;
        RECT 974.155 655.620 974.670 655.760 ;
        RECT 974.350 655.560 974.670 655.620 ;
        RECT 974.350 621.080 974.670 621.140 ;
        RECT 974.810 621.080 975.130 621.140 ;
        RECT 974.350 620.940 975.130 621.080 ;
        RECT 974.350 620.880 974.670 620.940 ;
        RECT 974.810 620.880 975.130 620.940 ;
        RECT 974.810 579.940 975.130 580.000 ;
        RECT 974.440 579.800 975.130 579.940 ;
        RECT 974.440 579.660 974.580 579.800 ;
        RECT 974.810 579.740 975.130 579.800 ;
        RECT 974.350 579.400 974.670 579.660 ;
        RECT 974.350 572.460 974.670 572.520 ;
        RECT 974.155 572.320 974.670 572.460 ;
        RECT 974.350 572.260 974.670 572.320 ;
        RECT 974.365 524.520 974.655 524.565 ;
        RECT 974.810 524.520 975.130 524.580 ;
        RECT 974.365 524.380 975.130 524.520 ;
        RECT 974.365 524.335 974.655 524.380 ;
        RECT 974.810 524.320 975.130 524.380 ;
        RECT 974.365 475.900 974.655 475.945 ;
        RECT 974.810 475.900 975.130 475.960 ;
        RECT 974.365 475.760 975.130 475.900 ;
        RECT 974.365 475.715 974.655 475.760 ;
        RECT 974.810 475.700 975.130 475.760 ;
        RECT 974.350 427.960 974.670 428.020 ;
        RECT 974.155 427.820 974.670 427.960 ;
        RECT 974.350 427.760 974.670 427.820 ;
        RECT 974.350 386.140 974.670 386.200 ;
        RECT 974.155 386.000 974.670 386.140 ;
        RECT 974.350 385.940 974.670 386.000 ;
        RECT 974.365 331.400 974.655 331.445 ;
        RECT 974.810 331.400 975.130 331.460 ;
        RECT 974.365 331.260 975.130 331.400 ;
        RECT 974.365 331.215 974.655 331.260 ;
        RECT 974.810 331.200 975.130 331.260 ;
        RECT 974.810 234.500 975.130 234.560 ;
        RECT 975.730 234.500 976.050 234.560 ;
        RECT 974.810 234.360 976.050 234.500 ;
        RECT 974.810 234.300 975.130 234.360 ;
        RECT 975.730 234.300 976.050 234.360 ;
        RECT 974.350 131.140 974.670 131.200 ;
        RECT 974.155 131.000 974.670 131.140 ;
        RECT 974.350 130.940 974.670 131.000 ;
        RECT 974.365 83.200 974.655 83.245 ;
        RECT 974.810 83.200 975.130 83.260 ;
        RECT 974.365 83.060 975.130 83.200 ;
        RECT 974.365 83.015 974.655 83.060 ;
        RECT 974.810 83.000 975.130 83.060 ;
        RECT 372.210 52.260 372.530 52.320 ;
        RECT 974.350 52.260 974.670 52.320 ;
        RECT 372.210 52.120 974.670 52.260 ;
        RECT 372.210 52.060 372.530 52.120 ;
        RECT 974.350 52.060 974.670 52.120 ;
      LAYER via ;
        RECT 973.460 1081.580 973.720 1081.840 ;
        RECT 977.600 1081.580 977.860 1081.840 ;
        RECT 973.460 1054.380 973.720 1054.640 ;
        RECT 975.760 1054.380 976.020 1054.640 ;
        RECT 974.840 862.620 975.100 862.880 ;
        RECT 975.300 862.620 975.560 862.880 ;
        RECT 974.840 703.500 975.100 703.760 ;
        RECT 974.380 655.560 974.640 655.820 ;
        RECT 974.380 620.880 974.640 621.140 ;
        RECT 974.840 620.880 975.100 621.140 ;
        RECT 974.840 579.740 975.100 580.000 ;
        RECT 974.380 579.400 974.640 579.660 ;
        RECT 974.380 572.260 974.640 572.520 ;
        RECT 974.840 524.320 975.100 524.580 ;
        RECT 974.840 475.700 975.100 475.960 ;
        RECT 974.380 427.760 974.640 428.020 ;
        RECT 974.380 385.940 974.640 386.200 ;
        RECT 974.840 331.200 975.100 331.460 ;
        RECT 974.840 234.300 975.100 234.560 ;
        RECT 975.760 234.300 976.020 234.560 ;
        RECT 974.380 130.940 974.640 131.200 ;
        RECT 974.840 83.000 975.100 83.260 ;
        RECT 372.240 52.060 372.500 52.320 ;
        RECT 974.380 52.060 974.640 52.320 ;
      LAYER met2 ;
        RECT 977.510 1100.580 977.790 1104.000 ;
        RECT 977.510 1100.000 977.800 1100.580 ;
        RECT 977.660 1081.870 977.800 1100.000 ;
        RECT 973.460 1081.550 973.720 1081.870 ;
        RECT 977.600 1081.550 977.860 1081.870 ;
        RECT 973.520 1054.670 973.660 1081.550 ;
        RECT 973.460 1054.350 973.720 1054.670 ;
        RECT 975.760 1054.350 976.020 1054.670 ;
        RECT 975.820 959.210 975.960 1054.350 ;
        RECT 974.900 959.070 975.960 959.210 ;
        RECT 974.900 934.730 975.040 959.070 ;
        RECT 974.900 934.590 975.500 934.730 ;
        RECT 975.360 862.910 975.500 934.590 ;
        RECT 974.840 862.590 975.100 862.910 ;
        RECT 975.300 862.590 975.560 862.910 ;
        RECT 974.900 773.685 975.040 862.590 ;
        RECT 974.830 773.315 975.110 773.685 ;
        RECT 974.830 772.635 975.110 773.005 ;
        RECT 974.900 717.925 975.040 772.635 ;
        RECT 974.830 717.555 975.110 717.925 ;
        RECT 974.830 710.755 975.110 711.125 ;
        RECT 974.900 703.790 975.040 710.755 ;
        RECT 974.840 703.470 975.100 703.790 ;
        RECT 974.380 655.530 974.640 655.850 ;
        RECT 974.440 621.170 974.580 655.530 ;
        RECT 974.380 620.850 974.640 621.170 ;
        RECT 974.840 620.850 975.100 621.170 ;
        RECT 974.900 580.030 975.040 620.850 ;
        RECT 974.840 579.710 975.100 580.030 ;
        RECT 974.380 579.370 974.640 579.690 ;
        RECT 974.440 572.550 974.580 579.370 ;
        RECT 974.380 572.230 974.640 572.550 ;
        RECT 974.840 524.290 975.100 524.610 ;
        RECT 974.900 475.990 975.040 524.290 ;
        RECT 974.840 475.670 975.100 475.990 ;
        RECT 974.380 427.730 974.640 428.050 ;
        RECT 974.440 386.230 974.580 427.730 ;
        RECT 974.380 385.910 974.640 386.230 ;
        RECT 974.840 331.170 975.100 331.490 ;
        RECT 974.900 331.005 975.040 331.170 ;
        RECT 974.830 330.635 975.110 331.005 ;
        RECT 974.370 289.155 974.650 289.525 ;
        RECT 974.440 265.610 974.580 289.155 ;
        RECT 974.440 265.470 975.040 265.610 ;
        RECT 974.900 234.590 975.040 265.470 ;
        RECT 974.840 234.270 975.100 234.590 ;
        RECT 975.760 234.270 976.020 234.590 ;
        RECT 975.820 186.845 975.960 234.270 ;
        RECT 975.750 186.475 976.030 186.845 ;
        RECT 974.370 185.795 974.650 186.165 ;
        RECT 974.440 131.230 974.580 185.795 ;
        RECT 974.380 130.910 974.640 131.230 ;
        RECT 974.840 82.970 975.100 83.290 ;
        RECT 974.900 62.290 975.040 82.970 ;
        RECT 974.440 62.150 975.040 62.290 ;
        RECT 974.440 52.350 974.580 62.150 ;
        RECT 372.240 52.030 372.500 52.350 ;
        RECT 974.380 52.030 974.640 52.350 ;
        RECT 372.300 17.410 372.440 52.030 ;
        RECT 371.380 17.270 372.440 17.410 ;
        RECT 371.380 2.000 371.520 17.270 ;
        RECT 371.170 -4.000 371.730 2.000 ;
      LAYER via2 ;
        RECT 974.830 773.360 975.110 773.640 ;
        RECT 974.830 772.680 975.110 772.960 ;
        RECT 974.830 717.600 975.110 717.880 ;
        RECT 974.830 710.800 975.110 711.080 ;
        RECT 974.830 330.680 975.110 330.960 ;
        RECT 974.370 289.200 974.650 289.480 ;
        RECT 975.750 186.520 976.030 186.800 ;
        RECT 974.370 185.840 974.650 186.120 ;
      LAYER met3 ;
        RECT 974.805 773.650 975.135 773.665 ;
        RECT 974.805 773.350 975.810 773.650 ;
        RECT 974.805 773.335 975.135 773.350 ;
        RECT 974.805 772.970 975.135 772.985 ;
        RECT 975.510 772.970 975.810 773.350 ;
        RECT 974.805 772.670 975.810 772.970 ;
        RECT 974.805 772.655 975.135 772.670 ;
        RECT 974.805 717.900 975.135 717.905 ;
        RECT 974.550 717.890 975.135 717.900 ;
        RECT 974.350 717.590 975.135 717.890 ;
        RECT 974.550 717.580 975.135 717.590 ;
        RECT 974.805 717.575 975.135 717.580 ;
        RECT 974.805 711.100 975.135 711.105 ;
        RECT 974.550 711.090 975.135 711.100 ;
        RECT 974.550 710.790 975.360 711.090 ;
        RECT 974.550 710.780 975.135 710.790 ;
        RECT 974.805 710.775 975.135 710.780 ;
        RECT 974.805 330.970 975.135 330.985 ;
        RECT 975.470 330.970 975.850 330.980 ;
        RECT 974.805 330.670 975.850 330.970 ;
        RECT 974.805 330.655 975.135 330.670 ;
        RECT 975.470 330.660 975.850 330.670 ;
        RECT 974.345 289.490 974.675 289.505 ;
        RECT 975.470 289.490 975.850 289.500 ;
        RECT 974.345 289.190 975.850 289.490 ;
        RECT 974.345 289.175 974.675 289.190 ;
        RECT 975.470 289.180 975.850 289.190 ;
        RECT 975.725 186.810 976.055 186.825 ;
        RECT 975.510 186.495 976.055 186.810 ;
        RECT 974.345 186.130 974.675 186.145 ;
        RECT 975.510 186.130 975.810 186.495 ;
        RECT 974.345 185.830 975.810 186.130 ;
        RECT 974.345 185.815 974.675 185.830 ;
      LAYER via3 ;
        RECT 974.580 717.580 974.900 717.900 ;
        RECT 974.580 710.780 974.900 711.100 ;
        RECT 975.500 330.660 975.820 330.980 ;
        RECT 975.500 289.180 975.820 289.500 ;
      LAYER met4 ;
        RECT 974.575 717.575 974.905 717.905 ;
        RECT 974.590 711.105 974.890 717.575 ;
        RECT 974.575 710.775 974.905 711.105 ;
        RECT 975.495 330.655 975.825 330.985 ;
        RECT 975.510 289.505 975.810 330.655 ;
        RECT 975.495 289.175 975.825 289.505 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 980.330 1028.400 980.650 1028.460 ;
        RECT 981.710 1028.400 982.030 1028.460 ;
        RECT 980.330 1028.260 982.030 1028.400 ;
        RECT 980.330 1028.200 980.650 1028.260 ;
        RECT 981.710 1028.200 982.030 1028.260 ;
        RECT 980.330 159.160 980.650 159.420 ;
        RECT 980.420 158.740 980.560 159.160 ;
        RECT 980.330 158.480 980.650 158.740 ;
        RECT 392.910 52.600 393.230 52.660 ;
        RECT 979.870 52.600 980.190 52.660 ;
        RECT 392.910 52.460 980.190 52.600 ;
        RECT 392.910 52.400 393.230 52.460 ;
        RECT 979.870 52.400 980.190 52.460 ;
        RECT 389.230 16.560 389.550 16.620 ;
        RECT 392.910 16.560 393.230 16.620 ;
        RECT 389.230 16.420 393.230 16.560 ;
        RECT 389.230 16.360 389.550 16.420 ;
        RECT 392.910 16.360 393.230 16.420 ;
      LAYER via ;
        RECT 980.360 1028.200 980.620 1028.460 ;
        RECT 981.740 1028.200 982.000 1028.460 ;
        RECT 980.360 159.160 980.620 159.420 ;
        RECT 980.360 158.480 980.620 158.740 ;
        RECT 392.940 52.400 393.200 52.660 ;
        RECT 979.900 52.400 980.160 52.660 ;
        RECT 389.260 16.360 389.520 16.620 ;
        RECT 392.940 16.360 393.200 16.620 ;
      LAYER met2 ;
        RECT 983.490 1100.650 983.770 1104.000 ;
        RECT 981.800 1100.510 983.770 1100.650 ;
        RECT 981.800 1028.490 981.940 1100.510 ;
        RECT 983.490 1100.000 983.770 1100.510 ;
        RECT 980.360 1028.170 980.620 1028.490 ;
        RECT 981.740 1028.170 982.000 1028.490 ;
        RECT 980.420 980.290 980.560 1028.170 ;
        RECT 979.960 980.150 980.560 980.290 ;
        RECT 979.960 979.610 980.100 980.150 ;
        RECT 979.960 979.470 980.560 979.610 ;
        RECT 980.420 835.450 980.560 979.470 ;
        RECT 979.960 835.310 980.560 835.450 ;
        RECT 979.960 834.770 980.100 835.310 ;
        RECT 979.960 834.630 980.560 834.770 ;
        RECT 980.420 738.890 980.560 834.630 ;
        RECT 979.960 738.750 980.560 738.890 ;
        RECT 979.960 738.210 980.100 738.750 ;
        RECT 979.960 738.070 980.560 738.210 ;
        RECT 980.420 642.330 980.560 738.070 ;
        RECT 979.960 642.190 980.560 642.330 ;
        RECT 979.960 641.650 980.100 642.190 ;
        RECT 979.960 641.510 980.560 641.650 ;
        RECT 980.420 545.770 980.560 641.510 ;
        RECT 979.960 545.630 980.560 545.770 ;
        RECT 979.960 545.090 980.100 545.630 ;
        RECT 979.960 544.950 980.560 545.090 ;
        RECT 980.420 449.210 980.560 544.950 ;
        RECT 979.960 449.070 980.560 449.210 ;
        RECT 979.960 448.530 980.100 449.070 ;
        RECT 979.960 448.390 980.560 448.530 ;
        RECT 980.420 351.970 980.560 448.390 ;
        RECT 979.960 351.830 980.560 351.970 ;
        RECT 979.960 351.290 980.100 351.830 ;
        RECT 979.960 351.150 980.560 351.290 ;
        RECT 980.420 255.410 980.560 351.150 ;
        RECT 979.960 255.270 980.560 255.410 ;
        RECT 979.960 254.730 980.100 255.270 ;
        RECT 979.960 254.590 980.560 254.730 ;
        RECT 980.420 159.450 980.560 254.590 ;
        RECT 980.360 159.130 980.620 159.450 ;
        RECT 980.360 158.450 980.620 158.770 ;
        RECT 980.420 62.290 980.560 158.450 ;
        RECT 979.960 62.150 980.560 62.290 ;
        RECT 979.960 52.690 980.100 62.150 ;
        RECT 392.940 52.370 393.200 52.690 ;
        RECT 979.900 52.370 980.160 52.690 ;
        RECT 393.000 16.650 393.140 52.370 ;
        RECT 389.260 16.330 389.520 16.650 ;
        RECT 392.940 16.330 393.200 16.650 ;
        RECT 389.320 2.000 389.460 16.330 ;
        RECT 389.110 -4.000 389.670 2.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 987.230 1028.740 987.550 1028.800 ;
        RECT 988.150 1028.740 988.470 1028.800 ;
        RECT 987.230 1028.600 988.470 1028.740 ;
        RECT 987.230 1028.540 987.550 1028.600 ;
        RECT 988.150 1028.540 988.470 1028.600 ;
        RECT 413.610 52.940 413.930 53.000 ;
        RECT 987.230 52.940 987.550 53.000 ;
        RECT 413.610 52.800 987.550 52.940 ;
        RECT 413.610 52.740 413.930 52.800 ;
        RECT 987.230 52.740 987.550 52.800 ;
        RECT 407.170 16.560 407.490 16.620 ;
        RECT 413.610 16.560 413.930 16.620 ;
        RECT 407.170 16.420 413.930 16.560 ;
        RECT 407.170 16.360 407.490 16.420 ;
        RECT 413.610 16.360 413.930 16.420 ;
      LAYER via ;
        RECT 987.260 1028.540 987.520 1028.800 ;
        RECT 988.180 1028.540 988.440 1028.800 ;
        RECT 413.640 52.740 413.900 53.000 ;
        RECT 987.260 52.740 987.520 53.000 ;
        RECT 407.200 16.360 407.460 16.620 ;
        RECT 413.640 16.360 413.900 16.620 ;
      LAYER met2 ;
        RECT 989.470 1100.650 989.750 1104.000 ;
        RECT 988.240 1100.510 989.750 1100.650 ;
        RECT 988.240 1028.830 988.380 1100.510 ;
        RECT 989.470 1100.000 989.750 1100.510 ;
        RECT 987.260 1028.510 987.520 1028.830 ;
        RECT 988.180 1028.510 988.440 1028.830 ;
        RECT 987.320 53.030 987.460 1028.510 ;
        RECT 413.640 52.710 413.900 53.030 ;
        RECT 987.260 52.710 987.520 53.030 ;
        RECT 413.700 16.650 413.840 52.710 ;
        RECT 407.200 16.330 407.460 16.650 ;
        RECT 413.640 16.330 413.900 16.650 ;
        RECT 407.260 2.000 407.400 16.330 ;
        RECT 407.050 -4.000 407.610 2.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 869.930 1076.680 870.250 1076.740 ;
        RECT 873.150 1076.680 873.470 1076.740 ;
        RECT 869.930 1076.540 873.470 1076.680 ;
        RECT 869.930 1076.480 870.250 1076.540 ;
        RECT 873.150 1076.480 873.470 1076.540 ;
        RECT 68.150 44.780 68.470 44.840 ;
        RECT 869.930 44.780 870.250 44.840 ;
        RECT 68.150 44.640 870.250 44.780 ;
        RECT 68.150 44.580 68.470 44.640 ;
        RECT 869.930 44.580 870.250 44.640 ;
      LAYER via ;
        RECT 869.960 1076.480 870.220 1076.740 ;
        RECT 873.180 1076.480 873.440 1076.740 ;
        RECT 68.180 44.580 68.440 44.840 ;
        RECT 869.960 44.580 870.220 44.840 ;
      LAYER met2 ;
        RECT 873.090 1100.580 873.370 1104.000 ;
        RECT 873.090 1100.000 873.380 1100.580 ;
        RECT 873.240 1076.770 873.380 1100.000 ;
        RECT 869.960 1076.450 870.220 1076.770 ;
        RECT 873.180 1076.450 873.440 1076.770 ;
        RECT 870.020 44.870 870.160 1076.450 ;
        RECT 68.180 44.550 68.440 44.870 ;
        RECT 869.960 44.550 870.220 44.870 ;
        RECT 68.240 2.000 68.380 44.550 ;
        RECT 68.030 -4.000 68.590 2.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 427.410 53.280 427.730 53.340 ;
        RECT 994.590 53.280 994.910 53.340 ;
        RECT 427.410 53.140 994.910 53.280 ;
        RECT 427.410 53.080 427.730 53.140 ;
        RECT 994.590 53.080 994.910 53.140 ;
        RECT 424.650 16.220 424.970 16.280 ;
        RECT 427.410 16.220 427.730 16.280 ;
        RECT 424.650 16.080 427.730 16.220 ;
        RECT 424.650 16.020 424.970 16.080 ;
        RECT 427.410 16.020 427.730 16.080 ;
      LAYER via ;
        RECT 427.440 53.080 427.700 53.340 ;
        RECT 994.620 53.080 994.880 53.340 ;
        RECT 424.680 16.020 424.940 16.280 ;
        RECT 427.440 16.020 427.700 16.280 ;
      LAYER met2 ;
        RECT 995.910 1100.650 996.190 1104.000 ;
        RECT 994.680 1100.510 996.190 1100.650 ;
        RECT 994.680 53.370 994.820 1100.510 ;
        RECT 995.910 1100.000 996.190 1100.510 ;
        RECT 427.440 53.050 427.700 53.370 ;
        RECT 994.620 53.050 994.880 53.370 ;
        RECT 427.500 16.310 427.640 53.050 ;
        RECT 424.680 15.990 424.940 16.310 ;
        RECT 427.440 15.990 427.700 16.310 ;
        RECT 424.740 2.000 424.880 15.990 ;
        RECT 424.530 -4.000 425.090 2.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 448.110 53.620 448.430 53.680 ;
        RECT 1001.030 53.620 1001.350 53.680 ;
        RECT 448.110 53.480 1001.350 53.620 ;
        RECT 448.110 53.420 448.430 53.480 ;
        RECT 1001.030 53.420 1001.350 53.480 ;
        RECT 442.590 15.880 442.910 15.940 ;
        RECT 448.110 15.880 448.430 15.940 ;
        RECT 442.590 15.740 448.430 15.880 ;
        RECT 442.590 15.680 442.910 15.740 ;
        RECT 448.110 15.680 448.430 15.740 ;
      LAYER via ;
        RECT 448.140 53.420 448.400 53.680 ;
        RECT 1001.060 53.420 1001.320 53.680 ;
        RECT 442.620 15.680 442.880 15.940 ;
        RECT 448.140 15.680 448.400 15.940 ;
      LAYER met2 ;
        RECT 1001.890 1100.650 1002.170 1104.000 ;
        RECT 1001.120 1100.510 1002.170 1100.650 ;
        RECT 1001.120 53.710 1001.260 1100.510 ;
        RECT 1001.890 1100.000 1002.170 1100.510 ;
        RECT 448.140 53.390 448.400 53.710 ;
        RECT 1001.060 53.390 1001.320 53.710 ;
        RECT 448.200 15.970 448.340 53.390 ;
        RECT 442.620 15.650 442.880 15.970 ;
        RECT 448.140 15.650 448.400 15.970 ;
        RECT 442.680 2.000 442.820 15.650 ;
        RECT 442.470 -4.000 443.030 2.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 461.910 53.960 462.230 54.020 ;
        RECT 1007.930 53.960 1008.250 54.020 ;
        RECT 461.910 53.820 1008.250 53.960 ;
        RECT 461.910 53.760 462.230 53.820 ;
        RECT 1007.930 53.760 1008.250 53.820 ;
      LAYER via ;
        RECT 461.940 53.760 462.200 54.020 ;
        RECT 1007.960 53.760 1008.220 54.020 ;
      LAYER met2 ;
        RECT 1007.870 1100.580 1008.150 1104.000 ;
        RECT 1007.870 1100.000 1008.160 1100.580 ;
        RECT 1008.020 54.050 1008.160 1100.000 ;
        RECT 461.940 53.730 462.200 54.050 ;
        RECT 1007.960 53.730 1008.220 54.050 ;
        RECT 462.000 16.730 462.140 53.730 ;
        RECT 460.620 16.590 462.140 16.730 ;
        RECT 460.620 2.000 460.760 16.590 ;
        RECT 460.410 -4.000 460.970 2.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1008.390 1052.200 1008.710 1052.260 ;
        RECT 1012.530 1052.200 1012.850 1052.260 ;
        RECT 1008.390 1052.060 1012.850 1052.200 ;
        RECT 1008.390 1052.000 1008.710 1052.060 ;
        RECT 1012.530 1052.000 1012.850 1052.060 ;
        RECT 482.610 54.300 482.930 54.360 ;
        RECT 1008.390 54.300 1008.710 54.360 ;
        RECT 482.610 54.160 1008.710 54.300 ;
        RECT 482.610 54.100 482.930 54.160 ;
        RECT 1008.390 54.100 1008.710 54.160 ;
        RECT 478.470 15.200 478.790 15.260 ;
        RECT 482.610 15.200 482.930 15.260 ;
        RECT 478.470 15.060 482.930 15.200 ;
        RECT 478.470 15.000 478.790 15.060 ;
        RECT 482.610 15.000 482.930 15.060 ;
      LAYER via ;
        RECT 1008.420 1052.000 1008.680 1052.260 ;
        RECT 1012.560 1052.000 1012.820 1052.260 ;
        RECT 482.640 54.100 482.900 54.360 ;
        RECT 1008.420 54.100 1008.680 54.360 ;
        RECT 478.500 15.000 478.760 15.260 ;
        RECT 482.640 15.000 482.900 15.260 ;
      LAYER met2 ;
        RECT 1013.850 1100.650 1014.130 1104.000 ;
        RECT 1012.620 1100.510 1014.130 1100.650 ;
        RECT 1012.620 1052.290 1012.760 1100.510 ;
        RECT 1013.850 1100.000 1014.130 1100.510 ;
        RECT 1008.420 1051.970 1008.680 1052.290 ;
        RECT 1012.560 1051.970 1012.820 1052.290 ;
        RECT 1008.480 54.390 1008.620 1051.970 ;
        RECT 482.640 54.070 482.900 54.390 ;
        RECT 1008.420 54.070 1008.680 54.390 ;
        RECT 482.700 15.290 482.840 54.070 ;
        RECT 478.500 14.970 478.760 15.290 ;
        RECT 482.640 14.970 482.900 15.290 ;
        RECT 478.560 2.000 478.700 14.970 ;
        RECT 478.350 -4.000 478.910 2.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1014.830 1052.200 1015.150 1052.260 ;
        RECT 1018.510 1052.200 1018.830 1052.260 ;
        RECT 1014.830 1052.060 1018.830 1052.200 ;
        RECT 1014.830 1052.000 1015.150 1052.060 ;
        RECT 1018.510 1052.000 1018.830 1052.060 ;
        RECT 496.410 54.640 496.730 54.700 ;
        RECT 1014.830 54.640 1015.150 54.700 ;
        RECT 496.410 54.500 1015.150 54.640 ;
        RECT 496.410 54.440 496.730 54.500 ;
        RECT 1014.830 54.440 1015.150 54.500 ;
      LAYER via ;
        RECT 1014.860 1052.000 1015.120 1052.260 ;
        RECT 1018.540 1052.000 1018.800 1052.260 ;
        RECT 496.440 54.440 496.700 54.700 ;
        RECT 1014.860 54.440 1015.120 54.700 ;
      LAYER met2 ;
        RECT 1020.290 1100.650 1020.570 1104.000 ;
        RECT 1018.600 1100.510 1020.570 1100.650 ;
        RECT 1018.600 1052.290 1018.740 1100.510 ;
        RECT 1020.290 1100.000 1020.570 1100.510 ;
        RECT 1014.860 1051.970 1015.120 1052.290 ;
        RECT 1018.540 1051.970 1018.800 1052.290 ;
        RECT 1014.920 54.730 1015.060 1051.970 ;
        RECT 496.440 54.410 496.700 54.730 ;
        RECT 1014.860 54.410 1015.120 54.730 ;
        RECT 496.500 2.000 496.640 54.410 ;
        RECT 496.290 -4.000 496.850 2.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1021.730 1052.200 1022.050 1052.260 ;
        RECT 1024.950 1052.200 1025.270 1052.260 ;
        RECT 1021.730 1052.060 1025.270 1052.200 ;
        RECT 1021.730 1052.000 1022.050 1052.060 ;
        RECT 1024.950 1052.000 1025.270 1052.060 ;
        RECT 517.110 54.980 517.430 55.040 ;
        RECT 1021.730 54.980 1022.050 55.040 ;
        RECT 517.110 54.840 1022.050 54.980 ;
        RECT 517.110 54.780 517.430 54.840 ;
        RECT 1021.730 54.780 1022.050 54.840 ;
        RECT 513.890 15.200 514.210 15.260 ;
        RECT 517.110 15.200 517.430 15.260 ;
        RECT 513.890 15.060 517.430 15.200 ;
        RECT 513.890 15.000 514.210 15.060 ;
        RECT 517.110 15.000 517.430 15.060 ;
      LAYER via ;
        RECT 1021.760 1052.000 1022.020 1052.260 ;
        RECT 1024.980 1052.000 1025.240 1052.260 ;
        RECT 517.140 54.780 517.400 55.040 ;
        RECT 1021.760 54.780 1022.020 55.040 ;
        RECT 513.920 15.000 514.180 15.260 ;
        RECT 517.140 15.000 517.400 15.260 ;
      LAYER met2 ;
        RECT 1026.270 1100.650 1026.550 1104.000 ;
        RECT 1025.040 1100.510 1026.550 1100.650 ;
        RECT 1025.040 1052.290 1025.180 1100.510 ;
        RECT 1026.270 1100.000 1026.550 1100.510 ;
        RECT 1021.760 1051.970 1022.020 1052.290 ;
        RECT 1024.980 1051.970 1025.240 1052.290 ;
        RECT 1021.820 55.070 1021.960 1051.970 ;
        RECT 517.140 54.750 517.400 55.070 ;
        RECT 1021.760 54.750 1022.020 55.070 ;
        RECT 517.200 15.290 517.340 54.750 ;
        RECT 513.920 14.970 514.180 15.290 ;
        RECT 517.140 14.970 517.400 15.290 ;
        RECT 513.980 2.000 514.120 14.970 ;
        RECT 513.770 -4.000 514.330 2.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1028.630 1072.940 1028.950 1073.000 ;
        RECT 1030.930 1072.940 1031.250 1073.000 ;
        RECT 1028.630 1072.800 1031.250 1072.940 ;
        RECT 1028.630 1072.740 1028.950 1072.800 ;
        RECT 1030.930 1072.740 1031.250 1072.800 ;
        RECT 537.810 51.240 538.130 51.300 ;
        RECT 1028.630 51.240 1028.950 51.300 ;
        RECT 537.810 51.100 1028.950 51.240 ;
        RECT 537.810 51.040 538.130 51.100 ;
        RECT 1028.630 51.040 1028.950 51.100 ;
        RECT 531.830 15.200 532.150 15.260 ;
        RECT 537.810 15.200 538.130 15.260 ;
        RECT 531.830 15.060 538.130 15.200 ;
        RECT 531.830 15.000 532.150 15.060 ;
        RECT 537.810 15.000 538.130 15.060 ;
      LAYER via ;
        RECT 1028.660 1072.740 1028.920 1073.000 ;
        RECT 1030.960 1072.740 1031.220 1073.000 ;
        RECT 537.840 51.040 538.100 51.300 ;
        RECT 1028.660 51.040 1028.920 51.300 ;
        RECT 531.860 15.000 532.120 15.260 ;
        RECT 537.840 15.000 538.100 15.260 ;
      LAYER met2 ;
        RECT 1032.250 1100.650 1032.530 1104.000 ;
        RECT 1031.020 1100.510 1032.530 1100.650 ;
        RECT 1031.020 1073.030 1031.160 1100.510 ;
        RECT 1032.250 1100.000 1032.530 1100.510 ;
        RECT 1028.660 1072.710 1028.920 1073.030 ;
        RECT 1030.960 1072.710 1031.220 1073.030 ;
        RECT 1028.720 51.330 1028.860 1072.710 ;
        RECT 537.840 51.010 538.100 51.330 ;
        RECT 1028.660 51.010 1028.920 51.330 ;
        RECT 537.900 15.290 538.040 51.010 ;
        RECT 531.860 14.970 532.120 15.290 ;
        RECT 537.840 14.970 538.100 15.290 ;
        RECT 531.920 2.000 532.060 14.970 ;
        RECT 531.710 -4.000 532.270 2.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1035.530 1049.140 1035.850 1049.200 ;
        RECT 1036.910 1049.140 1037.230 1049.200 ;
        RECT 1035.530 1049.000 1037.230 1049.140 ;
        RECT 1035.530 1048.940 1035.850 1049.000 ;
        RECT 1036.910 1048.940 1037.230 1049.000 ;
        RECT 551.610 50.900 551.930 50.960 ;
        RECT 1035.530 50.900 1035.850 50.960 ;
        RECT 551.610 50.760 1035.850 50.900 ;
        RECT 551.610 50.700 551.930 50.760 ;
        RECT 1035.530 50.700 1035.850 50.760 ;
      LAYER via ;
        RECT 1035.560 1048.940 1035.820 1049.200 ;
        RECT 1036.940 1048.940 1037.200 1049.200 ;
        RECT 551.640 50.700 551.900 50.960 ;
        RECT 1035.560 50.700 1035.820 50.960 ;
      LAYER met2 ;
        RECT 1038.690 1100.650 1038.970 1104.000 ;
        RECT 1037.000 1100.510 1038.970 1100.650 ;
        RECT 1037.000 1049.230 1037.140 1100.510 ;
        RECT 1038.690 1100.000 1038.970 1100.510 ;
        RECT 1035.560 1048.910 1035.820 1049.230 ;
        RECT 1036.940 1048.910 1037.200 1049.230 ;
        RECT 1035.620 50.990 1035.760 1048.910 ;
        RECT 551.640 50.670 551.900 50.990 ;
        RECT 1035.560 50.670 1035.820 50.990 ;
        RECT 551.700 17.410 551.840 50.670 ;
        RECT 549.860 17.270 551.840 17.410 ;
        RECT 549.860 2.000 550.000 17.270 ;
        RECT 549.650 -4.000 550.210 2.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1042.430 1072.940 1042.750 1073.000 ;
        RECT 1043.350 1072.940 1043.670 1073.000 ;
        RECT 1042.430 1072.800 1043.670 1072.940 ;
        RECT 1042.430 1072.740 1042.750 1072.800 ;
        RECT 1043.350 1072.740 1043.670 1072.800 ;
        RECT 572.310 50.560 572.630 50.620 ;
        RECT 1042.430 50.560 1042.750 50.620 ;
        RECT 572.310 50.420 1042.750 50.560 ;
        RECT 572.310 50.360 572.630 50.420 ;
        RECT 1042.430 50.360 1042.750 50.420 ;
        RECT 567.710 14.860 568.030 14.920 ;
        RECT 572.310 14.860 572.630 14.920 ;
        RECT 567.710 14.720 572.630 14.860 ;
        RECT 567.710 14.660 568.030 14.720 ;
        RECT 572.310 14.660 572.630 14.720 ;
      LAYER via ;
        RECT 1042.460 1072.740 1042.720 1073.000 ;
        RECT 1043.380 1072.740 1043.640 1073.000 ;
        RECT 572.340 50.360 572.600 50.620 ;
        RECT 1042.460 50.360 1042.720 50.620 ;
        RECT 567.740 14.660 568.000 14.920 ;
        RECT 572.340 14.660 572.600 14.920 ;
      LAYER met2 ;
        RECT 1044.670 1100.650 1044.950 1104.000 ;
        RECT 1043.440 1100.510 1044.950 1100.650 ;
        RECT 1043.440 1073.030 1043.580 1100.510 ;
        RECT 1044.670 1100.000 1044.950 1100.510 ;
        RECT 1042.460 1072.710 1042.720 1073.030 ;
        RECT 1043.380 1072.710 1043.640 1073.030 ;
        RECT 1042.520 50.650 1042.660 1072.710 ;
        RECT 572.340 50.330 572.600 50.650 ;
        RECT 1042.460 50.330 1042.720 50.650 ;
        RECT 572.400 14.950 572.540 50.330 ;
        RECT 567.740 14.630 568.000 14.950 ;
        RECT 572.340 14.630 572.600 14.950 ;
        RECT 567.800 2.000 567.940 14.630 ;
        RECT 567.590 -4.000 568.150 2.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 900.825 1062.585 900.995 1088.595 ;
        RECT 899.905 897.005 900.075 945.115 ;
        RECT 899.905 655.945 900.075 703.715 ;
        RECT 899.905 462.485 900.075 510.595 ;
        RECT 899.905 365.925 900.075 414.035 ;
        RECT 899.905 269.025 900.075 317.475 ;
        RECT 899.905 179.605 900.075 227.715 ;
        RECT 899.905 83.045 900.075 131.155 ;
      LAYER mcon ;
        RECT 900.825 1088.425 900.995 1088.595 ;
        RECT 899.905 944.945 900.075 945.115 ;
        RECT 899.905 703.545 900.075 703.715 ;
        RECT 899.905 510.425 900.075 510.595 ;
        RECT 899.905 413.865 900.075 414.035 ;
        RECT 899.905 317.305 900.075 317.475 ;
        RECT 899.905 227.545 900.075 227.715 ;
        RECT 899.905 130.985 900.075 131.155 ;
      LAYER met1 ;
        RECT 900.765 1088.580 901.055 1088.625 ;
        RECT 1050.710 1088.580 1051.030 1088.640 ;
        RECT 900.765 1088.440 1051.030 1088.580 ;
        RECT 900.765 1088.395 901.055 1088.440 ;
        RECT 1050.710 1088.380 1051.030 1088.440 ;
        RECT 900.750 1062.740 901.070 1062.800 ;
        RECT 900.555 1062.600 901.070 1062.740 ;
        RECT 900.750 1062.540 901.070 1062.600 ;
        RECT 900.290 976.040 900.610 976.100 ;
        RECT 900.750 976.040 901.070 976.100 ;
        RECT 900.290 975.900 901.070 976.040 ;
        RECT 900.290 975.840 900.610 975.900 ;
        RECT 900.750 975.840 901.070 975.900 ;
        RECT 899.845 945.100 900.135 945.145 ;
        RECT 900.290 945.100 900.610 945.160 ;
        RECT 899.845 944.960 900.610 945.100 ;
        RECT 899.845 944.915 900.135 944.960 ;
        RECT 900.290 944.900 900.610 944.960 ;
        RECT 899.830 897.160 900.150 897.220 ;
        RECT 899.635 897.020 900.150 897.160 ;
        RECT 899.830 896.960 900.150 897.020 ;
        RECT 899.370 759.120 899.690 759.180 ;
        RECT 899.830 759.120 900.150 759.180 ;
        RECT 899.370 758.980 900.150 759.120 ;
        RECT 899.370 758.920 899.690 758.980 ;
        RECT 899.830 758.920 900.150 758.980 ;
        RECT 899.830 703.700 900.150 703.760 ;
        RECT 899.635 703.560 900.150 703.700 ;
        RECT 899.830 703.500 900.150 703.560 ;
        RECT 899.845 656.100 900.135 656.145 ;
        RECT 899.845 655.960 900.980 656.100 ;
        RECT 899.845 655.915 900.135 655.960 ;
        RECT 900.840 655.820 900.980 655.960 ;
        RECT 900.750 655.560 901.070 655.820 ;
        RECT 899.830 638.420 900.150 638.480 ;
        RECT 900.750 638.420 901.070 638.480 ;
        RECT 899.830 638.280 901.070 638.420 ;
        RECT 899.830 638.220 900.150 638.280 ;
        RECT 900.750 638.220 901.070 638.280 ;
        RECT 899.830 510.580 900.150 510.640 ;
        RECT 899.635 510.440 900.150 510.580 ;
        RECT 899.830 510.380 900.150 510.440 ;
        RECT 899.830 462.640 900.150 462.700 ;
        RECT 899.635 462.500 900.150 462.640 ;
        RECT 899.830 462.440 900.150 462.500 ;
        RECT 899.830 414.020 900.150 414.080 ;
        RECT 899.635 413.880 900.150 414.020 ;
        RECT 899.830 413.820 900.150 413.880 ;
        RECT 899.830 366.080 900.150 366.140 ;
        RECT 899.635 365.940 900.150 366.080 ;
        RECT 899.830 365.880 900.150 365.940 ;
        RECT 899.830 317.460 900.150 317.520 ;
        RECT 899.635 317.320 900.150 317.460 ;
        RECT 899.830 317.260 900.150 317.320 ;
        RECT 899.830 269.180 900.150 269.240 ;
        RECT 899.635 269.040 900.150 269.180 ;
        RECT 899.830 268.980 900.150 269.040 ;
        RECT 899.830 228.180 900.150 228.440 ;
        RECT 899.920 227.745 900.060 228.180 ;
        RECT 899.845 227.515 900.135 227.745 ;
        RECT 899.845 179.760 900.135 179.805 ;
        RECT 900.290 179.760 900.610 179.820 ;
        RECT 899.845 179.620 900.610 179.760 ;
        RECT 899.845 179.575 900.135 179.620 ;
        RECT 900.290 179.560 900.610 179.620 ;
        RECT 900.290 159.020 900.610 159.080 ;
        RECT 899.920 158.880 900.610 159.020 ;
        RECT 899.920 158.740 900.060 158.880 ;
        RECT 900.290 158.820 900.610 158.880 ;
        RECT 899.830 158.480 900.150 158.740 ;
        RECT 899.830 131.140 900.150 131.200 ;
        RECT 899.635 131.000 900.150 131.140 ;
        RECT 899.830 130.940 900.150 131.000 ;
        RECT 899.830 83.200 900.150 83.260 ;
        RECT 899.635 83.060 900.150 83.200 ;
        RECT 899.830 83.000 900.150 83.060 ;
        RECT 585.650 43.420 585.970 43.480 ;
        RECT 899.830 43.420 900.150 43.480 ;
        RECT 585.650 43.280 900.150 43.420 ;
        RECT 585.650 43.220 585.970 43.280 ;
        RECT 899.830 43.220 900.150 43.280 ;
      LAYER via ;
        RECT 1050.740 1088.380 1051.000 1088.640 ;
        RECT 900.780 1062.540 901.040 1062.800 ;
        RECT 900.320 975.840 900.580 976.100 ;
        RECT 900.780 975.840 901.040 976.100 ;
        RECT 900.320 944.900 900.580 945.160 ;
        RECT 899.860 896.960 900.120 897.220 ;
        RECT 899.400 758.920 899.660 759.180 ;
        RECT 899.860 758.920 900.120 759.180 ;
        RECT 899.860 703.500 900.120 703.760 ;
        RECT 900.780 655.560 901.040 655.820 ;
        RECT 899.860 638.220 900.120 638.480 ;
        RECT 900.780 638.220 901.040 638.480 ;
        RECT 899.860 510.380 900.120 510.640 ;
        RECT 899.860 462.440 900.120 462.700 ;
        RECT 899.860 413.820 900.120 414.080 ;
        RECT 899.860 365.880 900.120 366.140 ;
        RECT 899.860 317.260 900.120 317.520 ;
        RECT 899.860 268.980 900.120 269.240 ;
        RECT 899.860 228.180 900.120 228.440 ;
        RECT 900.320 179.560 900.580 179.820 ;
        RECT 900.320 158.820 900.580 159.080 ;
        RECT 899.860 158.480 900.120 158.740 ;
        RECT 899.860 130.940 900.120 131.200 ;
        RECT 899.860 83.000 900.120 83.260 ;
        RECT 585.680 43.220 585.940 43.480 ;
        RECT 899.860 43.220 900.120 43.480 ;
      LAYER met2 ;
        RECT 1050.650 1100.580 1050.930 1104.000 ;
        RECT 1050.650 1100.000 1050.940 1100.580 ;
        RECT 1050.800 1088.670 1050.940 1100.000 ;
        RECT 1050.740 1088.350 1051.000 1088.670 ;
        RECT 900.780 1062.510 901.040 1062.830 ;
        RECT 900.840 976.130 900.980 1062.510 ;
        RECT 900.320 975.810 900.580 976.130 ;
        RECT 900.780 975.810 901.040 976.130 ;
        RECT 900.380 945.190 900.520 975.810 ;
        RECT 900.320 944.870 900.580 945.190 ;
        RECT 899.860 896.930 900.120 897.250 ;
        RECT 899.920 896.650 900.060 896.930 ;
        RECT 899.920 896.510 900.520 896.650 ;
        RECT 900.380 883.730 900.520 896.510 ;
        RECT 899.460 883.590 900.520 883.730 ;
        RECT 899.460 759.210 899.600 883.590 ;
        RECT 899.400 758.890 899.660 759.210 ;
        RECT 899.860 758.890 900.120 759.210 ;
        RECT 899.920 703.790 900.060 758.890 ;
        RECT 899.860 703.470 900.120 703.790 ;
        RECT 900.780 655.530 901.040 655.850 ;
        RECT 900.840 638.510 900.980 655.530 ;
        RECT 899.860 638.190 900.120 638.510 ;
        RECT 900.780 638.190 901.040 638.510 ;
        RECT 899.920 510.670 900.060 638.190 ;
        RECT 899.860 510.350 900.120 510.670 ;
        RECT 899.860 462.410 900.120 462.730 ;
        RECT 899.920 414.110 900.060 462.410 ;
        RECT 899.860 413.790 900.120 414.110 ;
        RECT 899.860 365.850 900.120 366.170 ;
        RECT 899.920 317.550 900.060 365.850 ;
        RECT 899.860 317.230 900.120 317.550 ;
        RECT 899.860 268.950 900.120 269.270 ;
        RECT 899.920 228.470 900.060 268.950 ;
        RECT 899.860 228.150 900.120 228.470 ;
        RECT 900.320 179.530 900.580 179.850 ;
        RECT 900.380 159.110 900.520 179.530 ;
        RECT 900.320 158.790 900.580 159.110 ;
        RECT 899.860 158.450 900.120 158.770 ;
        RECT 899.920 131.230 900.060 158.450 ;
        RECT 899.860 130.910 900.120 131.230 ;
        RECT 899.860 82.970 900.120 83.290 ;
        RECT 899.920 43.510 900.060 82.970 ;
        RECT 585.680 43.190 585.940 43.510 ;
        RECT 899.860 43.190 900.120 43.510 ;
        RECT 585.740 2.000 585.880 43.190 ;
        RECT 585.530 -4.000 586.090 2.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 876.830 1052.200 877.150 1052.260 ;
        RECT 880.050 1052.200 880.370 1052.260 ;
        RECT 876.830 1052.060 880.370 1052.200 ;
        RECT 876.830 1052.000 877.150 1052.060 ;
        RECT 880.050 1052.000 880.370 1052.060 ;
        RECT 91.610 45.120 91.930 45.180 ;
        RECT 876.830 45.120 877.150 45.180 ;
        RECT 91.610 44.980 877.150 45.120 ;
        RECT 91.610 44.920 91.930 44.980 ;
        RECT 876.830 44.920 877.150 44.980 ;
      LAYER via ;
        RECT 876.860 1052.000 877.120 1052.260 ;
        RECT 880.080 1052.000 880.340 1052.260 ;
        RECT 91.640 44.920 91.900 45.180 ;
        RECT 876.860 44.920 877.120 45.180 ;
      LAYER met2 ;
        RECT 881.370 1100.650 881.650 1104.000 ;
        RECT 880.140 1100.510 881.650 1100.650 ;
        RECT 880.140 1052.290 880.280 1100.510 ;
        RECT 881.370 1100.000 881.650 1100.510 ;
        RECT 876.860 1051.970 877.120 1052.290 ;
        RECT 880.080 1051.970 880.340 1052.290 ;
        RECT 876.920 45.210 877.060 1051.970 ;
        RECT 91.640 44.890 91.900 45.210 ;
        RECT 876.860 44.890 877.120 45.210 ;
        RECT 91.700 2.000 91.840 44.890 ;
        RECT 91.490 -4.000 92.050 2.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 606.810 59.060 607.130 59.120 ;
        RECT 1056.230 59.060 1056.550 59.120 ;
        RECT 606.810 58.920 1056.550 59.060 ;
        RECT 606.810 58.860 607.130 58.920 ;
        RECT 1056.230 58.860 1056.550 58.920 ;
        RECT 603.130 14.860 603.450 14.920 ;
        RECT 606.810 14.860 607.130 14.920 ;
        RECT 603.130 14.720 607.130 14.860 ;
        RECT 603.130 14.660 603.450 14.720 ;
        RECT 606.810 14.660 607.130 14.720 ;
      LAYER via ;
        RECT 606.840 58.860 607.100 59.120 ;
        RECT 1056.260 58.860 1056.520 59.120 ;
        RECT 603.160 14.660 603.420 14.920 ;
        RECT 606.840 14.660 607.100 14.920 ;
      LAYER met2 ;
        RECT 1057.090 1100.650 1057.370 1104.000 ;
        RECT 1056.320 1100.510 1057.370 1100.650 ;
        RECT 1056.320 59.150 1056.460 1100.510 ;
        RECT 1057.090 1100.000 1057.370 1100.510 ;
        RECT 606.840 58.830 607.100 59.150 ;
        RECT 1056.260 58.830 1056.520 59.150 ;
        RECT 606.900 14.950 607.040 58.830 ;
        RECT 603.160 14.630 603.420 14.950 ;
        RECT 606.840 14.630 607.100 14.950 ;
        RECT 603.220 2.000 603.360 14.630 ;
        RECT 603.010 -4.000 603.570 2.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 627.510 59.400 627.830 59.460 ;
        RECT 1063.590 59.400 1063.910 59.460 ;
        RECT 627.510 59.260 1063.910 59.400 ;
        RECT 627.510 59.200 627.830 59.260 ;
        RECT 1063.590 59.200 1063.910 59.260 ;
        RECT 621.070 14.180 621.390 14.240 ;
        RECT 627.510 14.180 627.830 14.240 ;
        RECT 621.070 14.040 627.830 14.180 ;
        RECT 621.070 13.980 621.390 14.040 ;
        RECT 627.510 13.980 627.830 14.040 ;
      LAYER via ;
        RECT 627.540 59.200 627.800 59.460 ;
        RECT 1063.620 59.200 1063.880 59.460 ;
        RECT 621.100 13.980 621.360 14.240 ;
        RECT 627.540 13.980 627.800 14.240 ;
      LAYER met2 ;
        RECT 1063.070 1100.650 1063.350 1104.000 ;
        RECT 1063.070 1100.510 1063.820 1100.650 ;
        RECT 1063.070 1100.000 1063.350 1100.510 ;
        RECT 1063.680 59.490 1063.820 1100.510 ;
        RECT 627.540 59.170 627.800 59.490 ;
        RECT 1063.620 59.170 1063.880 59.490 ;
        RECT 627.600 14.270 627.740 59.170 ;
        RECT 621.100 13.950 621.360 14.270 ;
        RECT 627.540 13.950 627.800 14.270 ;
        RECT 621.160 2.000 621.300 13.950 ;
        RECT 620.950 -4.000 621.510 2.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 884.725 865.725 884.895 896.835 ;
        RECT 885.645 793.645 885.815 841.755 ;
        RECT 885.645 697.425 885.815 745.195 ;
        RECT 885.645 648.805 885.815 696.915 ;
        RECT 885.185 462.485 885.355 510.595 ;
        RECT 885.185 289.425 885.355 317.475 ;
      LAYER mcon ;
        RECT 884.725 896.665 884.895 896.835 ;
        RECT 885.645 841.585 885.815 841.755 ;
        RECT 885.645 745.025 885.815 745.195 ;
        RECT 885.645 696.745 885.815 696.915 ;
        RECT 885.185 510.425 885.355 510.595 ;
        RECT 885.185 317.305 885.355 317.475 ;
      LAYER met1 ;
        RECT 886.490 1062.740 886.810 1062.800 ;
        RECT 889.710 1062.740 890.030 1062.800 ;
        RECT 886.490 1062.600 890.030 1062.740 ;
        RECT 886.490 1062.540 886.810 1062.600 ;
        RECT 889.710 1062.540 890.030 1062.600 ;
        RECT 884.665 896.820 884.955 896.865 ;
        RECT 885.570 896.820 885.890 896.880 ;
        RECT 884.665 896.680 885.890 896.820 ;
        RECT 884.665 896.635 884.955 896.680 ;
        RECT 885.570 896.620 885.890 896.680 ;
        RECT 884.665 865.880 884.955 865.925 ;
        RECT 885.570 865.880 885.890 865.940 ;
        RECT 884.665 865.740 885.890 865.880 ;
        RECT 884.665 865.695 884.955 865.740 ;
        RECT 885.570 865.680 885.890 865.740 ;
        RECT 885.570 841.740 885.890 841.800 ;
        RECT 885.375 841.600 885.890 841.740 ;
        RECT 885.570 841.540 885.890 841.600 ;
        RECT 885.570 793.800 885.890 793.860 ;
        RECT 885.375 793.660 885.890 793.800 ;
        RECT 885.570 793.600 885.890 793.660 ;
        RECT 885.570 745.180 885.890 745.240 ;
        RECT 885.375 745.040 885.890 745.180 ;
        RECT 885.570 744.980 885.890 745.040 ;
        RECT 885.570 697.580 885.890 697.640 ;
        RECT 885.375 697.440 885.890 697.580 ;
        RECT 885.570 697.380 885.890 697.440 ;
        RECT 885.570 696.900 885.890 696.960 ;
        RECT 885.375 696.760 885.890 696.900 ;
        RECT 885.570 696.700 885.890 696.760 ;
        RECT 885.570 648.960 885.890 649.020 ;
        RECT 885.375 648.820 885.890 648.960 ;
        RECT 885.570 648.760 885.890 648.820 ;
        RECT 884.650 552.400 884.970 552.460 ;
        RECT 885.570 552.400 885.890 552.460 ;
        RECT 884.650 552.260 885.890 552.400 ;
        RECT 884.650 552.200 884.970 552.260 ;
        RECT 885.570 552.200 885.890 552.260 ;
        RECT 884.650 524.520 884.970 524.580 ;
        RECT 885.110 524.520 885.430 524.580 ;
        RECT 884.650 524.380 885.430 524.520 ;
        RECT 884.650 524.320 884.970 524.380 ;
        RECT 885.110 524.320 885.430 524.380 ;
        RECT 885.110 510.580 885.430 510.640 ;
        RECT 884.915 510.440 885.430 510.580 ;
        RECT 885.110 510.380 885.430 510.440 ;
        RECT 885.125 462.640 885.415 462.685 ;
        RECT 885.570 462.640 885.890 462.700 ;
        RECT 885.125 462.500 885.890 462.640 ;
        RECT 885.125 462.455 885.415 462.500 ;
        RECT 885.570 462.440 885.890 462.500 ;
        RECT 885.110 427.960 885.430 428.020 ;
        RECT 885.570 427.960 885.890 428.020 ;
        RECT 885.110 427.820 885.890 427.960 ;
        RECT 885.110 427.760 885.430 427.820 ;
        RECT 885.570 427.760 885.890 427.820 ;
        RECT 885.110 317.460 885.430 317.520 ;
        RECT 884.915 317.320 885.430 317.460 ;
        RECT 885.110 317.260 885.430 317.320 ;
        RECT 885.125 289.580 885.415 289.625 ;
        RECT 885.570 289.580 885.890 289.640 ;
        RECT 885.125 289.440 885.890 289.580 ;
        RECT 885.125 289.395 885.415 289.440 ;
        RECT 885.570 289.380 885.890 289.440 ;
        RECT 885.570 83.540 885.890 83.600 ;
        RECT 885.200 83.400 885.890 83.540 ;
        RECT 885.200 83.260 885.340 83.400 ;
        RECT 885.570 83.340 885.890 83.400 ;
        RECT 885.110 83.000 885.430 83.260 ;
        RECT 115.530 45.460 115.850 45.520 ;
        RECT 885.110 45.460 885.430 45.520 ;
        RECT 115.530 45.320 885.430 45.460 ;
        RECT 115.530 45.260 115.850 45.320 ;
        RECT 885.110 45.260 885.430 45.320 ;
      LAYER via ;
        RECT 886.520 1062.540 886.780 1062.800 ;
        RECT 889.740 1062.540 890.000 1062.800 ;
        RECT 885.600 896.620 885.860 896.880 ;
        RECT 885.600 865.680 885.860 865.940 ;
        RECT 885.600 841.540 885.860 841.800 ;
        RECT 885.600 793.600 885.860 793.860 ;
        RECT 885.600 744.980 885.860 745.240 ;
        RECT 885.600 697.380 885.860 697.640 ;
        RECT 885.600 696.700 885.860 696.960 ;
        RECT 885.600 648.760 885.860 649.020 ;
        RECT 884.680 552.200 884.940 552.460 ;
        RECT 885.600 552.200 885.860 552.460 ;
        RECT 884.680 524.320 884.940 524.580 ;
        RECT 885.140 524.320 885.400 524.580 ;
        RECT 885.140 510.380 885.400 510.640 ;
        RECT 885.600 462.440 885.860 462.700 ;
        RECT 885.140 427.760 885.400 428.020 ;
        RECT 885.600 427.760 885.860 428.020 ;
        RECT 885.140 317.260 885.400 317.520 ;
        RECT 885.600 289.380 885.860 289.640 ;
        RECT 885.600 83.340 885.860 83.600 ;
        RECT 885.140 83.000 885.400 83.260 ;
        RECT 115.560 45.260 115.820 45.520 ;
        RECT 885.140 45.260 885.400 45.520 ;
      LAYER met2 ;
        RECT 889.650 1100.580 889.930 1104.000 ;
        RECT 889.650 1100.000 889.940 1100.580 ;
        RECT 889.800 1062.830 889.940 1100.000 ;
        RECT 886.520 1062.510 886.780 1062.830 ;
        RECT 889.740 1062.510 890.000 1062.830 ;
        RECT 886.580 976.210 886.720 1062.510 ;
        RECT 885.660 976.070 886.720 976.210 ;
        RECT 885.660 896.910 885.800 976.070 ;
        RECT 885.600 896.590 885.860 896.910 ;
        RECT 885.600 865.650 885.860 865.970 ;
        RECT 885.660 841.830 885.800 865.650 ;
        RECT 885.600 841.510 885.860 841.830 ;
        RECT 885.600 793.570 885.860 793.890 ;
        RECT 885.660 745.270 885.800 793.570 ;
        RECT 885.600 744.950 885.860 745.270 ;
        RECT 885.600 697.350 885.860 697.670 ;
        RECT 885.660 696.990 885.800 697.350 ;
        RECT 885.600 696.670 885.860 696.990 ;
        RECT 885.600 648.730 885.860 649.050 ;
        RECT 885.660 552.490 885.800 648.730 ;
        RECT 884.680 552.170 884.940 552.490 ;
        RECT 885.600 552.170 885.860 552.490 ;
        RECT 884.740 524.610 884.880 552.170 ;
        RECT 884.680 524.290 884.940 524.610 ;
        RECT 885.140 524.290 885.400 524.610 ;
        RECT 885.200 510.670 885.340 524.290 ;
        RECT 885.140 510.350 885.400 510.670 ;
        RECT 885.600 462.410 885.860 462.730 ;
        RECT 885.660 428.050 885.800 462.410 ;
        RECT 885.140 427.730 885.400 428.050 ;
        RECT 885.600 427.730 885.860 428.050 ;
        RECT 885.200 317.550 885.340 427.730 ;
        RECT 885.140 317.230 885.400 317.550 ;
        RECT 885.600 289.350 885.860 289.670 ;
        RECT 885.660 179.930 885.800 289.350 ;
        RECT 885.200 179.790 885.800 179.930 ;
        RECT 885.200 155.450 885.340 179.790 ;
        RECT 885.200 155.310 885.800 155.450 ;
        RECT 885.660 83.630 885.800 155.310 ;
        RECT 885.600 83.310 885.860 83.630 ;
        RECT 885.140 82.970 885.400 83.290 ;
        RECT 885.200 45.550 885.340 82.970 ;
        RECT 115.560 45.230 115.820 45.550 ;
        RECT 885.140 45.230 885.400 45.550 ;
        RECT 115.620 2.000 115.760 45.230 ;
        RECT 115.410 -4.000 115.970 2.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 144.510 51.580 144.830 51.640 ;
        RECT 897.990 51.580 898.310 51.640 ;
        RECT 144.510 51.440 898.310 51.580 ;
        RECT 144.510 51.380 144.830 51.440 ;
        RECT 897.990 51.380 898.310 51.440 ;
        RECT 139.450 16.900 139.770 16.960 ;
        RECT 144.510 16.900 144.830 16.960 ;
        RECT 139.450 16.760 144.830 16.900 ;
        RECT 139.450 16.700 139.770 16.760 ;
        RECT 144.510 16.700 144.830 16.760 ;
      LAYER via ;
        RECT 144.540 51.380 144.800 51.640 ;
        RECT 898.020 51.380 898.280 51.640 ;
        RECT 139.480 16.700 139.740 16.960 ;
        RECT 144.540 16.700 144.800 16.960 ;
      LAYER met2 ;
        RECT 897.930 1100.580 898.210 1104.000 ;
        RECT 897.930 1100.000 898.220 1100.580 ;
        RECT 898.080 51.670 898.220 1100.000 ;
        RECT 144.540 51.350 144.800 51.670 ;
        RECT 898.020 51.350 898.280 51.670 ;
        RECT 144.600 16.990 144.740 51.350 ;
        RECT 139.480 16.670 139.740 16.990 ;
        RECT 144.540 16.670 144.800 16.990 ;
        RECT 139.540 2.000 139.680 16.670 ;
        RECT 139.330 -4.000 139.890 2.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 158.310 58.720 158.630 58.780 ;
        RECT 904.890 58.720 905.210 58.780 ;
        RECT 158.310 58.580 905.210 58.720 ;
        RECT 158.310 58.520 158.630 58.580 ;
        RECT 904.890 58.520 905.210 58.580 ;
      LAYER via ;
        RECT 158.340 58.520 158.600 58.780 ;
        RECT 904.920 58.520 905.180 58.780 ;
      LAYER met2 ;
        RECT 903.910 1100.650 904.190 1104.000 ;
        RECT 903.910 1100.510 905.120 1100.650 ;
        RECT 903.910 1100.000 904.190 1100.510 ;
        RECT 904.980 58.810 905.120 1100.510 ;
        RECT 158.340 58.490 158.600 58.810 ;
        RECT 904.920 58.490 905.180 58.810 ;
        RECT 158.400 16.730 158.540 58.490 ;
        RECT 157.480 16.590 158.540 16.730 ;
        RECT 157.480 2.000 157.620 16.590 ;
        RECT 157.270 -4.000 157.830 2.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 905.425 848.725 905.595 896.835 ;
        RECT 905.425 758.965 905.595 807.075 ;
        RECT 905.425 662.745 905.595 710.515 ;
        RECT 905.425 614.125 905.595 662.235 ;
        RECT 904.965 559.385 905.135 607.155 ;
        RECT 905.885 606.985 906.055 613.615 ;
        RECT 905.425 511.105 905.595 558.875 ;
        RECT 906.345 324.445 906.515 372.555 ;
        RECT 905.425 269.025 905.595 293.335 ;
        RECT 905.425 131.325 905.595 220.575 ;
      LAYER mcon ;
        RECT 905.425 896.665 905.595 896.835 ;
        RECT 905.425 806.905 905.595 807.075 ;
        RECT 905.425 710.345 905.595 710.515 ;
        RECT 905.425 662.065 905.595 662.235 ;
        RECT 905.885 613.445 906.055 613.615 ;
        RECT 904.965 606.985 905.135 607.155 ;
        RECT 905.425 558.705 905.595 558.875 ;
        RECT 906.345 372.385 906.515 372.555 ;
        RECT 905.425 293.165 905.595 293.335 ;
        RECT 905.425 220.405 905.595 220.575 ;
      LAYER met1 ;
        RECT 906.730 1087.900 907.050 1087.960 ;
        RECT 909.490 1087.900 909.810 1087.960 ;
        RECT 906.730 1087.760 909.810 1087.900 ;
        RECT 906.730 1087.700 907.050 1087.760 ;
        RECT 909.490 1087.700 909.810 1087.760 ;
        RECT 905.810 931.840 906.130 931.900 ;
        RECT 905.440 931.700 906.130 931.840 ;
        RECT 905.440 931.560 905.580 931.700 ;
        RECT 905.810 931.640 906.130 931.700 ;
        RECT 905.350 931.300 905.670 931.560 ;
        RECT 905.350 896.820 905.670 896.880 ;
        RECT 905.155 896.680 905.670 896.820 ;
        RECT 905.350 896.620 905.670 896.680 ;
        RECT 905.365 848.880 905.655 848.925 ;
        RECT 906.730 848.880 907.050 848.940 ;
        RECT 905.365 848.740 907.050 848.880 ;
        RECT 905.365 848.695 905.655 848.740 ;
        RECT 906.730 848.680 907.050 848.740 ;
        RECT 905.350 807.060 905.670 807.120 ;
        RECT 905.155 806.920 905.670 807.060 ;
        RECT 905.350 806.860 905.670 806.920 ;
        RECT 905.350 759.120 905.670 759.180 ;
        RECT 905.155 758.980 905.670 759.120 ;
        RECT 905.350 758.920 905.670 758.980 ;
        RECT 905.350 710.500 905.670 710.560 ;
        RECT 905.155 710.360 905.670 710.500 ;
        RECT 905.350 710.300 905.670 710.360 ;
        RECT 905.365 662.900 905.655 662.945 ;
        RECT 905.810 662.900 906.130 662.960 ;
        RECT 905.365 662.760 906.130 662.900 ;
        RECT 905.365 662.715 905.655 662.760 ;
        RECT 905.810 662.700 906.130 662.760 ;
        RECT 905.365 662.220 905.655 662.265 ;
        RECT 905.810 662.220 906.130 662.280 ;
        RECT 905.365 662.080 906.130 662.220 ;
        RECT 905.365 662.035 905.655 662.080 ;
        RECT 905.810 662.020 906.130 662.080 ;
        RECT 905.350 614.280 905.670 614.340 ;
        RECT 905.155 614.140 905.670 614.280 ;
        RECT 905.350 614.080 905.670 614.140 ;
        RECT 905.350 613.600 905.670 613.660 ;
        RECT 905.825 613.600 906.115 613.645 ;
        RECT 905.350 613.460 906.115 613.600 ;
        RECT 905.350 613.400 905.670 613.460 ;
        RECT 905.825 613.415 906.115 613.460 ;
        RECT 904.905 607.140 905.195 607.185 ;
        RECT 905.825 607.140 906.115 607.185 ;
        RECT 904.905 607.000 906.115 607.140 ;
        RECT 904.905 606.955 905.195 607.000 ;
        RECT 905.825 606.955 906.115 607.000 ;
        RECT 904.905 559.540 905.195 559.585 ;
        RECT 905.350 559.540 905.670 559.600 ;
        RECT 904.905 559.400 905.670 559.540 ;
        RECT 904.905 559.355 905.195 559.400 ;
        RECT 905.350 559.340 905.670 559.400 ;
        RECT 905.350 558.860 905.670 558.920 ;
        RECT 905.155 558.720 905.670 558.860 ;
        RECT 905.350 558.660 905.670 558.720 ;
        RECT 905.350 511.260 905.670 511.320 ;
        RECT 905.155 511.120 905.670 511.260 ;
        RECT 905.350 511.060 905.670 511.120 ;
        RECT 905.350 510.580 905.670 510.640 ;
        RECT 907.190 510.580 907.510 510.640 ;
        RECT 905.350 510.440 907.510 510.580 ;
        RECT 905.350 510.380 905.670 510.440 ;
        RECT 907.190 510.380 907.510 510.440 ;
        RECT 906.270 372.540 906.590 372.600 ;
        RECT 906.075 372.400 906.590 372.540 ;
        RECT 906.270 372.340 906.590 372.400 ;
        RECT 905.350 324.600 905.670 324.660 ;
        RECT 906.285 324.600 906.575 324.645 ;
        RECT 905.350 324.460 906.575 324.600 ;
        RECT 905.350 324.400 905.670 324.460 ;
        RECT 906.285 324.415 906.575 324.460 ;
        RECT 905.350 293.320 905.670 293.380 ;
        RECT 905.155 293.180 905.670 293.320 ;
        RECT 905.350 293.120 905.670 293.180 ;
        RECT 905.365 269.180 905.655 269.225 ;
        RECT 905.810 269.180 906.130 269.240 ;
        RECT 905.365 269.040 906.130 269.180 ;
        RECT 905.365 268.995 905.655 269.040 ;
        RECT 905.810 268.980 906.130 269.040 ;
        RECT 905.810 228.380 906.130 228.440 ;
        RECT 905.440 228.240 906.130 228.380 ;
        RECT 905.440 228.100 905.580 228.240 ;
        RECT 905.810 228.180 906.130 228.240 ;
        RECT 905.350 227.840 905.670 228.100 ;
        RECT 905.365 220.560 905.655 220.605 ;
        RECT 906.730 220.560 907.050 220.620 ;
        RECT 905.365 220.420 907.050 220.560 ;
        RECT 905.365 220.375 905.655 220.420 ;
        RECT 906.730 220.360 907.050 220.420 ;
        RECT 905.350 131.480 905.670 131.540 ;
        RECT 905.155 131.340 905.670 131.480 ;
        RECT 905.350 131.280 905.670 131.340 ;
        RECT 905.810 130.800 906.130 130.860 ;
        RECT 906.730 130.800 907.050 130.860 ;
        RECT 905.810 130.660 907.050 130.800 ;
        RECT 905.810 130.600 906.130 130.660 ;
        RECT 906.730 130.600 907.050 130.660 ;
        RECT 905.350 41.720 905.670 41.780 ;
        RECT 906.270 41.720 906.590 41.780 ;
        RECT 905.350 41.580 906.590 41.720 ;
        RECT 905.350 41.520 905.670 41.580 ;
        RECT 906.270 41.520 906.590 41.580 ;
        RECT 174.870 18.940 175.190 19.000 ;
        RECT 905.350 18.940 905.670 19.000 ;
        RECT 174.870 18.800 905.670 18.940 ;
        RECT 174.870 18.740 175.190 18.800 ;
        RECT 905.350 18.740 905.670 18.800 ;
      LAYER via ;
        RECT 906.760 1087.700 907.020 1087.960 ;
        RECT 909.520 1087.700 909.780 1087.960 ;
        RECT 905.840 931.640 906.100 931.900 ;
        RECT 905.380 931.300 905.640 931.560 ;
        RECT 905.380 896.620 905.640 896.880 ;
        RECT 906.760 848.680 907.020 848.940 ;
        RECT 905.380 806.860 905.640 807.120 ;
        RECT 905.380 758.920 905.640 759.180 ;
        RECT 905.380 710.300 905.640 710.560 ;
        RECT 905.840 662.700 906.100 662.960 ;
        RECT 905.840 662.020 906.100 662.280 ;
        RECT 905.380 614.080 905.640 614.340 ;
        RECT 905.380 613.400 905.640 613.660 ;
        RECT 905.380 559.340 905.640 559.600 ;
        RECT 905.380 558.660 905.640 558.920 ;
        RECT 905.380 511.060 905.640 511.320 ;
        RECT 905.380 510.380 905.640 510.640 ;
        RECT 907.220 510.380 907.480 510.640 ;
        RECT 906.300 372.340 906.560 372.600 ;
        RECT 905.380 324.400 905.640 324.660 ;
        RECT 905.380 293.120 905.640 293.380 ;
        RECT 905.840 268.980 906.100 269.240 ;
        RECT 905.840 228.180 906.100 228.440 ;
        RECT 905.380 227.840 905.640 228.100 ;
        RECT 906.760 220.360 907.020 220.620 ;
        RECT 905.380 131.280 905.640 131.540 ;
        RECT 905.840 130.600 906.100 130.860 ;
        RECT 906.760 130.600 907.020 130.860 ;
        RECT 905.380 41.520 905.640 41.780 ;
        RECT 906.300 41.520 906.560 41.780 ;
        RECT 174.900 18.740 175.160 19.000 ;
        RECT 905.380 18.740 905.640 19.000 ;
      LAYER met2 ;
        RECT 909.890 1100.650 910.170 1104.000 ;
        RECT 909.580 1100.510 910.170 1100.650 ;
        RECT 909.580 1087.990 909.720 1100.510 ;
        RECT 909.890 1100.000 910.170 1100.510 ;
        RECT 906.760 1087.670 907.020 1087.990 ;
        RECT 909.520 1087.670 909.780 1087.990 ;
        RECT 906.820 1051.690 906.960 1087.670 ;
        RECT 905.900 1051.550 906.960 1051.690 ;
        RECT 905.900 931.930 906.040 1051.550 ;
        RECT 905.840 931.610 906.100 931.930 ;
        RECT 905.380 931.270 905.640 931.590 ;
        RECT 905.440 896.910 905.580 931.270 ;
        RECT 905.380 896.590 905.640 896.910 ;
        RECT 906.760 848.650 907.020 848.970 ;
        RECT 906.820 830.690 906.960 848.650 ;
        RECT 905.440 830.550 906.960 830.690 ;
        RECT 905.440 807.150 905.580 830.550 ;
        RECT 905.380 806.830 905.640 807.150 ;
        RECT 905.380 758.890 905.640 759.210 ;
        RECT 905.440 710.590 905.580 758.890 ;
        RECT 905.380 710.270 905.640 710.590 ;
        RECT 905.840 662.670 906.100 662.990 ;
        RECT 905.900 662.310 906.040 662.670 ;
        RECT 905.840 661.990 906.100 662.310 ;
        RECT 905.380 614.050 905.640 614.370 ;
        RECT 905.440 613.690 905.580 614.050 ;
        RECT 905.380 613.370 905.640 613.690 ;
        RECT 905.380 559.310 905.640 559.630 ;
        RECT 905.440 558.950 905.580 559.310 ;
        RECT 905.380 558.630 905.640 558.950 ;
        RECT 905.380 511.030 905.640 511.350 ;
        RECT 905.440 510.670 905.580 511.030 ;
        RECT 905.380 510.350 905.640 510.670 ;
        RECT 907.220 510.350 907.480 510.670 ;
        RECT 907.280 427.450 907.420 510.350 ;
        RECT 906.820 427.310 907.420 427.450 ;
        RECT 906.820 420.650 906.960 427.310 ;
        RECT 906.820 420.510 907.420 420.650 ;
        RECT 907.280 379.680 907.420 420.510 ;
        RECT 906.360 379.540 907.420 379.680 ;
        RECT 906.360 372.630 906.500 379.540 ;
        RECT 906.300 372.310 906.560 372.630 ;
        RECT 905.380 324.370 905.640 324.690 ;
        RECT 905.440 293.410 905.580 324.370 ;
        RECT 905.380 293.090 905.640 293.410 ;
        RECT 905.840 268.950 906.100 269.270 ;
        RECT 905.900 228.470 906.040 268.950 ;
        RECT 905.840 228.150 906.100 228.470 ;
        RECT 905.380 227.810 905.640 228.130 ;
        RECT 905.440 227.530 905.580 227.810 ;
        RECT 905.440 227.390 906.960 227.530 ;
        RECT 906.820 220.650 906.960 227.390 ;
        RECT 906.760 220.330 907.020 220.650 ;
        RECT 905.380 131.250 905.640 131.570 ;
        RECT 905.440 130.970 905.580 131.250 ;
        RECT 905.440 130.890 906.040 130.970 ;
        RECT 905.440 130.830 906.100 130.890 ;
        RECT 905.840 130.570 906.100 130.830 ;
        RECT 906.760 130.570 907.020 130.890 ;
        RECT 906.820 89.490 906.960 130.570 ;
        RECT 906.360 89.350 906.960 89.490 ;
        RECT 906.360 41.810 906.500 89.350 ;
        RECT 905.380 41.490 905.640 41.810 ;
        RECT 906.300 41.490 906.560 41.810 ;
        RECT 905.440 19.030 905.580 41.490 ;
        RECT 174.900 18.710 175.160 19.030 ;
        RECT 905.380 18.710 905.640 19.030 ;
        RECT 174.960 2.000 175.100 18.710 ;
        RECT 174.750 -4.000 175.310 2.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 854.365 1087.405 854.535 1088.595 ;
        RECT 339.625 15.045 339.795 16.575 ;
        RECT 347.905 16.405 348.995 16.575 ;
        RECT 347.905 15.045 348.075 16.405 ;
        RECT 348.825 16.065 348.995 16.405 ;
      LAYER mcon ;
        RECT 854.365 1088.425 854.535 1088.595 ;
        RECT 339.625 16.405 339.795 16.575 ;
      LAYER met1 ;
        RECT 355.190 1088.580 355.510 1088.640 ;
        RECT 854.305 1088.580 854.595 1088.625 ;
        RECT 355.190 1088.440 854.595 1088.580 ;
        RECT 355.190 1088.380 355.510 1088.440 ;
        RECT 854.305 1088.395 854.595 1088.440 ;
        RECT 854.305 1087.560 854.595 1087.605 ;
        RECT 915.930 1087.560 916.250 1087.620 ;
        RECT 854.305 1087.420 916.250 1087.560 ;
        RECT 854.305 1087.375 854.595 1087.420 ;
        RECT 915.930 1087.360 916.250 1087.420 ;
        RECT 192.810 16.560 193.130 16.620 ;
        RECT 339.565 16.560 339.855 16.605 ;
        RECT 192.810 16.420 339.855 16.560 ;
        RECT 192.810 16.360 193.130 16.420 ;
        RECT 339.565 16.375 339.855 16.420 ;
        RECT 348.765 16.220 349.055 16.265 ;
        RECT 355.190 16.220 355.510 16.280 ;
        RECT 348.765 16.080 355.510 16.220 ;
        RECT 348.765 16.035 349.055 16.080 ;
        RECT 355.190 16.020 355.510 16.080 ;
        RECT 339.565 15.200 339.855 15.245 ;
        RECT 347.845 15.200 348.135 15.245 ;
        RECT 339.565 15.060 348.135 15.200 ;
        RECT 339.565 15.015 339.855 15.060 ;
        RECT 347.845 15.015 348.135 15.060 ;
      LAYER via ;
        RECT 355.220 1088.380 355.480 1088.640 ;
        RECT 915.960 1087.360 916.220 1087.620 ;
        RECT 192.840 16.360 193.100 16.620 ;
        RECT 355.220 16.020 355.480 16.280 ;
      LAYER met2 ;
        RECT 915.870 1100.580 916.150 1104.000 ;
        RECT 915.870 1100.000 916.160 1100.580 ;
        RECT 355.220 1088.350 355.480 1088.670 ;
        RECT 192.840 16.330 193.100 16.650 ;
        RECT 192.900 2.000 193.040 16.330 ;
        RECT 355.280 16.310 355.420 1088.350 ;
        RECT 916.020 1087.650 916.160 1100.000 ;
        RECT 915.960 1087.330 916.220 1087.650 ;
        RECT 355.220 15.990 355.480 16.310 ;
        RECT 192.690 -4.000 193.250 2.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 920.145 544.085 920.315 579.615 ;
        RECT 920.145 331.245 920.315 379.355 ;
        RECT 919.685 227.885 919.855 275.995 ;
      LAYER mcon ;
        RECT 920.145 579.445 920.315 579.615 ;
        RECT 920.145 379.185 920.315 379.355 ;
        RECT 919.685 275.825 919.855 275.995 ;
      LAYER met1 ;
        RECT 920.070 1062.740 920.390 1062.800 ;
        RECT 922.370 1062.740 922.690 1062.800 ;
        RECT 920.070 1062.600 922.690 1062.740 ;
        RECT 920.070 1062.540 920.390 1062.600 ;
        RECT 922.370 1062.540 922.690 1062.600 ;
        RECT 920.530 1007.320 920.850 1007.380 ;
        RECT 921.450 1007.320 921.770 1007.380 ;
        RECT 920.530 1007.180 921.770 1007.320 ;
        RECT 920.530 1007.120 920.850 1007.180 ;
        RECT 921.450 1007.120 921.770 1007.180 ;
        RECT 920.070 918.240 920.390 918.300 ;
        RECT 920.530 918.240 920.850 918.300 ;
        RECT 920.070 918.100 920.850 918.240 ;
        RECT 920.070 918.040 920.390 918.100 ;
        RECT 920.530 918.040 920.850 918.100 ;
        RECT 920.530 910.760 920.850 910.820 ;
        RECT 920.990 910.760 921.310 910.820 ;
        RECT 920.530 910.620 921.310 910.760 ;
        RECT 920.530 910.560 920.850 910.620 ;
        RECT 920.990 910.560 921.310 910.620 ;
        RECT 920.070 821.000 920.390 821.060 ;
        RECT 920.530 821.000 920.850 821.060 ;
        RECT 920.070 820.860 920.850 821.000 ;
        RECT 920.070 820.800 920.390 820.860 ;
        RECT 920.530 820.800 920.850 820.860 ;
        RECT 920.070 738.520 920.390 738.780 ;
        RECT 920.160 738.100 920.300 738.520 ;
        RECT 920.070 737.840 920.390 738.100 ;
        RECT 919.610 676.160 919.930 676.220 ;
        RECT 920.070 676.160 920.390 676.220 ;
        RECT 919.610 676.020 920.390 676.160 ;
        RECT 919.610 675.960 919.930 676.020 ;
        RECT 920.070 675.960 920.390 676.020 ;
        RECT 919.610 627.880 919.930 627.940 ;
        RECT 920.530 627.880 920.850 627.940 ;
        RECT 919.610 627.740 920.850 627.880 ;
        RECT 919.610 627.680 919.930 627.740 ;
        RECT 920.530 627.680 920.850 627.740 ;
        RECT 920.070 579.600 920.390 579.660 ;
        RECT 919.875 579.460 920.390 579.600 ;
        RECT 920.070 579.400 920.390 579.460 ;
        RECT 920.085 544.240 920.375 544.285 ;
        RECT 920.530 544.240 920.850 544.300 ;
        RECT 920.085 544.100 920.850 544.240 ;
        RECT 920.085 544.055 920.375 544.100 ;
        RECT 920.530 544.040 920.850 544.100 ;
        RECT 920.070 379.340 920.390 379.400 ;
        RECT 919.875 379.200 920.390 379.340 ;
        RECT 920.070 379.140 920.390 379.200 ;
        RECT 920.085 331.400 920.375 331.445 ;
        RECT 920.530 331.400 920.850 331.460 ;
        RECT 920.085 331.260 920.850 331.400 ;
        RECT 920.085 331.215 920.375 331.260 ;
        RECT 920.530 331.200 920.850 331.260 ;
        RECT 919.610 289.580 919.930 289.640 ;
        RECT 920.530 289.580 920.850 289.640 ;
        RECT 919.610 289.440 920.850 289.580 ;
        RECT 919.610 289.380 919.930 289.440 ;
        RECT 920.530 289.380 920.850 289.440 ;
        RECT 919.610 275.980 919.930 276.040 ;
        RECT 919.415 275.840 919.930 275.980 ;
        RECT 919.610 275.780 919.930 275.840 ;
        RECT 919.610 228.040 919.930 228.100 ;
        RECT 919.415 227.900 919.930 228.040 ;
        RECT 919.610 227.840 919.930 227.900 ;
        RECT 920.070 144.740 920.390 144.800 ;
        RECT 920.530 144.740 920.850 144.800 ;
        RECT 920.070 144.600 920.850 144.740 ;
        RECT 920.070 144.540 920.390 144.600 ;
        RECT 920.530 144.540 920.850 144.600 ;
        RECT 210.750 19.620 211.070 19.680 ;
        RECT 919.610 19.620 919.930 19.680 ;
        RECT 210.750 19.480 919.930 19.620 ;
        RECT 210.750 19.420 211.070 19.480 ;
        RECT 919.610 19.420 919.930 19.480 ;
      LAYER via ;
        RECT 920.100 1062.540 920.360 1062.800 ;
        RECT 922.400 1062.540 922.660 1062.800 ;
        RECT 920.560 1007.120 920.820 1007.380 ;
        RECT 921.480 1007.120 921.740 1007.380 ;
        RECT 920.100 918.040 920.360 918.300 ;
        RECT 920.560 918.040 920.820 918.300 ;
        RECT 920.560 910.560 920.820 910.820 ;
        RECT 921.020 910.560 921.280 910.820 ;
        RECT 920.100 820.800 920.360 821.060 ;
        RECT 920.560 820.800 920.820 821.060 ;
        RECT 920.100 738.520 920.360 738.780 ;
        RECT 920.100 737.840 920.360 738.100 ;
        RECT 919.640 675.960 919.900 676.220 ;
        RECT 920.100 675.960 920.360 676.220 ;
        RECT 919.640 627.680 919.900 627.940 ;
        RECT 920.560 627.680 920.820 627.940 ;
        RECT 920.100 579.400 920.360 579.660 ;
        RECT 920.560 544.040 920.820 544.300 ;
        RECT 920.100 379.140 920.360 379.400 ;
        RECT 920.560 331.200 920.820 331.460 ;
        RECT 919.640 289.380 919.900 289.640 ;
        RECT 920.560 289.380 920.820 289.640 ;
        RECT 919.640 275.780 919.900 276.040 ;
        RECT 919.640 227.840 919.900 228.100 ;
        RECT 920.100 144.540 920.360 144.800 ;
        RECT 920.560 144.540 920.820 144.800 ;
        RECT 210.780 19.420 211.040 19.680 ;
        RECT 919.640 19.420 919.900 19.680 ;
      LAYER met2 ;
        RECT 922.310 1100.580 922.590 1104.000 ;
        RECT 922.310 1100.000 922.600 1100.580 ;
        RECT 922.460 1062.830 922.600 1100.000 ;
        RECT 920.100 1062.510 920.360 1062.830 ;
        RECT 922.400 1062.510 922.660 1062.830 ;
        RECT 920.160 1027.890 920.300 1062.510 ;
        RECT 920.160 1027.750 920.760 1027.890 ;
        RECT 920.620 1007.410 920.760 1027.750 ;
        RECT 920.560 1007.090 920.820 1007.410 ;
        RECT 921.480 1007.090 921.740 1007.410 ;
        RECT 921.540 959.325 921.680 1007.090 ;
        RECT 920.090 958.955 920.370 959.325 ;
        RECT 921.470 958.955 921.750 959.325 ;
        RECT 920.160 918.330 920.300 958.955 ;
        RECT 920.100 918.010 920.360 918.330 ;
        RECT 920.560 918.010 920.820 918.330 ;
        RECT 920.620 910.850 920.760 918.010 ;
        RECT 920.560 910.530 920.820 910.850 ;
        RECT 921.020 910.530 921.280 910.850 ;
        RECT 921.080 845.650 921.220 910.530 ;
        RECT 920.620 845.510 921.220 845.650 ;
        RECT 920.620 821.090 920.760 845.510 ;
        RECT 920.100 820.770 920.360 821.090 ;
        RECT 920.560 820.770 920.820 821.090 ;
        RECT 920.160 738.810 920.300 820.770 ;
        RECT 920.100 738.490 920.360 738.810 ;
        RECT 920.100 737.810 920.360 738.130 ;
        RECT 920.160 676.250 920.300 737.810 ;
        RECT 919.640 675.930 919.900 676.250 ;
        RECT 920.100 675.930 920.360 676.250 ;
        RECT 919.700 641.650 919.840 675.930 ;
        RECT 919.700 641.510 920.300 641.650 ;
        RECT 920.160 628.050 920.300 641.510 ;
        RECT 920.160 627.970 920.760 628.050 ;
        RECT 919.640 627.650 919.900 627.970 ;
        RECT 920.160 627.910 920.820 627.970 ;
        RECT 920.560 627.650 920.820 627.910 ;
        RECT 919.700 593.370 919.840 627.650 ;
        RECT 919.700 593.230 920.300 593.370 ;
        RECT 920.160 579.690 920.300 593.230 ;
        RECT 920.100 579.370 920.360 579.690 ;
        RECT 920.560 544.010 920.820 544.330 ;
        RECT 920.620 497.490 920.760 544.010 ;
        RECT 920.620 497.350 921.220 497.490 ;
        RECT 921.080 496.810 921.220 497.350 ;
        RECT 920.620 496.670 921.220 496.810 ;
        RECT 920.620 379.850 920.760 496.670 ;
        RECT 920.160 379.710 920.760 379.850 ;
        RECT 920.160 379.430 920.300 379.710 ;
        RECT 920.100 379.110 920.360 379.430 ;
        RECT 920.560 331.170 920.820 331.490 ;
        RECT 920.620 289.670 920.760 331.170 ;
        RECT 919.640 289.350 919.900 289.670 ;
        RECT 920.560 289.350 920.820 289.670 ;
        RECT 919.700 276.070 919.840 289.350 ;
        RECT 919.640 275.750 919.900 276.070 ;
        RECT 919.640 227.810 919.900 228.130 ;
        RECT 919.700 193.530 919.840 227.810 ;
        RECT 919.700 193.390 920.300 193.530 ;
        RECT 920.160 169.050 920.300 193.390 ;
        RECT 920.160 168.910 921.220 169.050 ;
        RECT 921.080 158.170 921.220 168.910 ;
        RECT 920.620 158.030 921.220 158.170 ;
        RECT 920.620 144.830 920.760 158.030 ;
        RECT 920.100 144.510 920.360 144.830 ;
        RECT 920.560 144.510 920.820 144.830 ;
        RECT 920.160 48.010 920.300 144.510 ;
        RECT 919.700 47.870 920.300 48.010 ;
        RECT 919.700 19.710 919.840 47.870 ;
        RECT 210.780 19.390 211.040 19.710 ;
        RECT 919.640 19.390 919.900 19.710 ;
        RECT 210.840 2.000 210.980 19.390 ;
        RECT 210.630 -4.000 211.190 2.000 ;
      LAYER via2 ;
        RECT 920.090 959.000 920.370 959.280 ;
        RECT 921.470 959.000 921.750 959.280 ;
      LAYER met3 ;
        RECT 920.065 959.290 920.395 959.305 ;
        RECT 921.445 959.290 921.775 959.305 ;
        RECT 920.065 958.990 921.775 959.290 ;
        RECT 920.065 958.975 920.395 958.990 ;
        RECT 921.445 958.975 921.775 958.990 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 348.365 14.025 348.535 16.235 ;
      LAYER mcon ;
        RECT 348.365 16.065 348.535 16.235 ;
      LAYER met1 ;
        RECT 375.890 1088.920 376.210 1088.980 ;
        RECT 928.350 1088.920 928.670 1088.980 ;
        RECT 375.890 1088.780 928.670 1088.920 ;
        RECT 375.890 1088.720 376.210 1088.780 ;
        RECT 928.350 1088.720 928.670 1088.780 ;
        RECT 228.690 16.220 229.010 16.280 ;
        RECT 348.305 16.220 348.595 16.265 ;
        RECT 228.690 16.080 348.595 16.220 ;
        RECT 228.690 16.020 229.010 16.080 ;
        RECT 348.305 16.035 348.595 16.080 ;
        RECT 348.305 14.180 348.595 14.225 ;
        RECT 375.890 14.180 376.210 14.240 ;
        RECT 348.305 14.040 376.210 14.180 ;
        RECT 348.305 13.995 348.595 14.040 ;
        RECT 375.890 13.980 376.210 14.040 ;
      LAYER via ;
        RECT 375.920 1088.720 376.180 1088.980 ;
        RECT 928.380 1088.720 928.640 1088.980 ;
        RECT 228.720 16.020 228.980 16.280 ;
        RECT 375.920 13.980 376.180 14.240 ;
      LAYER met2 ;
        RECT 928.290 1100.580 928.570 1104.000 ;
        RECT 928.290 1100.000 928.580 1100.580 ;
        RECT 928.440 1089.010 928.580 1100.000 ;
        RECT 375.920 1088.690 376.180 1089.010 ;
        RECT 928.380 1088.690 928.640 1089.010 ;
        RECT 228.720 15.990 228.980 16.310 ;
        RECT 228.780 2.000 228.920 15.990 ;
        RECT 375.980 14.270 376.120 1088.690 ;
        RECT 375.920 13.950 376.180 14.270 ;
        RECT 228.570 -4.000 229.130 2.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 50.210 17.240 50.530 17.300 ;
        RECT 864.410 17.240 864.730 17.300 ;
        RECT 50.210 17.100 864.730 17.240 ;
        RECT 50.210 17.040 50.530 17.100 ;
        RECT 864.410 17.040 864.730 17.100 ;
      LAYER via ;
        RECT 50.240 17.040 50.500 17.300 ;
        RECT 864.440 17.040 864.700 17.300 ;
      LAYER met2 ;
        RECT 867.110 1100.650 867.390 1104.000 ;
        RECT 865.880 1100.510 867.390 1100.650 ;
        RECT 865.880 1053.050 866.020 1100.510 ;
        RECT 867.110 1100.000 867.390 1100.510 ;
        RECT 864.500 1052.910 866.020 1053.050 ;
        RECT 864.500 17.330 864.640 1052.910 ;
        RECT 50.240 17.010 50.500 17.330 ;
        RECT 864.440 17.010 864.700 17.330 ;
        RECT 50.300 2.000 50.440 17.010 ;
        RECT 50.090 -4.000 50.650 2.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 389.690 1089.260 390.010 1089.320 ;
        RECT 936.630 1089.260 936.950 1089.320 ;
        RECT 389.690 1089.120 936.950 1089.260 ;
        RECT 389.690 1089.060 390.010 1089.120 ;
        RECT 936.630 1089.060 936.950 1089.120 ;
        RECT 252.610 15.540 252.930 15.600 ;
        RECT 389.690 15.540 390.010 15.600 ;
        RECT 252.610 15.400 390.010 15.540 ;
        RECT 252.610 15.340 252.930 15.400 ;
        RECT 389.690 15.340 390.010 15.400 ;
      LAYER via ;
        RECT 389.720 1089.060 389.980 1089.320 ;
        RECT 936.660 1089.060 936.920 1089.320 ;
        RECT 252.640 15.340 252.900 15.600 ;
        RECT 389.720 15.340 389.980 15.600 ;
      LAYER met2 ;
        RECT 936.570 1100.580 936.850 1104.000 ;
        RECT 936.570 1100.000 936.860 1100.580 ;
        RECT 936.720 1089.350 936.860 1100.000 ;
        RECT 389.720 1089.030 389.980 1089.350 ;
        RECT 936.660 1089.030 936.920 1089.350 ;
        RECT 389.780 15.630 389.920 1089.030 ;
        RECT 252.640 15.310 252.900 15.630 ;
        RECT 389.720 15.310 389.980 15.630 ;
        RECT 252.700 2.000 252.840 15.310 ;
        RECT 252.490 -4.000 253.050 2.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 927.890 1083.480 928.210 1083.540 ;
        RECT 942.610 1083.480 942.930 1083.540 ;
        RECT 927.890 1083.340 942.930 1083.480 ;
        RECT 927.890 1083.280 928.210 1083.340 ;
        RECT 942.610 1083.280 942.930 1083.340 ;
        RECT 270.090 20.300 270.410 20.360 ;
        RECT 927.890 20.300 928.210 20.360 ;
        RECT 270.090 20.160 928.210 20.300 ;
        RECT 270.090 20.100 270.410 20.160 ;
        RECT 927.890 20.100 928.210 20.160 ;
      LAYER via ;
        RECT 927.920 1083.280 928.180 1083.540 ;
        RECT 942.640 1083.280 942.900 1083.540 ;
        RECT 270.120 20.100 270.380 20.360 ;
        RECT 927.920 20.100 928.180 20.360 ;
      LAYER met2 ;
        RECT 942.550 1100.580 942.830 1104.000 ;
        RECT 942.550 1100.000 942.840 1100.580 ;
        RECT 942.700 1083.570 942.840 1100.000 ;
        RECT 927.920 1083.250 928.180 1083.570 ;
        RECT 942.640 1083.250 942.900 1083.570 ;
        RECT 927.980 20.390 928.120 1083.250 ;
        RECT 270.120 20.070 270.380 20.390 ;
        RECT 927.920 20.070 928.180 20.390 ;
        RECT 270.180 2.000 270.320 20.070 ;
        RECT 269.970 -4.000 270.530 2.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 397.125 14.705 397.295 15.895 ;
      LAYER mcon ;
        RECT 397.125 15.725 397.295 15.895 ;
      LAYER met1 ;
        RECT 424.190 1086.200 424.510 1086.260 ;
        RECT 948.590 1086.200 948.910 1086.260 ;
        RECT 424.190 1086.060 948.910 1086.200 ;
        RECT 424.190 1086.000 424.510 1086.060 ;
        RECT 948.590 1086.000 948.910 1086.060 ;
        RECT 288.030 15.880 288.350 15.940 ;
        RECT 397.065 15.880 397.355 15.925 ;
        RECT 288.030 15.740 397.355 15.880 ;
        RECT 288.030 15.680 288.350 15.740 ;
        RECT 397.065 15.695 397.355 15.740 ;
        RECT 397.065 14.860 397.355 14.905 ;
        RECT 424.190 14.860 424.510 14.920 ;
        RECT 397.065 14.720 424.510 14.860 ;
        RECT 397.065 14.675 397.355 14.720 ;
        RECT 424.190 14.660 424.510 14.720 ;
      LAYER via ;
        RECT 424.220 1086.000 424.480 1086.260 ;
        RECT 948.620 1086.000 948.880 1086.260 ;
        RECT 288.060 15.680 288.320 15.940 ;
        RECT 424.220 14.660 424.480 14.920 ;
      LAYER met2 ;
        RECT 948.530 1100.580 948.810 1104.000 ;
        RECT 948.530 1100.000 948.820 1100.580 ;
        RECT 948.680 1086.290 948.820 1100.000 ;
        RECT 424.220 1085.970 424.480 1086.290 ;
        RECT 948.620 1085.970 948.880 1086.290 ;
        RECT 288.060 15.650 288.320 15.970 ;
        RECT 288.120 2.000 288.260 15.650 ;
        RECT 424.280 14.950 424.420 1085.970 ;
        RECT 424.220 14.630 424.480 14.950 ;
        RECT 287.910 -4.000 288.470 2.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 934.790 1087.560 935.110 1087.620 ;
        RECT 955.030 1087.560 955.350 1087.620 ;
        RECT 934.790 1087.420 955.350 1087.560 ;
        RECT 934.790 1087.360 935.110 1087.420 ;
        RECT 955.030 1087.360 955.350 1087.420 ;
        RECT 305.970 20.640 306.290 20.700 ;
        RECT 934.790 20.640 935.110 20.700 ;
        RECT 305.970 20.500 935.110 20.640 ;
        RECT 305.970 20.440 306.290 20.500 ;
        RECT 934.790 20.440 935.110 20.500 ;
      LAYER via ;
        RECT 934.820 1087.360 935.080 1087.620 ;
        RECT 955.060 1087.360 955.320 1087.620 ;
        RECT 306.000 20.440 306.260 20.700 ;
        RECT 934.820 20.440 935.080 20.700 ;
      LAYER met2 ;
        RECT 954.970 1100.580 955.250 1104.000 ;
        RECT 954.970 1100.000 955.260 1100.580 ;
        RECT 955.120 1087.650 955.260 1100.000 ;
        RECT 934.820 1087.330 935.080 1087.650 ;
        RECT 955.060 1087.330 955.320 1087.650 ;
        RECT 934.880 20.730 935.020 1087.330 ;
        RECT 306.000 20.410 306.260 20.730 ;
        RECT 934.820 20.410 935.080 20.730 ;
        RECT 306.060 2.000 306.200 20.410 ;
        RECT 305.850 -4.000 306.410 2.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 907.265 1083.325 907.435 1086.555 ;
      LAYER mcon ;
        RECT 907.265 1086.385 907.435 1086.555 ;
      LAYER met1 ;
        RECT 907.205 1086.540 907.495 1086.585 ;
        RECT 961.010 1086.540 961.330 1086.600 ;
        RECT 907.205 1086.400 961.330 1086.540 ;
        RECT 907.205 1086.355 907.495 1086.400 ;
        RECT 961.010 1086.340 961.330 1086.400 ;
        RECT 534.590 1083.480 534.910 1083.540 ;
        RECT 907.205 1083.480 907.495 1083.525 ;
        RECT 534.590 1083.340 907.495 1083.480 ;
        RECT 534.590 1083.280 534.910 1083.340 ;
        RECT 907.205 1083.295 907.495 1083.340 ;
        RECT 323.910 14.520 324.230 14.580 ;
        RECT 534.590 14.520 534.910 14.580 ;
        RECT 323.910 14.380 534.910 14.520 ;
        RECT 323.910 14.320 324.230 14.380 ;
        RECT 534.590 14.320 534.910 14.380 ;
      LAYER via ;
        RECT 961.040 1086.340 961.300 1086.600 ;
        RECT 534.620 1083.280 534.880 1083.540 ;
        RECT 323.940 14.320 324.200 14.580 ;
        RECT 534.620 14.320 534.880 14.580 ;
      LAYER met2 ;
        RECT 960.950 1100.580 961.230 1104.000 ;
        RECT 960.950 1100.000 961.240 1100.580 ;
        RECT 961.100 1086.630 961.240 1100.000 ;
        RECT 961.040 1086.310 961.300 1086.630 ;
        RECT 534.620 1083.250 534.880 1083.570 ;
        RECT 534.680 14.610 534.820 1083.250 ;
        RECT 323.940 14.290 324.200 14.610 ;
        RECT 534.620 14.290 534.880 14.610 ;
        RECT 324.000 2.000 324.140 14.290 ;
        RECT 323.790 -4.000 324.350 2.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 941.690 1088.240 942.010 1088.300 ;
        RECT 966.990 1088.240 967.310 1088.300 ;
        RECT 941.690 1088.100 967.310 1088.240 ;
        RECT 941.690 1088.040 942.010 1088.100 ;
        RECT 966.990 1088.040 967.310 1088.100 ;
        RECT 941.690 16.900 942.010 16.960 ;
        RECT 358.960 16.760 942.010 16.900 ;
        RECT 341.390 16.560 341.710 16.620 ;
        RECT 358.960 16.560 359.100 16.760 ;
        RECT 941.690 16.700 942.010 16.760 ;
        RECT 341.390 16.420 359.100 16.560 ;
        RECT 341.390 16.360 341.710 16.420 ;
      LAYER via ;
        RECT 941.720 1088.040 941.980 1088.300 ;
        RECT 967.020 1088.040 967.280 1088.300 ;
        RECT 341.420 16.360 341.680 16.620 ;
        RECT 941.720 16.700 941.980 16.960 ;
      LAYER met2 ;
        RECT 966.930 1100.580 967.210 1104.000 ;
        RECT 966.930 1100.000 967.220 1100.580 ;
        RECT 967.080 1088.330 967.220 1100.000 ;
        RECT 941.720 1088.010 941.980 1088.330 ;
        RECT 967.020 1088.010 967.280 1088.330 ;
        RECT 941.780 16.990 941.920 1088.010 ;
        RECT 941.720 16.670 941.980 16.990 ;
        RECT 341.420 16.330 341.680 16.650 ;
        RECT 341.480 2.000 341.620 16.330 ;
        RECT 341.270 -4.000 341.830 2.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 396.665 14.025 396.835 14.875 ;
      LAYER mcon ;
        RECT 396.665 14.705 396.835 14.875 ;
      LAYER met1 ;
        RECT 431.090 1089.600 431.410 1089.660 ;
        RECT 973.430 1089.600 973.750 1089.660 ;
        RECT 431.090 1089.460 973.750 1089.600 ;
        RECT 431.090 1089.400 431.410 1089.460 ;
        RECT 973.430 1089.400 973.750 1089.460 ;
        RECT 359.330 14.860 359.650 14.920 ;
        RECT 396.605 14.860 396.895 14.905 ;
        RECT 359.330 14.720 396.895 14.860 ;
        RECT 359.330 14.660 359.650 14.720 ;
        RECT 396.605 14.675 396.895 14.720 ;
        RECT 396.605 14.180 396.895 14.225 ;
        RECT 431.090 14.180 431.410 14.240 ;
        RECT 396.605 14.040 431.410 14.180 ;
        RECT 396.605 13.995 396.895 14.040 ;
        RECT 431.090 13.980 431.410 14.040 ;
      LAYER via ;
        RECT 431.120 1089.400 431.380 1089.660 ;
        RECT 973.460 1089.400 973.720 1089.660 ;
        RECT 359.360 14.660 359.620 14.920 ;
        RECT 431.120 13.980 431.380 14.240 ;
      LAYER met2 ;
        RECT 973.370 1100.580 973.650 1104.000 ;
        RECT 973.370 1100.000 973.660 1100.580 ;
        RECT 973.520 1089.690 973.660 1100.000 ;
        RECT 431.120 1089.370 431.380 1089.690 ;
        RECT 973.460 1089.370 973.720 1089.690 ;
        RECT 359.360 14.630 359.620 14.950 ;
        RECT 359.420 2.000 359.560 14.630 ;
        RECT 431.180 14.270 431.320 1089.370 ;
        RECT 431.120 13.950 431.380 14.270 ;
        RECT 359.210 -4.000 359.770 2.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 955.565 372.725 955.735 420.835 ;
        RECT 412.765 16.405 414.315 16.575 ;
        RECT 397.585 13.685 397.755 15.895 ;
        RECT 412.765 15.725 412.935 16.405 ;
      LAYER mcon ;
        RECT 955.565 420.665 955.735 420.835 ;
        RECT 414.145 16.405 414.315 16.575 ;
        RECT 397.585 15.725 397.755 15.895 ;
      LAYER met1 ;
        RECT 955.950 1088.920 956.270 1088.980 ;
        RECT 979.410 1088.920 979.730 1088.980 ;
        RECT 955.950 1088.780 979.730 1088.920 ;
        RECT 955.950 1088.720 956.270 1088.780 ;
        RECT 979.410 1088.720 979.730 1088.780 ;
        RECT 955.490 765.920 955.810 765.980 ;
        RECT 955.950 765.920 956.270 765.980 ;
        RECT 955.490 765.780 956.270 765.920 ;
        RECT 955.490 765.720 955.810 765.780 ;
        RECT 955.950 765.720 956.270 765.780 ;
        RECT 955.490 642.160 955.810 642.220 ;
        RECT 955.120 642.020 955.810 642.160 ;
        RECT 955.120 641.540 955.260 642.020 ;
        RECT 955.490 641.960 955.810 642.020 ;
        RECT 955.030 641.280 955.350 641.540 ;
        RECT 955.030 627.880 955.350 627.940 ;
        RECT 955.950 627.880 956.270 627.940 ;
        RECT 955.030 627.740 956.270 627.880 ;
        RECT 955.030 627.680 955.350 627.740 ;
        RECT 955.950 627.680 956.270 627.740 ;
        RECT 955.030 476.240 955.350 476.300 ;
        RECT 955.950 476.240 956.270 476.300 ;
        RECT 955.030 476.100 956.270 476.240 ;
        RECT 955.030 476.040 955.350 476.100 ;
        RECT 955.950 476.040 956.270 476.100 ;
        RECT 955.950 435.100 956.270 435.160 ;
        RECT 955.580 434.960 956.270 435.100 ;
        RECT 955.580 434.820 955.720 434.960 ;
        RECT 955.950 434.900 956.270 434.960 ;
        RECT 955.490 434.560 955.810 434.820 ;
        RECT 955.490 420.820 955.810 420.880 ;
        RECT 955.295 420.680 955.810 420.820 ;
        RECT 955.490 420.620 955.810 420.680 ;
        RECT 955.505 372.880 955.795 372.925 ;
        RECT 956.410 372.880 956.730 372.940 ;
        RECT 955.505 372.740 956.730 372.880 ;
        RECT 955.505 372.695 955.795 372.740 ;
        RECT 956.410 372.680 956.730 372.740 ;
        RECT 954.570 220.900 954.890 220.960 ;
        RECT 955.490 220.900 955.810 220.960 ;
        RECT 954.570 220.760 955.810 220.900 ;
        RECT 954.570 220.700 954.890 220.760 ;
        RECT 955.490 220.700 955.810 220.760 ;
        RECT 955.950 193.360 956.270 193.420 ;
        RECT 955.580 193.220 956.270 193.360 ;
        RECT 955.580 193.080 955.720 193.220 ;
        RECT 955.950 193.160 956.270 193.220 ;
        RECT 955.490 192.820 955.810 193.080 ;
        RECT 414.085 16.560 414.375 16.605 ;
        RECT 955.030 16.560 955.350 16.620 ;
        RECT 414.085 16.420 955.350 16.560 ;
        RECT 414.085 16.375 414.375 16.420 ;
        RECT 955.030 16.360 955.350 16.420 ;
        RECT 397.525 15.880 397.815 15.925 ;
        RECT 412.705 15.880 412.995 15.925 ;
        RECT 397.525 15.740 412.995 15.880 ;
        RECT 397.525 15.695 397.815 15.740 ;
        RECT 412.705 15.695 412.995 15.740 ;
        RECT 377.270 14.180 377.590 14.240 ;
        RECT 377.270 14.040 396.360 14.180 ;
        RECT 377.270 13.980 377.590 14.040 ;
        RECT 396.220 13.840 396.360 14.040 ;
        RECT 397.525 13.840 397.815 13.885 ;
        RECT 396.220 13.700 397.815 13.840 ;
        RECT 397.525 13.655 397.815 13.700 ;
      LAYER via ;
        RECT 955.980 1088.720 956.240 1088.980 ;
        RECT 979.440 1088.720 979.700 1088.980 ;
        RECT 955.520 765.720 955.780 765.980 ;
        RECT 955.980 765.720 956.240 765.980 ;
        RECT 955.520 641.960 955.780 642.220 ;
        RECT 955.060 641.280 955.320 641.540 ;
        RECT 955.060 627.680 955.320 627.940 ;
        RECT 955.980 627.680 956.240 627.940 ;
        RECT 955.060 476.040 955.320 476.300 ;
        RECT 955.980 476.040 956.240 476.300 ;
        RECT 955.980 434.900 956.240 435.160 ;
        RECT 955.520 434.560 955.780 434.820 ;
        RECT 955.520 420.620 955.780 420.880 ;
        RECT 956.440 372.680 956.700 372.940 ;
        RECT 954.600 220.700 954.860 220.960 ;
        RECT 955.520 220.700 955.780 220.960 ;
        RECT 955.980 193.160 956.240 193.420 ;
        RECT 955.520 192.820 955.780 193.080 ;
        RECT 955.060 16.360 955.320 16.620 ;
        RECT 377.300 13.980 377.560 14.240 ;
      LAYER met2 ;
        RECT 979.350 1100.580 979.630 1104.000 ;
        RECT 979.350 1100.000 979.640 1100.580 ;
        RECT 979.500 1089.010 979.640 1100.000 ;
        RECT 955.980 1088.690 956.240 1089.010 ;
        RECT 979.440 1088.690 979.700 1089.010 ;
        RECT 956.040 1041.490 956.180 1088.690 ;
        RECT 955.580 1041.350 956.180 1041.490 ;
        RECT 955.580 980.290 955.720 1041.350 ;
        RECT 955.120 980.150 955.720 980.290 ;
        RECT 955.120 979.610 955.260 980.150 ;
        RECT 955.120 979.470 955.720 979.610 ;
        RECT 955.580 835.450 955.720 979.470 ;
        RECT 955.120 835.310 955.720 835.450 ;
        RECT 955.120 834.770 955.260 835.310 ;
        RECT 955.120 834.630 955.720 834.770 ;
        RECT 955.580 773.685 955.720 834.630 ;
        RECT 955.510 773.315 955.790 773.685 ;
        RECT 955.510 772.635 955.790 773.005 ;
        RECT 955.580 766.010 955.720 772.635 ;
        RECT 955.520 765.690 955.780 766.010 ;
        RECT 955.980 765.690 956.240 766.010 ;
        RECT 956.040 699.450 956.180 765.690 ;
        RECT 955.580 699.310 956.180 699.450 ;
        RECT 955.580 642.250 955.720 699.310 ;
        RECT 955.520 641.930 955.780 642.250 ;
        RECT 955.060 641.250 955.320 641.570 ;
        RECT 955.120 627.970 955.260 641.250 ;
        RECT 955.060 627.650 955.320 627.970 ;
        RECT 955.980 627.650 956.240 627.970 ;
        RECT 956.040 602.890 956.180 627.650 ;
        RECT 955.580 602.750 956.180 602.890 ;
        RECT 955.580 532.285 955.720 602.750 ;
        RECT 955.510 531.915 955.790 532.285 ;
        RECT 955.050 531.235 955.330 531.605 ;
        RECT 955.120 476.330 955.260 531.235 ;
        RECT 955.060 476.010 955.320 476.330 ;
        RECT 955.980 476.010 956.240 476.330 ;
        RECT 956.040 435.190 956.180 476.010 ;
        RECT 955.980 434.870 956.240 435.190 ;
        RECT 955.520 434.530 955.780 434.850 ;
        RECT 955.580 420.910 955.720 434.530 ;
        RECT 955.520 420.590 955.780 420.910 ;
        RECT 956.440 372.650 956.700 372.970 ;
        RECT 956.500 372.370 956.640 372.650 ;
        RECT 955.580 372.230 956.640 372.370 ;
        RECT 955.580 325.565 955.720 372.230 ;
        RECT 955.510 325.195 955.790 325.565 ;
        RECT 955.050 324.770 955.330 324.885 ;
        RECT 955.050 324.630 955.720 324.770 ;
        RECT 955.050 324.515 955.330 324.630 ;
        RECT 955.580 270.485 955.720 324.630 ;
        RECT 955.510 270.115 955.790 270.485 ;
        RECT 955.510 269.435 955.790 269.805 ;
        RECT 955.580 269.125 955.720 269.435 ;
        RECT 954.590 268.755 954.870 269.125 ;
        RECT 955.510 268.755 955.790 269.125 ;
        RECT 954.660 220.990 954.800 268.755 ;
        RECT 955.580 220.990 955.720 221.145 ;
        RECT 954.600 220.670 954.860 220.990 ;
        RECT 955.520 220.730 955.780 220.990 ;
        RECT 955.520 220.670 956.180 220.730 ;
        RECT 955.580 220.590 956.180 220.670 ;
        RECT 956.040 193.450 956.180 220.590 ;
        RECT 955.980 193.130 956.240 193.450 ;
        RECT 955.520 192.790 955.780 193.110 ;
        RECT 955.580 62.290 955.720 192.790 ;
        RECT 955.120 62.150 955.720 62.290 ;
        RECT 955.120 16.650 955.260 62.150 ;
        RECT 955.060 16.330 955.320 16.650 ;
        RECT 377.300 13.950 377.560 14.270 ;
        RECT 377.360 2.000 377.500 13.950 ;
        RECT 377.150 -4.000 377.710 2.000 ;
      LAYER via2 ;
        RECT 955.510 773.360 955.790 773.640 ;
        RECT 955.510 772.680 955.790 772.960 ;
        RECT 955.510 531.960 955.790 532.240 ;
        RECT 955.050 531.280 955.330 531.560 ;
        RECT 955.510 325.240 955.790 325.520 ;
        RECT 955.050 324.560 955.330 324.840 ;
        RECT 955.510 270.160 955.790 270.440 ;
        RECT 955.510 269.480 955.790 269.760 ;
        RECT 954.590 268.800 954.870 269.080 ;
        RECT 955.510 268.800 955.790 269.080 ;
      LAYER met3 ;
        RECT 955.485 773.650 955.815 773.665 ;
        RECT 955.270 773.335 955.815 773.650 ;
        RECT 955.270 772.985 955.570 773.335 ;
        RECT 955.270 772.670 955.815 772.985 ;
        RECT 955.485 772.655 955.815 772.670 ;
        RECT 955.485 532.250 955.815 532.265 ;
        RECT 955.270 531.935 955.815 532.250 ;
        RECT 955.270 531.585 955.570 531.935 ;
        RECT 955.025 531.270 955.570 531.585 ;
        RECT 955.025 531.255 955.355 531.270 ;
        RECT 955.485 325.530 955.815 325.545 ;
        RECT 955.270 325.215 955.815 325.530 ;
        RECT 955.270 324.865 955.570 325.215 ;
        RECT 955.025 324.550 955.570 324.865 ;
        RECT 955.025 324.535 955.355 324.550 ;
        RECT 955.485 270.450 955.815 270.465 ;
        RECT 955.485 270.150 956.490 270.450 ;
        RECT 955.485 270.135 955.815 270.150 ;
        RECT 955.485 269.770 955.815 269.785 ;
        RECT 956.190 269.770 956.490 270.150 ;
        RECT 955.485 269.470 956.490 269.770 ;
        RECT 955.485 269.455 955.815 269.470 ;
        RECT 954.565 269.090 954.895 269.105 ;
        RECT 955.485 269.090 955.815 269.105 ;
        RECT 954.565 268.790 955.815 269.090 ;
        RECT 954.565 268.775 954.895 268.790 ;
        RECT 955.485 268.775 955.815 268.790 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 430.245 14.705 430.415 15.555 ;
      LAYER mcon ;
        RECT 430.245 15.385 430.415 15.555 ;
      LAYER met1 ;
        RECT 444.890 1089.940 445.210 1090.000 ;
        RECT 985.390 1089.940 985.710 1090.000 ;
        RECT 444.890 1089.800 985.710 1089.940 ;
        RECT 444.890 1089.740 445.210 1089.800 ;
        RECT 985.390 1089.740 985.710 1089.800 ;
        RECT 395.210 15.540 395.530 15.600 ;
        RECT 430.185 15.540 430.475 15.585 ;
        RECT 395.210 15.400 430.475 15.540 ;
        RECT 395.210 15.340 395.530 15.400 ;
        RECT 430.185 15.355 430.475 15.400 ;
        RECT 430.185 14.860 430.475 14.905 ;
        RECT 444.890 14.860 445.210 14.920 ;
        RECT 430.185 14.720 445.210 14.860 ;
        RECT 430.185 14.675 430.475 14.720 ;
        RECT 444.890 14.660 445.210 14.720 ;
      LAYER via ;
        RECT 444.920 1089.740 445.180 1090.000 ;
        RECT 985.420 1089.740 985.680 1090.000 ;
        RECT 395.240 15.340 395.500 15.600 ;
        RECT 444.920 14.660 445.180 14.920 ;
      LAYER met2 ;
        RECT 985.330 1100.580 985.610 1104.000 ;
        RECT 985.330 1100.000 985.620 1100.580 ;
        RECT 985.480 1090.030 985.620 1100.000 ;
        RECT 444.920 1089.710 445.180 1090.030 ;
        RECT 985.420 1089.710 985.680 1090.030 ;
        RECT 395.240 15.310 395.500 15.630 ;
        RECT 395.300 2.000 395.440 15.310 ;
        RECT 444.980 14.950 445.120 1089.710 ;
        RECT 444.920 14.630 445.180 14.950 ;
        RECT 395.090 -4.000 395.650 2.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 962.850 1086.200 963.170 1086.260 ;
        RECT 991.830 1086.200 992.150 1086.260 ;
        RECT 962.850 1086.060 992.150 1086.200 ;
        RECT 962.850 1086.000 963.170 1086.060 ;
        RECT 991.830 1086.000 992.150 1086.060 ;
        RECT 962.850 16.220 963.170 16.280 ;
        RECT 438.540 16.080 963.170 16.220 ;
        RECT 413.150 15.880 413.470 15.940 ;
        RECT 438.540 15.880 438.680 16.080 ;
        RECT 962.850 16.020 963.170 16.080 ;
        RECT 413.150 15.740 438.680 15.880 ;
        RECT 413.150 15.680 413.470 15.740 ;
      LAYER via ;
        RECT 962.880 1086.000 963.140 1086.260 ;
        RECT 991.860 1086.000 992.120 1086.260 ;
        RECT 413.180 15.680 413.440 15.940 ;
        RECT 962.880 16.020 963.140 16.280 ;
      LAYER met2 ;
        RECT 991.770 1100.580 992.050 1104.000 ;
        RECT 991.770 1100.000 992.060 1100.580 ;
        RECT 991.920 1086.290 992.060 1100.000 ;
        RECT 962.880 1085.970 963.140 1086.290 ;
        RECT 991.860 1085.970 992.120 1086.290 ;
        RECT 962.940 16.310 963.080 1085.970 ;
        RECT 962.880 15.990 963.140 16.310 ;
        RECT 413.180 15.650 413.440 15.970 ;
        RECT 413.240 2.000 413.380 15.650 ;
        RECT 413.030 -4.000 413.590 2.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 875.450 1086.880 875.770 1086.940 ;
        RECT 835.980 1086.740 875.770 1086.880 ;
        RECT 86.090 1086.540 86.410 1086.600 ;
        RECT 835.980 1086.540 836.120 1086.740 ;
        RECT 875.450 1086.680 875.770 1086.740 ;
        RECT 86.090 1086.400 836.120 1086.540 ;
        RECT 86.090 1086.340 86.410 1086.400 ;
        RECT 74.130 19.960 74.450 20.020 ;
        RECT 86.090 19.960 86.410 20.020 ;
        RECT 74.130 19.820 86.410 19.960 ;
        RECT 74.130 19.760 74.450 19.820 ;
        RECT 86.090 19.760 86.410 19.820 ;
      LAYER via ;
        RECT 86.120 1086.340 86.380 1086.600 ;
        RECT 875.480 1086.680 875.740 1086.940 ;
        RECT 74.160 19.760 74.420 20.020 ;
        RECT 86.120 19.760 86.380 20.020 ;
      LAYER met2 ;
        RECT 875.390 1100.580 875.670 1104.000 ;
        RECT 875.390 1100.000 875.680 1100.580 ;
        RECT 875.540 1086.970 875.680 1100.000 ;
        RECT 875.480 1086.650 875.740 1086.970 ;
        RECT 86.120 1086.310 86.380 1086.630 ;
        RECT 86.180 20.050 86.320 1086.310 ;
        RECT 74.160 19.730 74.420 20.050 ;
        RECT 86.120 19.730 86.380 20.050 ;
        RECT 74.220 2.000 74.360 19.730 ;
        RECT 74.010 -4.000 74.570 2.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 962.390 1086.540 962.710 1086.600 ;
        RECT 997.810 1086.540 998.130 1086.600 ;
        RECT 962.390 1086.400 998.130 1086.540 ;
        RECT 962.390 1086.340 962.710 1086.400 ;
        RECT 997.810 1086.340 998.130 1086.400 ;
        RECT 962.390 15.880 962.710 15.940 ;
        RECT 448.660 15.740 962.710 15.880 ;
        RECT 430.630 15.540 430.950 15.600 ;
        RECT 448.660 15.540 448.800 15.740 ;
        RECT 962.390 15.680 962.710 15.740 ;
        RECT 430.630 15.400 448.800 15.540 ;
        RECT 430.630 15.340 430.950 15.400 ;
      LAYER via ;
        RECT 962.420 1086.340 962.680 1086.600 ;
        RECT 997.840 1086.340 998.100 1086.600 ;
        RECT 430.660 15.340 430.920 15.600 ;
        RECT 962.420 15.680 962.680 15.940 ;
      LAYER met2 ;
        RECT 997.750 1100.580 998.030 1104.000 ;
        RECT 997.750 1100.000 998.040 1100.580 ;
        RECT 997.900 1086.630 998.040 1100.000 ;
        RECT 962.420 1086.310 962.680 1086.630 ;
        RECT 997.840 1086.310 998.100 1086.630 ;
        RECT 962.480 15.970 962.620 1086.310 ;
        RECT 962.420 15.650 962.680 15.970 ;
        RECT 430.660 15.310 430.920 15.630 ;
        RECT 430.720 2.000 430.860 15.310 ;
        RECT 430.510 -4.000 431.070 2.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 479.390 1085.860 479.710 1085.920 ;
        RECT 1003.790 1085.860 1004.110 1085.920 ;
        RECT 479.390 1085.720 1004.110 1085.860 ;
        RECT 479.390 1085.660 479.710 1085.720 ;
        RECT 1003.790 1085.660 1004.110 1085.720 ;
        RECT 448.570 14.860 448.890 14.920 ;
        RECT 479.390 14.860 479.710 14.920 ;
        RECT 448.570 14.720 479.710 14.860 ;
        RECT 448.570 14.660 448.890 14.720 ;
        RECT 479.390 14.660 479.710 14.720 ;
      LAYER via ;
        RECT 479.420 1085.660 479.680 1085.920 ;
        RECT 1003.820 1085.660 1004.080 1085.920 ;
        RECT 448.600 14.660 448.860 14.920 ;
        RECT 479.420 14.660 479.680 14.920 ;
      LAYER met2 ;
        RECT 1003.730 1100.580 1004.010 1104.000 ;
        RECT 1003.730 1100.000 1004.020 1100.580 ;
        RECT 1003.880 1085.950 1004.020 1100.000 ;
        RECT 479.420 1085.630 479.680 1085.950 ;
        RECT 1003.820 1085.630 1004.080 1085.950 ;
        RECT 479.480 14.950 479.620 1085.630 ;
        RECT 448.600 14.630 448.860 14.950 ;
        RECT 479.420 14.630 479.680 14.950 ;
        RECT 448.660 2.000 448.800 14.630 ;
        RECT 448.450 -4.000 449.010 2.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 969.290 1064.440 969.610 1064.500 ;
        RECT 1010.230 1064.440 1010.550 1064.500 ;
        RECT 969.290 1064.300 1010.550 1064.440 ;
        RECT 969.290 1064.240 969.610 1064.300 ;
        RECT 1010.230 1064.240 1010.550 1064.300 ;
        RECT 466.510 15.540 466.830 15.600 ;
        RECT 969.290 15.540 969.610 15.600 ;
        RECT 466.510 15.400 969.610 15.540 ;
        RECT 466.510 15.340 466.830 15.400 ;
        RECT 969.290 15.340 969.610 15.400 ;
      LAYER via ;
        RECT 969.320 1064.240 969.580 1064.500 ;
        RECT 1010.260 1064.240 1010.520 1064.500 ;
        RECT 466.540 15.340 466.800 15.600 ;
        RECT 969.320 15.340 969.580 15.600 ;
      LAYER met2 ;
        RECT 1010.170 1100.580 1010.450 1104.000 ;
        RECT 1010.170 1100.000 1010.460 1100.580 ;
        RECT 1010.320 1064.530 1010.460 1100.000 ;
        RECT 969.320 1064.210 969.580 1064.530 ;
        RECT 1010.260 1064.210 1010.520 1064.530 ;
        RECT 969.380 15.630 969.520 1064.210 ;
        RECT 466.540 15.310 466.800 15.630 ;
        RECT 969.320 15.310 969.580 15.630 ;
        RECT 466.600 2.000 466.740 15.310 ;
        RECT 466.390 -4.000 466.950 2.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 513.890 1085.180 514.210 1085.240 ;
        RECT 1016.210 1085.180 1016.530 1085.240 ;
        RECT 513.890 1085.040 1016.530 1085.180 ;
        RECT 513.890 1084.980 514.210 1085.040 ;
        RECT 1016.210 1084.980 1016.530 1085.040 ;
        RECT 484.450 15.200 484.770 15.260 ;
        RECT 512.970 15.200 513.290 15.260 ;
        RECT 484.450 15.060 513.290 15.200 ;
        RECT 484.450 15.000 484.770 15.060 ;
        RECT 512.970 15.000 513.290 15.060 ;
      LAYER via ;
        RECT 513.920 1084.980 514.180 1085.240 ;
        RECT 1016.240 1084.980 1016.500 1085.240 ;
        RECT 484.480 15.000 484.740 15.260 ;
        RECT 513.000 15.000 513.260 15.260 ;
      LAYER met2 ;
        RECT 1016.150 1100.580 1016.430 1104.000 ;
        RECT 1016.150 1100.000 1016.440 1100.580 ;
        RECT 1016.300 1085.270 1016.440 1100.000 ;
        RECT 513.920 1084.950 514.180 1085.270 ;
        RECT 1016.240 1084.950 1016.500 1085.270 ;
        RECT 513.980 16.050 514.120 1084.950 ;
        RECT 513.060 15.910 514.120 16.050 ;
        RECT 513.060 15.290 513.200 15.910 ;
        RECT 484.480 14.970 484.740 15.290 ;
        RECT 513.000 14.970 513.260 15.290 ;
        RECT 484.540 2.000 484.680 14.970 ;
        RECT 484.330 -4.000 484.890 2.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 976.650 1087.560 976.970 1087.620 ;
        RECT 1022.190 1087.560 1022.510 1087.620 ;
        RECT 976.650 1087.420 1022.510 1087.560 ;
        RECT 976.650 1087.360 976.970 1087.420 ;
        RECT 1022.190 1087.360 1022.510 1087.420 ;
        RECT 976.650 15.200 976.970 15.260 ;
        RECT 559.060 15.060 976.970 15.200 ;
        RECT 502.390 14.860 502.710 14.920 ;
        RECT 559.060 14.860 559.200 15.060 ;
        RECT 976.650 15.000 976.970 15.060 ;
        RECT 502.390 14.720 559.200 14.860 ;
        RECT 502.390 14.660 502.710 14.720 ;
      LAYER via ;
        RECT 976.680 1087.360 976.940 1087.620 ;
        RECT 1022.220 1087.360 1022.480 1087.620 ;
        RECT 502.420 14.660 502.680 14.920 ;
        RECT 976.680 15.000 976.940 15.260 ;
      LAYER met2 ;
        RECT 1022.130 1100.580 1022.410 1104.000 ;
        RECT 1022.130 1100.000 1022.420 1100.580 ;
        RECT 1022.280 1087.650 1022.420 1100.000 ;
        RECT 976.680 1087.330 976.940 1087.650 ;
        RECT 1022.220 1087.330 1022.480 1087.650 ;
        RECT 976.740 15.290 976.880 1087.330 ;
        RECT 976.680 14.970 976.940 15.290 ;
        RECT 502.420 14.630 502.680 14.950 ;
        RECT 502.480 2.000 502.620 14.630 ;
        RECT 502.270 -4.000 502.830 2.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 524.010 1085.520 524.330 1085.580 ;
        RECT 1028.170 1085.520 1028.490 1085.580 ;
        RECT 524.010 1085.380 1028.490 1085.520 ;
        RECT 524.010 1085.320 524.330 1085.380 ;
        RECT 1028.170 1085.320 1028.490 1085.380 ;
        RECT 519.870 15.200 520.190 15.260 ;
        RECT 524.010 15.200 524.330 15.260 ;
        RECT 519.870 15.060 524.330 15.200 ;
        RECT 519.870 15.000 520.190 15.060 ;
        RECT 524.010 15.000 524.330 15.060 ;
      LAYER via ;
        RECT 524.040 1085.320 524.300 1085.580 ;
        RECT 1028.200 1085.320 1028.460 1085.580 ;
        RECT 519.900 15.000 520.160 15.260 ;
        RECT 524.040 15.000 524.300 15.260 ;
      LAYER met2 ;
        RECT 1028.110 1100.580 1028.390 1104.000 ;
        RECT 1028.110 1100.000 1028.400 1100.580 ;
        RECT 1028.260 1085.610 1028.400 1100.000 ;
        RECT 524.040 1085.290 524.300 1085.610 ;
        RECT 1028.200 1085.290 1028.460 1085.610 ;
        RECT 524.100 15.290 524.240 1085.290 ;
        RECT 519.900 14.970 520.160 15.290 ;
        RECT 524.040 14.970 524.300 15.290 ;
        RECT 519.960 2.000 520.100 14.970 ;
        RECT 519.750 -4.000 520.310 2.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 976.190 1087.900 976.510 1087.960 ;
        RECT 1034.610 1087.900 1034.930 1087.960 ;
        RECT 976.190 1087.760 1034.930 1087.900 ;
        RECT 976.190 1087.700 976.510 1087.760 ;
        RECT 1034.610 1087.700 1034.930 1087.760 ;
        RECT 976.190 14.860 976.510 14.920 ;
        RECT 607.820 14.720 976.510 14.860 ;
        RECT 537.810 14.180 538.130 14.240 ;
        RECT 607.820 14.180 607.960 14.720 ;
        RECT 976.190 14.660 976.510 14.720 ;
        RECT 537.810 14.040 607.960 14.180 ;
        RECT 537.810 13.980 538.130 14.040 ;
      LAYER via ;
        RECT 976.220 1087.700 976.480 1087.960 ;
        RECT 1034.640 1087.700 1034.900 1087.960 ;
        RECT 537.840 13.980 538.100 14.240 ;
        RECT 976.220 14.660 976.480 14.920 ;
      LAYER met2 ;
        RECT 1034.550 1100.580 1034.830 1104.000 ;
        RECT 1034.550 1100.000 1034.840 1100.580 ;
        RECT 1034.700 1087.990 1034.840 1100.000 ;
        RECT 976.220 1087.670 976.480 1087.990 ;
        RECT 1034.640 1087.670 1034.900 1087.990 ;
        RECT 976.280 14.950 976.420 1087.670 ;
        RECT 976.220 14.630 976.480 14.950 ;
        RECT 537.840 13.950 538.100 14.270 ;
        RECT 537.900 2.000 538.040 13.950 ;
        RECT 537.690 -4.000 538.250 2.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 558.510 1084.840 558.830 1084.900 ;
        RECT 1040.590 1084.840 1040.910 1084.900 ;
        RECT 558.510 1084.700 1040.910 1084.840 ;
        RECT 558.510 1084.640 558.830 1084.700 ;
        RECT 1040.590 1084.640 1040.910 1084.700 ;
        RECT 555.750 15.200 556.070 15.260 ;
        RECT 558.510 15.200 558.830 15.260 ;
        RECT 555.750 15.060 558.830 15.200 ;
        RECT 555.750 15.000 556.070 15.060 ;
        RECT 558.510 15.000 558.830 15.060 ;
      LAYER via ;
        RECT 558.540 1084.640 558.800 1084.900 ;
        RECT 1040.620 1084.640 1040.880 1084.900 ;
        RECT 555.780 15.000 556.040 15.260 ;
        RECT 558.540 15.000 558.800 15.260 ;
      LAYER met2 ;
        RECT 1040.530 1100.580 1040.810 1104.000 ;
        RECT 1040.530 1100.000 1040.820 1100.580 ;
        RECT 1040.680 1084.930 1040.820 1100.000 ;
        RECT 558.540 1084.610 558.800 1084.930 ;
        RECT 1040.620 1084.610 1040.880 1084.930 ;
        RECT 558.600 15.290 558.740 1084.610 ;
        RECT 555.780 14.970 556.040 15.290 ;
        RECT 558.540 14.970 558.800 15.290 ;
        RECT 555.840 2.000 555.980 14.970 ;
        RECT 555.630 -4.000 556.190 2.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 607.345 14.365 608.435 14.535 ;
      LAYER mcon ;
        RECT 608.265 14.365 608.435 14.535 ;
      LAYER met1 ;
        RECT 977.110 1088.240 977.430 1088.300 ;
        RECT 1046.570 1088.240 1046.890 1088.300 ;
        RECT 977.110 1088.100 1046.890 1088.240 ;
        RECT 977.110 1088.040 977.430 1088.100 ;
        RECT 1046.570 1088.040 1046.890 1088.100 ;
        RECT 573.690 14.520 574.010 14.580 ;
        RECT 607.285 14.520 607.575 14.565 ;
        RECT 573.690 14.380 607.575 14.520 ;
        RECT 573.690 14.320 574.010 14.380 ;
        RECT 607.285 14.335 607.575 14.380 ;
        RECT 608.205 14.520 608.495 14.565 ;
        RECT 977.110 14.520 977.430 14.580 ;
        RECT 608.205 14.380 977.430 14.520 ;
        RECT 608.205 14.335 608.495 14.380 ;
        RECT 977.110 14.320 977.430 14.380 ;
      LAYER via ;
        RECT 977.140 1088.040 977.400 1088.300 ;
        RECT 1046.600 1088.040 1046.860 1088.300 ;
        RECT 573.720 14.320 573.980 14.580 ;
        RECT 977.140 14.320 977.400 14.580 ;
      LAYER met2 ;
        RECT 1046.510 1100.580 1046.790 1104.000 ;
        RECT 1046.510 1100.000 1046.800 1100.580 ;
        RECT 1046.660 1088.330 1046.800 1100.000 ;
        RECT 977.140 1088.010 977.400 1088.330 ;
        RECT 1046.600 1088.010 1046.860 1088.330 ;
        RECT 977.200 14.610 977.340 1088.010 ;
        RECT 573.720 14.290 573.980 14.610 ;
        RECT 977.140 14.290 977.400 14.610 ;
        RECT 573.780 2.000 573.920 14.290 ;
        RECT 573.570 -4.000 574.130 2.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 593.010 1084.500 593.330 1084.560 ;
        RECT 1053.010 1084.500 1053.330 1084.560 ;
        RECT 593.010 1084.360 1053.330 1084.500 ;
        RECT 593.010 1084.300 593.330 1084.360 ;
        RECT 1053.010 1084.300 1053.330 1084.360 ;
      LAYER via ;
        RECT 593.040 1084.300 593.300 1084.560 ;
        RECT 1053.040 1084.300 1053.300 1084.560 ;
      LAYER met2 ;
        RECT 1052.950 1100.580 1053.230 1104.000 ;
        RECT 1052.950 1100.000 1053.240 1100.580 ;
        RECT 1053.100 1084.590 1053.240 1100.000 ;
        RECT 593.040 1084.270 593.300 1084.590 ;
        RECT 1053.040 1084.270 1053.300 1084.590 ;
        RECT 593.100 2.450 593.240 1084.270 ;
        RECT 591.260 2.310 593.240 2.450 ;
        RECT 591.260 2.000 591.400 2.310 ;
        RECT 591.050 -4.000 591.610 2.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 97.590 17.920 97.910 17.980 ;
        RECT 883.270 17.920 883.590 17.980 ;
        RECT 97.590 17.780 883.590 17.920 ;
        RECT 97.590 17.720 97.910 17.780 ;
        RECT 883.270 17.720 883.590 17.780 ;
      LAYER via ;
        RECT 97.620 17.720 97.880 17.980 ;
        RECT 883.300 17.720 883.560 17.980 ;
      LAYER met2 ;
        RECT 883.210 1100.580 883.490 1104.000 ;
        RECT 883.210 1100.000 883.500 1100.580 ;
        RECT 883.360 18.010 883.500 1100.000 ;
        RECT 97.620 17.690 97.880 18.010 ;
        RECT 883.300 17.690 883.560 18.010 ;
        RECT 97.680 2.000 97.820 17.690 ;
        RECT 97.470 -4.000 98.030 2.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 613.710 1084.160 614.030 1084.220 ;
        RECT 1057.610 1084.160 1057.930 1084.220 ;
        RECT 613.710 1084.020 1057.930 1084.160 ;
        RECT 613.710 1083.960 614.030 1084.020 ;
        RECT 1057.610 1083.960 1057.930 1084.020 ;
        RECT 609.110 14.180 609.430 14.240 ;
        RECT 613.710 14.180 614.030 14.240 ;
        RECT 609.110 14.040 614.030 14.180 ;
        RECT 609.110 13.980 609.430 14.040 ;
        RECT 613.710 13.980 614.030 14.040 ;
      LAYER via ;
        RECT 613.740 1083.960 614.000 1084.220 ;
        RECT 1057.640 1083.960 1057.900 1084.220 ;
        RECT 609.140 13.980 609.400 14.240 ;
        RECT 613.740 13.980 614.000 14.240 ;
      LAYER met2 ;
        RECT 1058.930 1100.650 1059.210 1104.000 ;
        RECT 1057.700 1100.510 1059.210 1100.650 ;
        RECT 1057.700 1084.250 1057.840 1100.510 ;
        RECT 1058.930 1100.000 1059.210 1100.510 ;
        RECT 613.740 1083.930 614.000 1084.250 ;
        RECT 1057.640 1083.930 1057.900 1084.250 ;
        RECT 613.800 14.270 613.940 1083.930 ;
        RECT 609.140 13.950 609.400 14.270 ;
        RECT 613.740 13.950 614.000 14.270 ;
        RECT 609.200 2.000 609.340 13.950 ;
        RECT 608.990 -4.000 609.550 2.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 983.090 1089.600 983.410 1089.660 ;
        RECT 1064.970 1089.600 1065.290 1089.660 ;
        RECT 983.090 1089.460 1065.290 1089.600 ;
        RECT 983.090 1089.400 983.410 1089.460 ;
        RECT 1064.970 1089.400 1065.290 1089.460 ;
        RECT 983.090 14.180 983.410 14.240 ;
        RECT 628.060 14.040 983.410 14.180 ;
        RECT 627.050 13.840 627.370 13.900 ;
        RECT 628.060 13.840 628.200 14.040 ;
        RECT 983.090 13.980 983.410 14.040 ;
        RECT 627.050 13.700 628.200 13.840 ;
        RECT 627.050 13.640 627.370 13.700 ;
      LAYER via ;
        RECT 983.120 1089.400 983.380 1089.660 ;
        RECT 1065.000 1089.400 1065.260 1089.660 ;
        RECT 627.080 13.640 627.340 13.900 ;
        RECT 983.120 13.980 983.380 14.240 ;
      LAYER met2 ;
        RECT 1064.910 1100.580 1065.190 1104.000 ;
        RECT 1064.910 1100.000 1065.200 1100.580 ;
        RECT 1065.060 1089.690 1065.200 1100.000 ;
        RECT 983.120 1089.370 983.380 1089.690 ;
        RECT 1065.000 1089.370 1065.260 1089.690 ;
        RECT 983.180 14.270 983.320 1089.370 ;
        RECT 983.120 13.950 983.380 14.270 ;
        RECT 627.080 13.610 627.340 13.930 ;
        RECT 627.140 2.000 627.280 13.610 ;
        RECT 626.930 -4.000 627.490 2.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 835.505 1086.555 835.675 1086.895 ;
        RECT 835.505 1086.385 836.595 1086.555 ;
      LAYER mcon ;
        RECT 835.505 1086.725 835.675 1086.895 ;
        RECT 836.425 1086.385 836.595 1086.555 ;
      LAYER met1 ;
        RECT 155.090 1087.220 155.410 1087.280 ;
        RECT 155.090 1087.080 835.660 1087.220 ;
        RECT 155.090 1087.020 155.410 1087.080 ;
        RECT 835.520 1086.925 835.660 1087.080 ;
        RECT 835.445 1086.695 835.735 1086.925 ;
        RECT 836.365 1086.540 836.655 1086.585 ;
        RECT 891.550 1086.540 891.870 1086.600 ;
        RECT 836.365 1086.400 891.870 1086.540 ;
        RECT 836.365 1086.355 836.655 1086.400 ;
        RECT 891.550 1086.340 891.870 1086.400 ;
        RECT 121.510 19.280 121.830 19.340 ;
        RECT 155.090 19.280 155.410 19.340 ;
        RECT 121.510 19.140 155.410 19.280 ;
        RECT 121.510 19.080 121.830 19.140 ;
        RECT 155.090 19.080 155.410 19.140 ;
      LAYER via ;
        RECT 155.120 1087.020 155.380 1087.280 ;
        RECT 891.580 1086.340 891.840 1086.600 ;
        RECT 121.540 19.080 121.800 19.340 ;
        RECT 155.120 19.080 155.380 19.340 ;
      LAYER met2 ;
        RECT 891.490 1100.580 891.770 1104.000 ;
        RECT 891.490 1100.000 891.780 1100.580 ;
        RECT 155.120 1086.990 155.380 1087.310 ;
        RECT 155.180 19.370 155.320 1086.990 ;
        RECT 891.640 1086.630 891.780 1100.000 ;
        RECT 891.580 1086.310 891.840 1086.630 ;
        RECT 121.540 19.050 121.800 19.370 ;
        RECT 155.120 19.050 155.380 19.370 ;
        RECT 121.600 2.000 121.740 19.050 ;
        RECT 121.390 -4.000 121.950 2.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 897.070 1069.200 897.390 1069.260 ;
        RECT 899.830 1069.200 900.150 1069.260 ;
        RECT 897.070 1069.060 900.150 1069.200 ;
        RECT 897.070 1069.000 897.390 1069.060 ;
        RECT 899.830 1069.000 900.150 1069.060 ;
        RECT 145.430 18.600 145.750 18.660 ;
        RECT 897.070 18.600 897.390 18.660 ;
        RECT 145.430 18.460 897.390 18.600 ;
        RECT 145.430 18.400 145.750 18.460 ;
        RECT 897.070 18.400 897.390 18.460 ;
      LAYER via ;
        RECT 897.100 1069.000 897.360 1069.260 ;
        RECT 899.860 1069.000 900.120 1069.260 ;
        RECT 145.460 18.400 145.720 18.660 ;
        RECT 897.100 18.400 897.360 18.660 ;
      LAYER met2 ;
        RECT 899.770 1100.580 900.050 1104.000 ;
        RECT 899.770 1100.000 900.060 1100.580 ;
        RECT 899.920 1069.290 900.060 1100.000 ;
        RECT 897.100 1068.970 897.360 1069.290 ;
        RECT 899.860 1068.970 900.120 1069.290 ;
        RECT 897.160 18.690 897.300 1068.970 ;
        RECT 145.460 18.370 145.720 18.690 ;
        RECT 897.100 18.370 897.360 18.690 ;
        RECT 145.520 2.000 145.660 18.370 ;
        RECT 145.310 -4.000 145.870 2.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 175.790 1087.900 176.110 1087.960 ;
        RECT 905.810 1087.900 906.130 1087.960 ;
        RECT 175.790 1087.760 906.130 1087.900 ;
        RECT 175.790 1087.700 176.110 1087.760 ;
        RECT 905.810 1087.700 906.130 1087.760 ;
        RECT 163.370 16.900 163.690 16.960 ;
        RECT 175.790 16.900 176.110 16.960 ;
        RECT 163.370 16.760 176.110 16.900 ;
        RECT 163.370 16.700 163.690 16.760 ;
        RECT 175.790 16.700 176.110 16.760 ;
      LAYER via ;
        RECT 175.820 1087.700 176.080 1087.960 ;
        RECT 905.840 1087.700 906.100 1087.960 ;
        RECT 163.400 16.700 163.660 16.960 ;
        RECT 175.820 16.700 176.080 16.960 ;
      LAYER met2 ;
        RECT 905.750 1100.580 906.030 1104.000 ;
        RECT 905.750 1100.000 906.040 1100.580 ;
        RECT 905.900 1087.990 906.040 1100.000 ;
        RECT 175.820 1087.670 176.080 1087.990 ;
        RECT 905.840 1087.670 906.100 1087.990 ;
        RECT 175.880 16.990 176.020 1087.670 ;
        RECT 163.400 16.670 163.660 16.990 ;
        RECT 175.820 16.670 176.080 16.990 ;
        RECT 163.460 2.000 163.600 16.670 ;
        RECT 163.250 -4.000 163.810 2.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 911.865 88.825 912.035 90.015 ;
      LAYER mcon ;
        RECT 911.865 89.845 912.035 90.015 ;
      LAYER met1 ;
        RECT 911.790 385.940 912.110 386.200 ;
        RECT 911.880 385.520 912.020 385.940 ;
        RECT 911.790 385.260 912.110 385.520 ;
        RECT 911.790 90.000 912.110 90.060 ;
        RECT 911.595 89.860 912.110 90.000 ;
        RECT 911.790 89.800 912.110 89.860 ;
        RECT 911.790 88.980 912.110 89.040 ;
        RECT 911.595 88.840 912.110 88.980 ;
        RECT 911.790 88.780 912.110 88.840 ;
        RECT 180.850 19.280 181.170 19.340 ;
        RECT 911.790 19.280 912.110 19.340 ;
        RECT 180.850 19.140 912.110 19.280 ;
        RECT 180.850 19.080 181.170 19.140 ;
        RECT 911.790 19.080 912.110 19.140 ;
      LAYER via ;
        RECT 911.820 385.940 912.080 386.200 ;
        RECT 911.820 385.260 912.080 385.520 ;
        RECT 911.820 89.800 912.080 90.060 ;
        RECT 911.820 88.780 912.080 89.040 ;
        RECT 180.880 19.080 181.140 19.340 ;
        RECT 911.820 19.080 912.080 19.340 ;
      LAYER met2 ;
        RECT 912.190 1100.650 912.470 1104.000 ;
        RECT 911.880 1100.510 912.470 1100.650 ;
        RECT 911.880 386.230 912.020 1100.510 ;
        RECT 912.190 1100.000 912.470 1100.510 ;
        RECT 911.820 385.910 912.080 386.230 ;
        RECT 911.820 385.230 912.080 385.550 ;
        RECT 911.880 90.090 912.020 385.230 ;
        RECT 911.820 89.770 912.080 90.090 ;
        RECT 911.820 88.750 912.080 89.070 ;
        RECT 911.880 19.370 912.020 88.750 ;
        RECT 180.880 19.050 181.140 19.370 ;
        RECT 911.820 19.050 912.080 19.370 ;
        RECT 180.940 2.000 181.080 19.050 ;
        RECT 180.730 -4.000 181.290 2.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 210.290 1088.240 210.610 1088.300 ;
        RECT 918.230 1088.240 918.550 1088.300 ;
        RECT 210.290 1088.100 918.550 1088.240 ;
        RECT 210.290 1088.040 210.610 1088.100 ;
        RECT 918.230 1088.040 918.550 1088.100 ;
        RECT 198.790 16.900 199.110 16.960 ;
        RECT 210.290 16.900 210.610 16.960 ;
        RECT 198.790 16.760 210.610 16.900 ;
        RECT 198.790 16.700 199.110 16.760 ;
        RECT 210.290 16.700 210.610 16.760 ;
      LAYER via ;
        RECT 210.320 1088.040 210.580 1088.300 ;
        RECT 918.260 1088.040 918.520 1088.300 ;
        RECT 198.820 16.700 199.080 16.960 ;
        RECT 210.320 16.700 210.580 16.960 ;
      LAYER met2 ;
        RECT 918.170 1100.580 918.450 1104.000 ;
        RECT 918.170 1100.000 918.460 1100.580 ;
        RECT 918.320 1088.330 918.460 1100.000 ;
        RECT 210.320 1088.010 210.580 1088.330 ;
        RECT 918.260 1088.010 918.520 1088.330 ;
        RECT 210.380 16.990 210.520 1088.010 ;
        RECT 198.820 16.670 199.080 16.990 ;
        RECT 210.320 16.670 210.580 16.990 ;
        RECT 198.880 2.000 199.020 16.670 ;
        RECT 198.670 -4.000 199.230 2.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 919.150 1042.000 919.470 1042.060 ;
        RECT 922.830 1042.000 923.150 1042.060 ;
        RECT 919.150 1041.860 923.150 1042.000 ;
        RECT 919.150 1041.800 919.470 1041.860 ;
        RECT 922.830 1041.800 923.150 1041.860 ;
        RECT 216.730 19.960 217.050 20.020 ;
        RECT 919.150 19.960 919.470 20.020 ;
        RECT 216.730 19.820 919.470 19.960 ;
        RECT 216.730 19.760 217.050 19.820 ;
        RECT 919.150 19.760 919.470 19.820 ;
      LAYER via ;
        RECT 919.180 1041.800 919.440 1042.060 ;
        RECT 922.860 1041.800 923.120 1042.060 ;
        RECT 216.760 19.760 217.020 20.020 ;
        RECT 919.180 19.760 919.440 20.020 ;
      LAYER met2 ;
        RECT 924.150 1100.650 924.430 1104.000 ;
        RECT 922.920 1100.510 924.430 1100.650 ;
        RECT 922.920 1042.090 923.060 1100.510 ;
        RECT 924.150 1100.000 924.430 1100.510 ;
        RECT 919.180 1041.770 919.440 1042.090 ;
        RECT 922.860 1041.770 923.120 1042.090 ;
        RECT 919.240 20.050 919.380 1041.770 ;
        RECT 216.760 19.730 217.020 20.050 ;
        RECT 919.180 19.730 919.440 20.050 ;
        RECT 216.820 2.000 216.960 19.730 ;
        RECT 216.610 -4.000 217.170 2.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 324.445 14.025 324.615 14.875 ;
        RECT 348.825 13.685 348.995 15.215 ;
        RECT 372.745 15.045 372.915 16.575 ;
        RECT 388.845 15.555 389.015 16.575 ;
        RECT 388.845 15.385 390.395 15.555 ;
        RECT 394.825 15.385 394.995 16.575 ;
        RECT 406.785 13.685 406.955 16.575 ;
        RECT 420.585 13.685 420.755 15.215 ;
        RECT 477.625 14.025 477.795 15.215 ;
      LAYER mcon ;
        RECT 372.745 16.405 372.915 16.575 ;
        RECT 388.845 16.405 389.015 16.575 ;
        RECT 394.825 16.405 394.995 16.575 ;
        RECT 390.225 15.385 390.395 15.555 ;
        RECT 406.785 16.405 406.955 16.575 ;
        RECT 348.825 15.045 348.995 15.215 ;
        RECT 324.445 14.705 324.615 14.875 ;
        RECT 420.585 15.045 420.755 15.215 ;
        RECT 477.625 15.045 477.795 15.215 ;
      LAYER met1 ;
        RECT 486.290 1083.820 486.610 1083.880 ;
        RECT 930.650 1083.820 930.970 1083.880 ;
        RECT 486.290 1083.680 930.970 1083.820 ;
        RECT 486.290 1083.620 486.610 1083.680 ;
        RECT 930.650 1083.620 930.970 1083.680 ;
        RECT 372.685 16.560 372.975 16.605 ;
        RECT 388.785 16.560 389.075 16.605 ;
        RECT 372.685 16.420 389.075 16.560 ;
        RECT 372.685 16.375 372.975 16.420 ;
        RECT 388.785 16.375 389.075 16.420 ;
        RECT 394.765 16.560 395.055 16.605 ;
        RECT 406.725 16.560 407.015 16.605 ;
        RECT 394.765 16.420 407.015 16.560 ;
        RECT 394.765 16.375 395.055 16.420 ;
        RECT 406.725 16.375 407.015 16.420 ;
        RECT 390.165 15.540 390.455 15.585 ;
        RECT 394.765 15.540 395.055 15.585 ;
        RECT 390.165 15.400 395.055 15.540 ;
        RECT 390.165 15.355 390.455 15.400 ;
        RECT 394.765 15.355 395.055 15.400 ;
        RECT 348.765 15.200 349.055 15.245 ;
        RECT 372.685 15.200 372.975 15.245 ;
        RECT 348.765 15.060 372.975 15.200 ;
        RECT 348.765 15.015 349.055 15.060 ;
        RECT 372.685 15.015 372.975 15.060 ;
        RECT 420.525 15.200 420.815 15.245 ;
        RECT 477.565 15.200 477.855 15.245 ;
        RECT 420.525 15.060 477.855 15.200 ;
        RECT 420.525 15.015 420.815 15.060 ;
        RECT 477.565 15.015 477.855 15.060 ;
        RECT 234.670 14.860 234.990 14.920 ;
        RECT 324.385 14.860 324.675 14.905 ;
        RECT 234.670 14.720 324.675 14.860 ;
        RECT 234.670 14.660 234.990 14.720 ;
        RECT 324.385 14.675 324.675 14.720 ;
        RECT 324.385 14.180 324.675 14.225 ;
        RECT 477.565 14.180 477.855 14.225 ;
        RECT 486.290 14.180 486.610 14.240 ;
        RECT 324.385 14.040 348.060 14.180 ;
        RECT 324.385 13.995 324.675 14.040 ;
        RECT 347.920 13.840 348.060 14.040 ;
        RECT 477.565 14.040 486.610 14.180 ;
        RECT 477.565 13.995 477.855 14.040 ;
        RECT 486.290 13.980 486.610 14.040 ;
        RECT 348.765 13.840 349.055 13.885 ;
        RECT 347.920 13.700 349.055 13.840 ;
        RECT 348.765 13.655 349.055 13.700 ;
        RECT 406.725 13.840 407.015 13.885 ;
        RECT 420.525 13.840 420.815 13.885 ;
        RECT 406.725 13.700 420.815 13.840 ;
        RECT 406.725 13.655 407.015 13.700 ;
        RECT 420.525 13.655 420.815 13.700 ;
      LAYER via ;
        RECT 486.320 1083.620 486.580 1083.880 ;
        RECT 930.680 1083.620 930.940 1083.880 ;
        RECT 234.700 14.660 234.960 14.920 ;
        RECT 486.320 13.980 486.580 14.240 ;
      LAYER met2 ;
        RECT 930.590 1100.580 930.870 1104.000 ;
        RECT 930.590 1100.000 930.880 1100.580 ;
        RECT 930.740 1083.910 930.880 1100.000 ;
        RECT 486.320 1083.590 486.580 1083.910 ;
        RECT 930.680 1083.590 930.940 1083.910 ;
        RECT 234.700 14.630 234.960 14.950 ;
        RECT 234.760 2.000 234.900 14.630 ;
        RECT 486.380 14.270 486.520 1083.590 ;
        RECT 486.320 13.950 486.580 14.270 ;
        RECT 234.550 -4.000 235.110 2.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 865.405 579.785 865.575 627.895 ;
        RECT 865.405 483.225 865.575 531.335 ;
        RECT 865.405 386.325 865.575 434.775 ;
        RECT 865.405 289.765 865.575 337.875 ;
      LAYER mcon ;
        RECT 865.405 627.725 865.575 627.895 ;
        RECT 865.405 531.165 865.575 531.335 ;
        RECT 865.405 434.605 865.575 434.775 ;
        RECT 865.405 337.705 865.575 337.875 ;
      LAYER met1 ;
        RECT 866.250 1062.740 866.570 1062.800 ;
        RECT 869.010 1062.740 869.330 1062.800 ;
        RECT 866.250 1062.600 869.330 1062.740 ;
        RECT 866.250 1062.540 866.570 1062.600 ;
        RECT 869.010 1062.540 869.330 1062.600 ;
        RECT 866.710 1014.460 867.030 1014.520 ;
        RECT 867.170 1014.460 867.490 1014.520 ;
        RECT 866.710 1014.320 867.490 1014.460 ;
        RECT 866.710 1014.260 867.030 1014.320 ;
        RECT 867.170 1014.260 867.490 1014.320 ;
        RECT 865.790 966.180 866.110 966.240 ;
        RECT 867.630 966.180 867.950 966.240 ;
        RECT 865.790 966.040 867.950 966.180 ;
        RECT 865.790 965.980 866.110 966.040 ;
        RECT 867.630 965.980 867.950 966.040 ;
        RECT 865.330 869.620 865.650 869.680 ;
        RECT 865.790 869.620 866.110 869.680 ;
        RECT 865.330 869.480 866.110 869.620 ;
        RECT 865.330 869.420 865.650 869.480 ;
        RECT 865.790 869.420 866.110 869.480 ;
        RECT 865.330 821.000 865.650 821.060 ;
        RECT 866.250 821.000 866.570 821.060 ;
        RECT 865.330 820.860 866.570 821.000 ;
        RECT 865.330 820.800 865.650 820.860 ;
        RECT 866.250 820.800 866.570 820.860 ;
        RECT 865.330 724.440 865.650 724.500 ;
        RECT 866.250 724.440 866.570 724.500 ;
        RECT 865.330 724.300 866.570 724.440 ;
        RECT 865.330 724.240 865.650 724.300 ;
        RECT 866.250 724.240 866.570 724.300 ;
        RECT 865.330 627.880 865.650 627.940 ;
        RECT 865.135 627.740 865.650 627.880 ;
        RECT 865.330 627.680 865.650 627.740 ;
        RECT 865.330 579.940 865.650 580.000 ;
        RECT 865.135 579.800 865.650 579.940 ;
        RECT 865.330 579.740 865.650 579.800 ;
        RECT 865.330 531.320 865.650 531.380 ;
        RECT 865.135 531.180 865.650 531.320 ;
        RECT 865.330 531.120 865.650 531.180 ;
        RECT 865.330 483.380 865.650 483.440 ;
        RECT 865.135 483.240 865.650 483.380 ;
        RECT 865.330 483.180 865.650 483.240 ;
        RECT 865.330 434.760 865.650 434.820 ;
        RECT 865.135 434.620 865.650 434.760 ;
        RECT 865.330 434.560 865.650 434.620 ;
        RECT 865.330 386.480 865.650 386.540 ;
        RECT 865.135 386.340 865.650 386.480 ;
        RECT 865.330 386.280 865.650 386.340 ;
        RECT 865.330 337.860 865.650 337.920 ;
        RECT 865.135 337.720 865.650 337.860 ;
        RECT 865.330 337.660 865.650 337.720 ;
        RECT 865.330 289.920 865.650 289.980 ;
        RECT 865.135 289.780 865.650 289.920 ;
        RECT 865.330 289.720 865.650 289.780 ;
        RECT 865.330 144.740 865.650 144.800 ;
        RECT 865.790 144.740 866.110 144.800 ;
        RECT 865.330 144.600 866.110 144.740 ;
        RECT 865.330 144.540 865.650 144.600 ;
        RECT 865.790 144.540 866.110 144.600 ;
        RECT 56.190 17.580 56.510 17.640 ;
        RECT 865.790 17.580 866.110 17.640 ;
        RECT 56.190 17.440 866.110 17.580 ;
        RECT 56.190 17.380 56.510 17.440 ;
        RECT 865.790 17.380 866.110 17.440 ;
      LAYER via ;
        RECT 866.280 1062.540 866.540 1062.800 ;
        RECT 869.040 1062.540 869.300 1062.800 ;
        RECT 866.740 1014.260 867.000 1014.520 ;
        RECT 867.200 1014.260 867.460 1014.520 ;
        RECT 865.820 965.980 866.080 966.240 ;
        RECT 867.660 965.980 867.920 966.240 ;
        RECT 865.360 869.420 865.620 869.680 ;
        RECT 865.820 869.420 866.080 869.680 ;
        RECT 865.360 820.800 865.620 821.060 ;
        RECT 866.280 820.800 866.540 821.060 ;
        RECT 865.360 724.240 865.620 724.500 ;
        RECT 866.280 724.240 866.540 724.500 ;
        RECT 865.360 627.680 865.620 627.940 ;
        RECT 865.360 579.740 865.620 580.000 ;
        RECT 865.360 531.120 865.620 531.380 ;
        RECT 865.360 483.180 865.620 483.440 ;
        RECT 865.360 434.560 865.620 434.820 ;
        RECT 865.360 386.280 865.620 386.540 ;
        RECT 865.360 337.660 865.620 337.920 ;
        RECT 865.360 289.720 865.620 289.980 ;
        RECT 865.360 144.540 865.620 144.800 ;
        RECT 865.820 144.540 866.080 144.800 ;
        RECT 56.220 17.380 56.480 17.640 ;
        RECT 865.820 17.380 866.080 17.640 ;
      LAYER met2 ;
        RECT 868.950 1100.580 869.230 1104.000 ;
        RECT 868.950 1100.000 869.240 1100.580 ;
        RECT 869.100 1062.830 869.240 1100.000 ;
        RECT 866.280 1062.685 866.540 1062.830 ;
        RECT 866.270 1062.315 866.550 1062.685 ;
        RECT 867.190 1062.315 867.470 1062.685 ;
        RECT 869.040 1062.510 869.300 1062.830 ;
        RECT 866.800 1014.550 866.940 1014.705 ;
        RECT 867.260 1014.550 867.400 1062.315 ;
        RECT 866.740 1014.290 867.000 1014.550 ;
        RECT 867.200 1014.290 867.460 1014.550 ;
        RECT 866.740 1014.230 867.860 1014.290 ;
        RECT 866.800 1014.150 867.860 1014.230 ;
        RECT 867.720 966.270 867.860 1014.150 ;
        RECT 865.820 965.950 866.080 966.270 ;
        RECT 867.660 965.950 867.920 966.270 ;
        RECT 865.880 869.710 866.020 965.950 ;
        RECT 865.360 869.390 865.620 869.710 ;
        RECT 865.820 869.390 866.080 869.710 ;
        RECT 865.420 821.090 865.560 869.390 ;
        RECT 865.360 820.770 865.620 821.090 ;
        RECT 866.280 820.770 866.540 821.090 ;
        RECT 866.340 773.005 866.480 820.770 ;
        RECT 865.350 772.635 865.630 773.005 ;
        RECT 866.270 772.635 866.550 773.005 ;
        RECT 865.420 724.530 865.560 772.635 ;
        RECT 865.360 724.210 865.620 724.530 ;
        RECT 866.280 724.210 866.540 724.530 ;
        RECT 866.340 676.445 866.480 724.210 ;
        RECT 865.350 676.075 865.630 676.445 ;
        RECT 866.270 676.075 866.550 676.445 ;
        RECT 865.420 627.970 865.560 676.075 ;
        RECT 865.360 627.650 865.620 627.970 ;
        RECT 865.360 579.710 865.620 580.030 ;
        RECT 865.420 531.410 865.560 579.710 ;
        RECT 865.360 531.090 865.620 531.410 ;
        RECT 865.360 483.150 865.620 483.470 ;
        RECT 865.420 434.850 865.560 483.150 ;
        RECT 865.360 434.530 865.620 434.850 ;
        RECT 865.360 386.250 865.620 386.570 ;
        RECT 865.420 337.950 865.560 386.250 ;
        RECT 865.360 337.630 865.620 337.950 ;
        RECT 865.360 289.690 865.620 290.010 ;
        RECT 865.420 144.830 865.560 289.690 ;
        RECT 865.360 144.510 865.620 144.830 ;
        RECT 865.820 144.510 866.080 144.830 ;
        RECT 865.880 17.670 866.020 144.510 ;
        RECT 56.220 17.350 56.480 17.670 ;
        RECT 865.820 17.350 866.080 17.670 ;
        RECT 56.280 2.000 56.420 17.350 ;
        RECT 56.070 -4.000 56.630 2.000 ;
      LAYER via2 ;
        RECT 866.270 1062.360 866.550 1062.640 ;
        RECT 867.190 1062.360 867.470 1062.640 ;
        RECT 865.350 772.680 865.630 772.960 ;
        RECT 866.270 772.680 866.550 772.960 ;
        RECT 865.350 676.120 865.630 676.400 ;
        RECT 866.270 676.120 866.550 676.400 ;
      LAYER met3 ;
        RECT 866.245 1062.650 866.575 1062.665 ;
        RECT 867.165 1062.650 867.495 1062.665 ;
        RECT 866.245 1062.350 867.495 1062.650 ;
        RECT 866.245 1062.335 866.575 1062.350 ;
        RECT 867.165 1062.335 867.495 1062.350 ;
        RECT 865.325 772.970 865.655 772.985 ;
        RECT 866.245 772.970 866.575 772.985 ;
        RECT 865.325 772.670 866.575 772.970 ;
        RECT 865.325 772.655 865.655 772.670 ;
        RECT 866.245 772.655 866.575 772.670 ;
        RECT 865.325 676.410 865.655 676.425 ;
        RECT 866.245 676.410 866.575 676.425 ;
        RECT 865.325 676.110 866.575 676.410 ;
        RECT 865.325 676.095 865.655 676.110 ;
        RECT 866.245 676.095 866.575 676.110 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 853.905 1087.235 854.075 1087.575 ;
        RECT 854.825 1087.235 854.995 1088.595 ;
        RECT 835.045 1087.065 836.135 1087.235 ;
        RECT 853.905 1087.065 854.995 1087.235 ;
        RECT 835.045 1086.725 835.215 1087.065 ;
      LAYER mcon ;
        RECT 854.825 1088.425 854.995 1088.595 ;
        RECT 853.905 1087.405 854.075 1087.575 ;
        RECT 835.965 1087.065 836.135 1087.235 ;
      LAYER met1 ;
        RECT 854.765 1088.580 855.055 1088.625 ;
        RECT 877.290 1088.580 877.610 1088.640 ;
        RECT 854.765 1088.440 877.610 1088.580 ;
        RECT 854.765 1088.395 855.055 1088.440 ;
        RECT 877.290 1088.380 877.610 1088.440 ;
        RECT 853.845 1087.560 854.135 1087.605 ;
        RECT 841.960 1087.420 854.135 1087.560 ;
        RECT 835.905 1087.220 836.195 1087.265 ;
        RECT 841.960 1087.220 842.100 1087.420 ;
        RECT 853.845 1087.375 854.135 1087.420 ;
        RECT 835.905 1087.080 842.100 1087.220 ;
        RECT 835.905 1087.035 836.195 1087.080 ;
        RECT 120.590 1086.880 120.910 1086.940 ;
        RECT 834.985 1086.880 835.275 1086.925 ;
        RECT 120.590 1086.740 835.275 1086.880 ;
        RECT 120.590 1086.680 120.910 1086.740 ;
        RECT 834.985 1086.695 835.275 1086.740 ;
        RECT 80.110 18.600 80.430 18.660 ;
        RECT 120.590 18.600 120.910 18.660 ;
        RECT 80.110 18.460 120.910 18.600 ;
        RECT 80.110 18.400 80.430 18.460 ;
        RECT 120.590 18.400 120.910 18.460 ;
      LAYER via ;
        RECT 877.320 1088.380 877.580 1088.640 ;
        RECT 120.620 1086.680 120.880 1086.940 ;
        RECT 80.140 18.400 80.400 18.660 ;
        RECT 120.620 18.400 120.880 18.660 ;
      LAYER met2 ;
        RECT 877.230 1100.580 877.510 1104.000 ;
        RECT 877.230 1100.000 877.520 1100.580 ;
        RECT 877.380 1088.670 877.520 1100.000 ;
        RECT 877.320 1088.350 877.580 1088.670 ;
        RECT 120.620 1086.650 120.880 1086.970 ;
        RECT 120.680 18.690 120.820 1086.650 ;
        RECT 80.140 18.370 80.400 18.690 ;
        RECT 120.620 18.370 120.880 18.690 ;
        RECT 80.200 2.000 80.340 18.370 ;
        RECT 79.990 -4.000 80.550 2.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 103.570 18.260 103.890 18.320 ;
        RECT 883.730 18.260 884.050 18.320 ;
        RECT 103.570 18.120 884.050 18.260 ;
        RECT 103.570 18.060 103.890 18.120 ;
        RECT 883.730 18.060 884.050 18.120 ;
      LAYER via ;
        RECT 103.600 18.060 103.860 18.320 ;
        RECT 883.760 18.060 884.020 18.320 ;
      LAYER met2 ;
        RECT 885.510 1100.650 885.790 1104.000 ;
        RECT 883.820 1100.510 885.790 1100.650 ;
        RECT 883.820 18.350 883.960 1100.510 ;
        RECT 885.510 1100.000 885.790 1100.510 ;
        RECT 103.600 18.030 103.860 18.350 ;
        RECT 883.760 18.030 884.020 18.350 ;
        RECT 103.660 2.000 103.800 18.030 ;
        RECT 103.450 -4.000 104.010 2.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 841.485 1087.235 841.655 1087.575 ;
        RECT 841.485 1087.065 842.575 1087.235 ;
      LAYER mcon ;
        RECT 841.485 1087.405 841.655 1087.575 ;
        RECT 842.405 1087.065 842.575 1087.235 ;
      LAYER met1 ;
        RECT 161.990 1087.560 162.310 1087.620 ;
        RECT 841.425 1087.560 841.715 1087.605 ;
        RECT 161.990 1087.420 841.715 1087.560 ;
        RECT 161.990 1087.360 162.310 1087.420 ;
        RECT 841.425 1087.375 841.715 1087.420 ;
        RECT 842.345 1087.220 842.635 1087.265 ;
        RECT 893.850 1087.220 894.170 1087.280 ;
        RECT 842.345 1087.080 894.170 1087.220 ;
        RECT 842.345 1087.035 842.635 1087.080 ;
        RECT 893.850 1087.020 894.170 1087.080 ;
        RECT 127.490 18.940 127.810 19.000 ;
        RECT 161.990 18.940 162.310 19.000 ;
        RECT 127.490 18.800 162.310 18.940 ;
        RECT 127.490 18.740 127.810 18.800 ;
        RECT 161.990 18.740 162.310 18.800 ;
      LAYER via ;
        RECT 162.020 1087.360 162.280 1087.620 ;
        RECT 893.880 1087.020 894.140 1087.280 ;
        RECT 127.520 18.740 127.780 19.000 ;
        RECT 162.020 18.740 162.280 19.000 ;
      LAYER met2 ;
        RECT 893.790 1100.580 894.070 1104.000 ;
        RECT 893.790 1100.000 894.080 1100.580 ;
        RECT 162.020 1087.330 162.280 1087.650 ;
        RECT 162.080 19.030 162.220 1087.330 ;
        RECT 893.940 1087.310 894.080 1100.000 ;
        RECT 893.880 1086.990 894.140 1087.310 ;
        RECT 127.520 18.710 127.780 19.030 ;
        RECT 162.020 18.710 162.280 19.030 ;
        RECT 127.580 2.000 127.720 18.710 ;
        RECT 127.370 -4.000 127.930 2.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 857.585 966.025 857.755 980.135 ;
        RECT 857.125 579.785 857.295 627.895 ;
        RECT 857.125 483.225 857.295 531.335 ;
        RECT 857.125 386.325 857.295 434.775 ;
        RECT 857.125 289.765 857.295 337.875 ;
        RECT 857.125 193.205 857.295 241.315 ;
        RECT 856.665 96.645 856.835 144.755 ;
      LAYER mcon ;
        RECT 857.585 979.965 857.755 980.135 ;
        RECT 857.125 627.725 857.295 627.895 ;
        RECT 857.125 531.165 857.295 531.335 ;
        RECT 857.125 434.605 857.295 434.775 ;
        RECT 857.125 337.705 857.295 337.875 ;
        RECT 857.125 241.145 857.295 241.315 ;
        RECT 856.665 144.585 856.835 144.755 ;
      LAYER met1 ;
        RECT 857.050 1062.740 857.370 1062.800 ;
        RECT 858.890 1062.740 859.210 1062.800 ;
        RECT 857.050 1062.600 859.210 1062.740 ;
        RECT 857.050 1062.540 857.370 1062.600 ;
        RECT 858.890 1062.540 859.210 1062.600 ;
        RECT 857.050 1028.060 857.370 1028.120 ;
        RECT 857.970 1028.060 858.290 1028.120 ;
        RECT 857.050 1027.920 858.290 1028.060 ;
        RECT 857.050 1027.860 857.370 1027.920 ;
        RECT 857.970 1027.860 858.290 1027.920 ;
        RECT 857.510 980.120 857.830 980.180 ;
        RECT 857.315 979.980 857.830 980.120 ;
        RECT 857.510 979.920 857.830 979.980 ;
        RECT 857.510 966.180 857.830 966.240 ;
        RECT 857.315 966.040 857.830 966.180 ;
        RECT 857.510 965.980 857.830 966.040 ;
        RECT 857.050 821.000 857.370 821.060 ;
        RECT 857.970 821.000 858.290 821.060 ;
        RECT 857.050 820.860 858.290 821.000 ;
        RECT 857.050 820.800 857.370 820.860 ;
        RECT 857.970 820.800 858.290 820.860 ;
        RECT 857.050 724.440 857.370 724.500 ;
        RECT 857.970 724.440 858.290 724.500 ;
        RECT 857.050 724.300 858.290 724.440 ;
        RECT 857.050 724.240 857.370 724.300 ;
        RECT 857.970 724.240 858.290 724.300 ;
        RECT 857.050 627.880 857.370 627.940 ;
        RECT 856.855 627.740 857.370 627.880 ;
        RECT 857.050 627.680 857.370 627.740 ;
        RECT 857.050 579.940 857.370 580.000 ;
        RECT 856.855 579.800 857.370 579.940 ;
        RECT 857.050 579.740 857.370 579.800 ;
        RECT 857.050 531.320 857.370 531.380 ;
        RECT 856.855 531.180 857.370 531.320 ;
        RECT 857.050 531.120 857.370 531.180 ;
        RECT 857.050 483.380 857.370 483.440 ;
        RECT 856.855 483.240 857.370 483.380 ;
        RECT 857.050 483.180 857.370 483.240 ;
        RECT 857.050 434.760 857.370 434.820 ;
        RECT 856.855 434.620 857.370 434.760 ;
        RECT 857.050 434.560 857.370 434.620 ;
        RECT 857.050 386.480 857.370 386.540 ;
        RECT 856.855 386.340 857.370 386.480 ;
        RECT 857.050 386.280 857.370 386.340 ;
        RECT 857.050 337.860 857.370 337.920 ;
        RECT 856.855 337.720 857.370 337.860 ;
        RECT 857.050 337.660 857.370 337.720 ;
        RECT 857.050 289.920 857.370 289.980 ;
        RECT 856.855 289.780 857.370 289.920 ;
        RECT 857.050 289.720 857.370 289.780 ;
        RECT 857.050 241.300 857.370 241.360 ;
        RECT 856.855 241.160 857.370 241.300 ;
        RECT 857.050 241.100 857.370 241.160 ;
        RECT 857.050 193.360 857.370 193.420 ;
        RECT 856.855 193.220 857.370 193.360 ;
        RECT 857.050 193.160 857.370 193.220 ;
        RECT 856.605 144.740 856.895 144.785 ;
        RECT 857.050 144.740 857.370 144.800 ;
        RECT 856.605 144.600 857.370 144.740 ;
        RECT 856.605 144.555 856.895 144.600 ;
        RECT 857.050 144.540 857.370 144.600 ;
        RECT 856.590 96.800 856.910 96.860 ;
        RECT 856.395 96.660 856.910 96.800 ;
        RECT 856.590 96.600 856.910 96.660 ;
        RECT 855.670 62.120 855.990 62.180 ;
        RECT 856.590 62.120 856.910 62.180 ;
        RECT 855.670 61.980 856.910 62.120 ;
        RECT 855.670 61.920 855.990 61.980 ;
        RECT 856.590 61.920 856.910 61.980 ;
      LAYER via ;
        RECT 857.080 1062.540 857.340 1062.800 ;
        RECT 858.920 1062.540 859.180 1062.800 ;
        RECT 857.080 1027.860 857.340 1028.120 ;
        RECT 858.000 1027.860 858.260 1028.120 ;
        RECT 857.540 979.920 857.800 980.180 ;
        RECT 857.540 965.980 857.800 966.240 ;
        RECT 857.080 820.800 857.340 821.060 ;
        RECT 858.000 820.800 858.260 821.060 ;
        RECT 857.080 724.240 857.340 724.500 ;
        RECT 858.000 724.240 858.260 724.500 ;
        RECT 857.080 627.680 857.340 627.940 ;
        RECT 857.080 579.740 857.340 580.000 ;
        RECT 857.080 531.120 857.340 531.380 ;
        RECT 857.080 483.180 857.340 483.440 ;
        RECT 857.080 434.560 857.340 434.820 ;
        RECT 857.080 386.280 857.340 386.540 ;
        RECT 857.080 337.660 857.340 337.920 ;
        RECT 857.080 289.720 857.340 289.980 ;
        RECT 857.080 241.100 857.340 241.360 ;
        RECT 857.080 193.160 857.340 193.420 ;
        RECT 857.080 144.540 857.340 144.800 ;
        RECT 856.620 96.600 856.880 96.860 ;
        RECT 855.700 61.920 855.960 62.180 ;
        RECT 856.620 61.920 856.880 62.180 ;
      LAYER met2 ;
        RECT 858.830 1100.580 859.110 1104.000 ;
        RECT 858.830 1100.000 859.120 1100.580 ;
        RECT 858.980 1062.830 859.120 1100.000 ;
        RECT 857.080 1062.510 857.340 1062.830 ;
        RECT 858.920 1062.510 859.180 1062.830 ;
        RECT 857.140 1028.150 857.280 1062.510 ;
        RECT 857.080 1027.830 857.340 1028.150 ;
        RECT 858.000 1027.830 858.260 1028.150 ;
        RECT 858.060 1014.290 858.200 1027.830 ;
        RECT 857.600 1014.150 858.200 1014.290 ;
        RECT 857.600 980.210 857.740 1014.150 ;
        RECT 857.540 979.890 857.800 980.210 ;
        RECT 857.540 965.950 857.800 966.270 ;
        RECT 857.600 882.370 857.740 965.950 ;
        RECT 857.140 882.230 857.740 882.370 ;
        RECT 857.140 821.090 857.280 882.230 ;
        RECT 857.080 820.770 857.340 821.090 ;
        RECT 858.000 820.770 858.260 821.090 ;
        RECT 858.060 773.005 858.200 820.770 ;
        RECT 857.070 772.635 857.350 773.005 ;
        RECT 857.990 772.635 858.270 773.005 ;
        RECT 857.140 724.530 857.280 772.635 ;
        RECT 857.080 724.210 857.340 724.530 ;
        RECT 858.000 724.210 858.260 724.530 ;
        RECT 858.060 676.445 858.200 724.210 ;
        RECT 857.070 676.075 857.350 676.445 ;
        RECT 857.990 676.075 858.270 676.445 ;
        RECT 857.140 627.970 857.280 676.075 ;
        RECT 857.080 627.650 857.340 627.970 ;
        RECT 857.080 579.710 857.340 580.030 ;
        RECT 857.140 531.410 857.280 579.710 ;
        RECT 857.080 531.090 857.340 531.410 ;
        RECT 857.080 483.150 857.340 483.470 ;
        RECT 857.140 434.850 857.280 483.150 ;
        RECT 857.080 434.530 857.340 434.850 ;
        RECT 857.080 386.250 857.340 386.570 ;
        RECT 857.140 337.950 857.280 386.250 ;
        RECT 857.080 337.630 857.340 337.950 ;
        RECT 857.080 289.690 857.340 290.010 ;
        RECT 857.140 241.390 857.280 289.690 ;
        RECT 857.080 241.070 857.340 241.390 ;
        RECT 857.080 193.130 857.340 193.450 ;
        RECT 857.140 144.830 857.280 193.130 ;
        RECT 857.080 144.510 857.340 144.830 ;
        RECT 856.620 96.570 856.880 96.890 ;
        RECT 856.680 62.210 856.820 96.570 ;
        RECT 855.700 61.890 855.960 62.210 ;
        RECT 856.620 61.890 856.880 62.210 ;
        RECT 855.760 16.845 855.900 61.890 ;
        RECT 26.310 16.475 26.590 16.845 ;
        RECT 855.690 16.475 855.970 16.845 ;
        RECT 26.380 2.000 26.520 16.475 ;
        RECT 26.170 -4.000 26.730 2.000 ;
      LAYER via2 ;
        RECT 857.070 772.680 857.350 772.960 ;
        RECT 857.990 772.680 858.270 772.960 ;
        RECT 857.070 676.120 857.350 676.400 ;
        RECT 857.990 676.120 858.270 676.400 ;
        RECT 26.310 16.520 26.590 16.800 ;
        RECT 855.690 16.520 855.970 16.800 ;
      LAYER met3 ;
        RECT 857.045 772.970 857.375 772.985 ;
        RECT 857.965 772.970 858.295 772.985 ;
        RECT 857.045 772.670 858.295 772.970 ;
        RECT 857.045 772.655 857.375 772.670 ;
        RECT 857.965 772.655 858.295 772.670 ;
        RECT 857.045 676.410 857.375 676.425 ;
        RECT 857.965 676.410 858.295 676.425 ;
        RECT 857.045 676.110 858.295 676.410 ;
        RECT 857.045 676.095 857.375 676.110 ;
        RECT 857.965 676.095 858.295 676.110 ;
        RECT 26.285 16.810 26.615 16.825 ;
        RECT 855.665 16.810 855.995 16.825 ;
        RECT 26.285 16.510 855.995 16.810 ;
        RECT 26.285 16.495 26.615 16.510 ;
        RECT 855.665 16.495 855.995 16.510 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 32.270 17.580 32.590 17.640 ;
        RECT 51.590 17.580 51.910 17.640 ;
        RECT 32.270 17.440 51.910 17.580 ;
        RECT 32.270 17.380 32.590 17.440 ;
        RECT 51.590 17.380 51.910 17.440 ;
      LAYER via ;
        RECT 32.300 17.380 32.560 17.640 ;
        RECT 51.620 17.380 51.880 17.640 ;
      LAYER met2 ;
        RECT 861.130 1100.580 861.410 1104.000 ;
        RECT 861.130 1100.000 861.420 1100.580 ;
        RECT 861.280 1086.485 861.420 1100.000 ;
        RECT 51.610 1086.115 51.890 1086.485 ;
        RECT 861.210 1086.115 861.490 1086.485 ;
        RECT 51.680 17.670 51.820 1086.115 ;
        RECT 32.300 17.350 32.560 17.670 ;
        RECT 51.620 17.350 51.880 17.670 ;
        RECT 32.360 2.000 32.500 17.350 ;
        RECT 32.150 -4.000 32.710 2.000 ;
      LAYER via2 ;
        RECT 51.610 1086.160 51.890 1086.440 ;
        RECT 861.210 1086.160 861.490 1086.440 ;
      LAYER met3 ;
        RECT 51.585 1086.450 51.915 1086.465 ;
        RECT 861.185 1086.450 861.515 1086.465 ;
        RECT 51.585 1086.150 861.515 1086.450 ;
        RECT 51.585 1086.135 51.915 1086.150 ;
        RECT 861.185 1086.135 861.515 1086.150 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -9.980 -4.620 -6.980 3524.300 ;
        RECT 4.020 -9.220 7.020 3528.900 ;
        RECT 184.020 -9.220 187.020 3528.900 ;
        RECT 364.020 -9.220 367.020 3528.900 ;
        RECT 544.020 -9.220 547.020 3528.900 ;
        RECT 724.020 -9.220 727.020 3528.900 ;
        RECT 904.020 -9.220 907.020 3528.900 ;
        RECT 1084.020 -9.220 1087.020 3528.900 ;
        RECT 1264.020 -9.220 1267.020 3528.900 ;
        RECT 1444.020 -9.220 1447.020 3528.900 ;
        RECT 1624.020 -9.220 1627.020 3528.900 ;
        RECT 1804.020 -9.220 1807.020 3528.900 ;
        RECT 1984.020 -9.220 1987.020 3528.900 ;
        RECT 2164.020 -9.220 2167.020 3528.900 ;
        RECT 2344.020 -9.220 2347.020 3528.900 ;
        RECT 2524.020 -9.220 2527.020 3528.900 ;
        RECT 2704.020 -9.220 2707.020 3528.900 ;
        RECT 2884.020 -9.220 2887.020 3528.900 ;
        RECT 2926.600 -4.620 2929.600 3524.300 ;
      LAYER via4 ;
        RECT -9.070 3523.010 -7.890 3524.190 ;
        RECT -9.070 3521.410 -7.890 3522.590 ;
        RECT -9.070 3431.090 -7.890 3432.270 ;
        RECT -9.070 3429.490 -7.890 3430.670 ;
        RECT -9.070 3251.090 -7.890 3252.270 ;
        RECT -9.070 3249.490 -7.890 3250.670 ;
        RECT -9.070 3071.090 -7.890 3072.270 ;
        RECT -9.070 3069.490 -7.890 3070.670 ;
        RECT -9.070 2891.090 -7.890 2892.270 ;
        RECT -9.070 2889.490 -7.890 2890.670 ;
        RECT -9.070 2711.090 -7.890 2712.270 ;
        RECT -9.070 2709.490 -7.890 2710.670 ;
        RECT -9.070 2531.090 -7.890 2532.270 ;
        RECT -9.070 2529.490 -7.890 2530.670 ;
        RECT -9.070 2351.090 -7.890 2352.270 ;
        RECT -9.070 2349.490 -7.890 2350.670 ;
        RECT -9.070 2171.090 -7.890 2172.270 ;
        RECT -9.070 2169.490 -7.890 2170.670 ;
        RECT -9.070 1991.090 -7.890 1992.270 ;
        RECT -9.070 1989.490 -7.890 1990.670 ;
        RECT -9.070 1811.090 -7.890 1812.270 ;
        RECT -9.070 1809.490 -7.890 1810.670 ;
        RECT -9.070 1631.090 -7.890 1632.270 ;
        RECT -9.070 1629.490 -7.890 1630.670 ;
        RECT -9.070 1451.090 -7.890 1452.270 ;
        RECT -9.070 1449.490 -7.890 1450.670 ;
        RECT -9.070 1271.090 -7.890 1272.270 ;
        RECT -9.070 1269.490 -7.890 1270.670 ;
        RECT -9.070 1091.090 -7.890 1092.270 ;
        RECT -9.070 1089.490 -7.890 1090.670 ;
        RECT -9.070 911.090 -7.890 912.270 ;
        RECT -9.070 909.490 -7.890 910.670 ;
        RECT -9.070 731.090 -7.890 732.270 ;
        RECT -9.070 729.490 -7.890 730.670 ;
        RECT -9.070 551.090 -7.890 552.270 ;
        RECT -9.070 549.490 -7.890 550.670 ;
        RECT -9.070 371.090 -7.890 372.270 ;
        RECT -9.070 369.490 -7.890 370.670 ;
        RECT -9.070 191.090 -7.890 192.270 ;
        RECT -9.070 189.490 -7.890 190.670 ;
        RECT -9.070 11.090 -7.890 12.270 ;
        RECT -9.070 9.490 -7.890 10.670 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 4.930 3523.010 6.110 3524.190 ;
        RECT 4.930 3521.410 6.110 3522.590 ;
        RECT 4.930 3431.090 6.110 3432.270 ;
        RECT 4.930 3429.490 6.110 3430.670 ;
        RECT 4.930 3251.090 6.110 3252.270 ;
        RECT 4.930 3249.490 6.110 3250.670 ;
        RECT 4.930 3071.090 6.110 3072.270 ;
        RECT 4.930 3069.490 6.110 3070.670 ;
        RECT 4.930 2891.090 6.110 2892.270 ;
        RECT 4.930 2889.490 6.110 2890.670 ;
        RECT 4.930 2711.090 6.110 2712.270 ;
        RECT 4.930 2709.490 6.110 2710.670 ;
        RECT 4.930 2531.090 6.110 2532.270 ;
        RECT 4.930 2529.490 6.110 2530.670 ;
        RECT 4.930 2351.090 6.110 2352.270 ;
        RECT 4.930 2349.490 6.110 2350.670 ;
        RECT 4.930 2171.090 6.110 2172.270 ;
        RECT 4.930 2169.490 6.110 2170.670 ;
        RECT 4.930 1991.090 6.110 1992.270 ;
        RECT 4.930 1989.490 6.110 1990.670 ;
        RECT 4.930 1811.090 6.110 1812.270 ;
        RECT 4.930 1809.490 6.110 1810.670 ;
        RECT 4.930 1631.090 6.110 1632.270 ;
        RECT 4.930 1629.490 6.110 1630.670 ;
        RECT 4.930 1451.090 6.110 1452.270 ;
        RECT 4.930 1449.490 6.110 1450.670 ;
        RECT 4.930 1271.090 6.110 1272.270 ;
        RECT 4.930 1269.490 6.110 1270.670 ;
        RECT 4.930 1091.090 6.110 1092.270 ;
        RECT 4.930 1089.490 6.110 1090.670 ;
        RECT 4.930 911.090 6.110 912.270 ;
        RECT 4.930 909.490 6.110 910.670 ;
        RECT 4.930 731.090 6.110 732.270 ;
        RECT 4.930 729.490 6.110 730.670 ;
        RECT 4.930 551.090 6.110 552.270 ;
        RECT 4.930 549.490 6.110 550.670 ;
        RECT 4.930 371.090 6.110 372.270 ;
        RECT 4.930 369.490 6.110 370.670 ;
        RECT 4.930 191.090 6.110 192.270 ;
        RECT 4.930 189.490 6.110 190.670 ;
        RECT 4.930 11.090 6.110 12.270 ;
        RECT 4.930 9.490 6.110 10.670 ;
        RECT 4.930 -2.910 6.110 -1.730 ;
        RECT 4.930 -4.510 6.110 -3.330 ;
        RECT 184.930 3523.010 186.110 3524.190 ;
        RECT 184.930 3521.410 186.110 3522.590 ;
        RECT 184.930 3431.090 186.110 3432.270 ;
        RECT 184.930 3429.490 186.110 3430.670 ;
        RECT 184.930 3251.090 186.110 3252.270 ;
        RECT 184.930 3249.490 186.110 3250.670 ;
        RECT 184.930 3071.090 186.110 3072.270 ;
        RECT 184.930 3069.490 186.110 3070.670 ;
        RECT 184.930 2891.090 186.110 2892.270 ;
        RECT 184.930 2889.490 186.110 2890.670 ;
        RECT 184.930 2711.090 186.110 2712.270 ;
        RECT 184.930 2709.490 186.110 2710.670 ;
        RECT 184.930 2531.090 186.110 2532.270 ;
        RECT 184.930 2529.490 186.110 2530.670 ;
        RECT 184.930 2351.090 186.110 2352.270 ;
        RECT 184.930 2349.490 186.110 2350.670 ;
        RECT 184.930 2171.090 186.110 2172.270 ;
        RECT 184.930 2169.490 186.110 2170.670 ;
        RECT 184.930 1991.090 186.110 1992.270 ;
        RECT 184.930 1989.490 186.110 1990.670 ;
        RECT 184.930 1811.090 186.110 1812.270 ;
        RECT 184.930 1809.490 186.110 1810.670 ;
        RECT 184.930 1631.090 186.110 1632.270 ;
        RECT 184.930 1629.490 186.110 1630.670 ;
        RECT 184.930 1451.090 186.110 1452.270 ;
        RECT 184.930 1449.490 186.110 1450.670 ;
        RECT 184.930 1271.090 186.110 1272.270 ;
        RECT 184.930 1269.490 186.110 1270.670 ;
        RECT 184.930 1091.090 186.110 1092.270 ;
        RECT 184.930 1089.490 186.110 1090.670 ;
        RECT 184.930 911.090 186.110 912.270 ;
        RECT 184.930 909.490 186.110 910.670 ;
        RECT 184.930 731.090 186.110 732.270 ;
        RECT 184.930 729.490 186.110 730.670 ;
        RECT 184.930 551.090 186.110 552.270 ;
        RECT 184.930 549.490 186.110 550.670 ;
        RECT 184.930 371.090 186.110 372.270 ;
        RECT 184.930 369.490 186.110 370.670 ;
        RECT 184.930 191.090 186.110 192.270 ;
        RECT 184.930 189.490 186.110 190.670 ;
        RECT 184.930 11.090 186.110 12.270 ;
        RECT 184.930 9.490 186.110 10.670 ;
        RECT 184.930 -2.910 186.110 -1.730 ;
        RECT 184.930 -4.510 186.110 -3.330 ;
        RECT 364.930 3523.010 366.110 3524.190 ;
        RECT 364.930 3521.410 366.110 3522.590 ;
        RECT 364.930 3431.090 366.110 3432.270 ;
        RECT 364.930 3429.490 366.110 3430.670 ;
        RECT 364.930 3251.090 366.110 3252.270 ;
        RECT 364.930 3249.490 366.110 3250.670 ;
        RECT 364.930 3071.090 366.110 3072.270 ;
        RECT 364.930 3069.490 366.110 3070.670 ;
        RECT 364.930 2891.090 366.110 2892.270 ;
        RECT 364.930 2889.490 366.110 2890.670 ;
        RECT 364.930 2711.090 366.110 2712.270 ;
        RECT 364.930 2709.490 366.110 2710.670 ;
        RECT 364.930 2531.090 366.110 2532.270 ;
        RECT 364.930 2529.490 366.110 2530.670 ;
        RECT 364.930 2351.090 366.110 2352.270 ;
        RECT 364.930 2349.490 366.110 2350.670 ;
        RECT 364.930 2171.090 366.110 2172.270 ;
        RECT 364.930 2169.490 366.110 2170.670 ;
        RECT 364.930 1991.090 366.110 1992.270 ;
        RECT 364.930 1989.490 366.110 1990.670 ;
        RECT 364.930 1811.090 366.110 1812.270 ;
        RECT 364.930 1809.490 366.110 1810.670 ;
        RECT 364.930 1631.090 366.110 1632.270 ;
        RECT 364.930 1629.490 366.110 1630.670 ;
        RECT 364.930 1451.090 366.110 1452.270 ;
        RECT 364.930 1449.490 366.110 1450.670 ;
        RECT 364.930 1271.090 366.110 1272.270 ;
        RECT 364.930 1269.490 366.110 1270.670 ;
        RECT 364.930 1091.090 366.110 1092.270 ;
        RECT 364.930 1089.490 366.110 1090.670 ;
        RECT 364.930 911.090 366.110 912.270 ;
        RECT 364.930 909.490 366.110 910.670 ;
        RECT 364.930 731.090 366.110 732.270 ;
        RECT 364.930 729.490 366.110 730.670 ;
        RECT 364.930 551.090 366.110 552.270 ;
        RECT 364.930 549.490 366.110 550.670 ;
        RECT 364.930 371.090 366.110 372.270 ;
        RECT 364.930 369.490 366.110 370.670 ;
        RECT 364.930 191.090 366.110 192.270 ;
        RECT 364.930 189.490 366.110 190.670 ;
        RECT 364.930 11.090 366.110 12.270 ;
        RECT 364.930 9.490 366.110 10.670 ;
        RECT 364.930 -2.910 366.110 -1.730 ;
        RECT 364.930 -4.510 366.110 -3.330 ;
        RECT 544.930 3523.010 546.110 3524.190 ;
        RECT 544.930 3521.410 546.110 3522.590 ;
        RECT 544.930 3431.090 546.110 3432.270 ;
        RECT 544.930 3429.490 546.110 3430.670 ;
        RECT 544.930 3251.090 546.110 3252.270 ;
        RECT 544.930 3249.490 546.110 3250.670 ;
        RECT 544.930 3071.090 546.110 3072.270 ;
        RECT 544.930 3069.490 546.110 3070.670 ;
        RECT 544.930 2891.090 546.110 2892.270 ;
        RECT 544.930 2889.490 546.110 2890.670 ;
        RECT 544.930 2711.090 546.110 2712.270 ;
        RECT 544.930 2709.490 546.110 2710.670 ;
        RECT 544.930 2531.090 546.110 2532.270 ;
        RECT 544.930 2529.490 546.110 2530.670 ;
        RECT 544.930 2351.090 546.110 2352.270 ;
        RECT 544.930 2349.490 546.110 2350.670 ;
        RECT 544.930 2171.090 546.110 2172.270 ;
        RECT 544.930 2169.490 546.110 2170.670 ;
        RECT 544.930 1991.090 546.110 1992.270 ;
        RECT 544.930 1989.490 546.110 1990.670 ;
        RECT 544.930 1811.090 546.110 1812.270 ;
        RECT 544.930 1809.490 546.110 1810.670 ;
        RECT 544.930 1631.090 546.110 1632.270 ;
        RECT 544.930 1629.490 546.110 1630.670 ;
        RECT 544.930 1451.090 546.110 1452.270 ;
        RECT 544.930 1449.490 546.110 1450.670 ;
        RECT 544.930 1271.090 546.110 1272.270 ;
        RECT 544.930 1269.490 546.110 1270.670 ;
        RECT 544.930 1091.090 546.110 1092.270 ;
        RECT 544.930 1089.490 546.110 1090.670 ;
        RECT 544.930 911.090 546.110 912.270 ;
        RECT 544.930 909.490 546.110 910.670 ;
        RECT 544.930 731.090 546.110 732.270 ;
        RECT 544.930 729.490 546.110 730.670 ;
        RECT 544.930 551.090 546.110 552.270 ;
        RECT 544.930 549.490 546.110 550.670 ;
        RECT 544.930 371.090 546.110 372.270 ;
        RECT 544.930 369.490 546.110 370.670 ;
        RECT 544.930 191.090 546.110 192.270 ;
        RECT 544.930 189.490 546.110 190.670 ;
        RECT 544.930 11.090 546.110 12.270 ;
        RECT 544.930 9.490 546.110 10.670 ;
        RECT 544.930 -2.910 546.110 -1.730 ;
        RECT 544.930 -4.510 546.110 -3.330 ;
        RECT 724.930 3523.010 726.110 3524.190 ;
        RECT 724.930 3521.410 726.110 3522.590 ;
        RECT 724.930 3431.090 726.110 3432.270 ;
        RECT 724.930 3429.490 726.110 3430.670 ;
        RECT 724.930 3251.090 726.110 3252.270 ;
        RECT 724.930 3249.490 726.110 3250.670 ;
        RECT 724.930 3071.090 726.110 3072.270 ;
        RECT 724.930 3069.490 726.110 3070.670 ;
        RECT 724.930 2891.090 726.110 2892.270 ;
        RECT 724.930 2889.490 726.110 2890.670 ;
        RECT 724.930 2711.090 726.110 2712.270 ;
        RECT 724.930 2709.490 726.110 2710.670 ;
        RECT 724.930 2531.090 726.110 2532.270 ;
        RECT 724.930 2529.490 726.110 2530.670 ;
        RECT 724.930 2351.090 726.110 2352.270 ;
        RECT 724.930 2349.490 726.110 2350.670 ;
        RECT 724.930 2171.090 726.110 2172.270 ;
        RECT 724.930 2169.490 726.110 2170.670 ;
        RECT 724.930 1991.090 726.110 1992.270 ;
        RECT 724.930 1989.490 726.110 1990.670 ;
        RECT 724.930 1811.090 726.110 1812.270 ;
        RECT 724.930 1809.490 726.110 1810.670 ;
        RECT 724.930 1631.090 726.110 1632.270 ;
        RECT 724.930 1629.490 726.110 1630.670 ;
        RECT 724.930 1451.090 726.110 1452.270 ;
        RECT 724.930 1449.490 726.110 1450.670 ;
        RECT 724.930 1271.090 726.110 1272.270 ;
        RECT 724.930 1269.490 726.110 1270.670 ;
        RECT 724.930 1091.090 726.110 1092.270 ;
        RECT 724.930 1089.490 726.110 1090.670 ;
        RECT 724.930 911.090 726.110 912.270 ;
        RECT 724.930 909.490 726.110 910.670 ;
        RECT 724.930 731.090 726.110 732.270 ;
        RECT 724.930 729.490 726.110 730.670 ;
        RECT 724.930 551.090 726.110 552.270 ;
        RECT 724.930 549.490 726.110 550.670 ;
        RECT 724.930 371.090 726.110 372.270 ;
        RECT 724.930 369.490 726.110 370.670 ;
        RECT 724.930 191.090 726.110 192.270 ;
        RECT 724.930 189.490 726.110 190.670 ;
        RECT 724.930 11.090 726.110 12.270 ;
        RECT 724.930 9.490 726.110 10.670 ;
        RECT 724.930 -2.910 726.110 -1.730 ;
        RECT 724.930 -4.510 726.110 -3.330 ;
        RECT 904.930 3523.010 906.110 3524.190 ;
        RECT 904.930 3521.410 906.110 3522.590 ;
        RECT 904.930 3431.090 906.110 3432.270 ;
        RECT 904.930 3429.490 906.110 3430.670 ;
        RECT 904.930 3251.090 906.110 3252.270 ;
        RECT 904.930 3249.490 906.110 3250.670 ;
        RECT 904.930 3071.090 906.110 3072.270 ;
        RECT 904.930 3069.490 906.110 3070.670 ;
        RECT 904.930 2891.090 906.110 2892.270 ;
        RECT 904.930 2889.490 906.110 2890.670 ;
        RECT 904.930 2711.090 906.110 2712.270 ;
        RECT 904.930 2709.490 906.110 2710.670 ;
        RECT 904.930 2531.090 906.110 2532.270 ;
        RECT 904.930 2529.490 906.110 2530.670 ;
        RECT 904.930 2351.090 906.110 2352.270 ;
        RECT 904.930 2349.490 906.110 2350.670 ;
        RECT 904.930 2171.090 906.110 2172.270 ;
        RECT 904.930 2169.490 906.110 2170.670 ;
        RECT 904.930 1991.090 906.110 1992.270 ;
        RECT 904.930 1989.490 906.110 1990.670 ;
        RECT 904.930 1811.090 906.110 1812.270 ;
        RECT 904.930 1809.490 906.110 1810.670 ;
        RECT 904.930 1631.090 906.110 1632.270 ;
        RECT 904.930 1629.490 906.110 1630.670 ;
        RECT 904.930 1451.090 906.110 1452.270 ;
        RECT 904.930 1449.490 906.110 1450.670 ;
        RECT 904.930 1271.090 906.110 1272.270 ;
        RECT 904.930 1269.490 906.110 1270.670 ;
        RECT 904.930 1091.090 906.110 1092.270 ;
        RECT 904.930 1089.490 906.110 1090.670 ;
        RECT 904.930 911.090 906.110 912.270 ;
        RECT 904.930 909.490 906.110 910.670 ;
        RECT 904.930 731.090 906.110 732.270 ;
        RECT 904.930 729.490 906.110 730.670 ;
        RECT 904.930 551.090 906.110 552.270 ;
        RECT 904.930 549.490 906.110 550.670 ;
        RECT 904.930 371.090 906.110 372.270 ;
        RECT 904.930 369.490 906.110 370.670 ;
        RECT 904.930 191.090 906.110 192.270 ;
        RECT 904.930 189.490 906.110 190.670 ;
        RECT 904.930 11.090 906.110 12.270 ;
        RECT 904.930 9.490 906.110 10.670 ;
        RECT 904.930 -2.910 906.110 -1.730 ;
        RECT 904.930 -4.510 906.110 -3.330 ;
        RECT 1084.930 3523.010 1086.110 3524.190 ;
        RECT 1084.930 3521.410 1086.110 3522.590 ;
        RECT 1084.930 3431.090 1086.110 3432.270 ;
        RECT 1084.930 3429.490 1086.110 3430.670 ;
        RECT 1084.930 3251.090 1086.110 3252.270 ;
        RECT 1084.930 3249.490 1086.110 3250.670 ;
        RECT 1084.930 3071.090 1086.110 3072.270 ;
        RECT 1084.930 3069.490 1086.110 3070.670 ;
        RECT 1084.930 2891.090 1086.110 2892.270 ;
        RECT 1084.930 2889.490 1086.110 2890.670 ;
        RECT 1084.930 2711.090 1086.110 2712.270 ;
        RECT 1084.930 2709.490 1086.110 2710.670 ;
        RECT 1084.930 2531.090 1086.110 2532.270 ;
        RECT 1084.930 2529.490 1086.110 2530.670 ;
        RECT 1084.930 2351.090 1086.110 2352.270 ;
        RECT 1084.930 2349.490 1086.110 2350.670 ;
        RECT 1084.930 2171.090 1086.110 2172.270 ;
        RECT 1084.930 2169.490 1086.110 2170.670 ;
        RECT 1084.930 1991.090 1086.110 1992.270 ;
        RECT 1084.930 1989.490 1086.110 1990.670 ;
        RECT 1084.930 1811.090 1086.110 1812.270 ;
        RECT 1084.930 1809.490 1086.110 1810.670 ;
        RECT 1084.930 1631.090 1086.110 1632.270 ;
        RECT 1084.930 1629.490 1086.110 1630.670 ;
        RECT 1084.930 1451.090 1086.110 1452.270 ;
        RECT 1084.930 1449.490 1086.110 1450.670 ;
        RECT 1084.930 1271.090 1086.110 1272.270 ;
        RECT 1084.930 1269.490 1086.110 1270.670 ;
        RECT 1084.930 1091.090 1086.110 1092.270 ;
        RECT 1084.930 1089.490 1086.110 1090.670 ;
        RECT 1084.930 911.090 1086.110 912.270 ;
        RECT 1084.930 909.490 1086.110 910.670 ;
        RECT 1084.930 731.090 1086.110 732.270 ;
        RECT 1084.930 729.490 1086.110 730.670 ;
        RECT 1084.930 551.090 1086.110 552.270 ;
        RECT 1084.930 549.490 1086.110 550.670 ;
        RECT 1084.930 371.090 1086.110 372.270 ;
        RECT 1084.930 369.490 1086.110 370.670 ;
        RECT 1084.930 191.090 1086.110 192.270 ;
        RECT 1084.930 189.490 1086.110 190.670 ;
        RECT 1084.930 11.090 1086.110 12.270 ;
        RECT 1084.930 9.490 1086.110 10.670 ;
        RECT 1084.930 -2.910 1086.110 -1.730 ;
        RECT 1084.930 -4.510 1086.110 -3.330 ;
        RECT 1264.930 3523.010 1266.110 3524.190 ;
        RECT 1264.930 3521.410 1266.110 3522.590 ;
        RECT 1264.930 3431.090 1266.110 3432.270 ;
        RECT 1264.930 3429.490 1266.110 3430.670 ;
        RECT 1264.930 3251.090 1266.110 3252.270 ;
        RECT 1264.930 3249.490 1266.110 3250.670 ;
        RECT 1264.930 3071.090 1266.110 3072.270 ;
        RECT 1264.930 3069.490 1266.110 3070.670 ;
        RECT 1264.930 2891.090 1266.110 2892.270 ;
        RECT 1264.930 2889.490 1266.110 2890.670 ;
        RECT 1264.930 2711.090 1266.110 2712.270 ;
        RECT 1264.930 2709.490 1266.110 2710.670 ;
        RECT 1264.930 2531.090 1266.110 2532.270 ;
        RECT 1264.930 2529.490 1266.110 2530.670 ;
        RECT 1264.930 2351.090 1266.110 2352.270 ;
        RECT 1264.930 2349.490 1266.110 2350.670 ;
        RECT 1264.930 2171.090 1266.110 2172.270 ;
        RECT 1264.930 2169.490 1266.110 2170.670 ;
        RECT 1264.930 1991.090 1266.110 1992.270 ;
        RECT 1264.930 1989.490 1266.110 1990.670 ;
        RECT 1264.930 1811.090 1266.110 1812.270 ;
        RECT 1264.930 1809.490 1266.110 1810.670 ;
        RECT 1264.930 1631.090 1266.110 1632.270 ;
        RECT 1264.930 1629.490 1266.110 1630.670 ;
        RECT 1264.930 1451.090 1266.110 1452.270 ;
        RECT 1264.930 1449.490 1266.110 1450.670 ;
        RECT 1264.930 1271.090 1266.110 1272.270 ;
        RECT 1264.930 1269.490 1266.110 1270.670 ;
        RECT 1264.930 1091.090 1266.110 1092.270 ;
        RECT 1264.930 1089.490 1266.110 1090.670 ;
        RECT 1264.930 911.090 1266.110 912.270 ;
        RECT 1264.930 909.490 1266.110 910.670 ;
        RECT 1264.930 731.090 1266.110 732.270 ;
        RECT 1264.930 729.490 1266.110 730.670 ;
        RECT 1264.930 551.090 1266.110 552.270 ;
        RECT 1264.930 549.490 1266.110 550.670 ;
        RECT 1264.930 371.090 1266.110 372.270 ;
        RECT 1264.930 369.490 1266.110 370.670 ;
        RECT 1264.930 191.090 1266.110 192.270 ;
        RECT 1264.930 189.490 1266.110 190.670 ;
        RECT 1264.930 11.090 1266.110 12.270 ;
        RECT 1264.930 9.490 1266.110 10.670 ;
        RECT 1264.930 -2.910 1266.110 -1.730 ;
        RECT 1264.930 -4.510 1266.110 -3.330 ;
        RECT 1444.930 3523.010 1446.110 3524.190 ;
        RECT 1444.930 3521.410 1446.110 3522.590 ;
        RECT 1444.930 3431.090 1446.110 3432.270 ;
        RECT 1444.930 3429.490 1446.110 3430.670 ;
        RECT 1444.930 3251.090 1446.110 3252.270 ;
        RECT 1444.930 3249.490 1446.110 3250.670 ;
        RECT 1444.930 3071.090 1446.110 3072.270 ;
        RECT 1444.930 3069.490 1446.110 3070.670 ;
        RECT 1444.930 2891.090 1446.110 2892.270 ;
        RECT 1444.930 2889.490 1446.110 2890.670 ;
        RECT 1444.930 2711.090 1446.110 2712.270 ;
        RECT 1444.930 2709.490 1446.110 2710.670 ;
        RECT 1444.930 2531.090 1446.110 2532.270 ;
        RECT 1444.930 2529.490 1446.110 2530.670 ;
        RECT 1444.930 2351.090 1446.110 2352.270 ;
        RECT 1444.930 2349.490 1446.110 2350.670 ;
        RECT 1444.930 2171.090 1446.110 2172.270 ;
        RECT 1444.930 2169.490 1446.110 2170.670 ;
        RECT 1444.930 1991.090 1446.110 1992.270 ;
        RECT 1444.930 1989.490 1446.110 1990.670 ;
        RECT 1444.930 1811.090 1446.110 1812.270 ;
        RECT 1444.930 1809.490 1446.110 1810.670 ;
        RECT 1444.930 1631.090 1446.110 1632.270 ;
        RECT 1444.930 1629.490 1446.110 1630.670 ;
        RECT 1444.930 1451.090 1446.110 1452.270 ;
        RECT 1444.930 1449.490 1446.110 1450.670 ;
        RECT 1444.930 1271.090 1446.110 1272.270 ;
        RECT 1444.930 1269.490 1446.110 1270.670 ;
        RECT 1444.930 1091.090 1446.110 1092.270 ;
        RECT 1444.930 1089.490 1446.110 1090.670 ;
        RECT 1444.930 911.090 1446.110 912.270 ;
        RECT 1444.930 909.490 1446.110 910.670 ;
        RECT 1444.930 731.090 1446.110 732.270 ;
        RECT 1444.930 729.490 1446.110 730.670 ;
        RECT 1444.930 551.090 1446.110 552.270 ;
        RECT 1444.930 549.490 1446.110 550.670 ;
        RECT 1444.930 371.090 1446.110 372.270 ;
        RECT 1444.930 369.490 1446.110 370.670 ;
        RECT 1444.930 191.090 1446.110 192.270 ;
        RECT 1444.930 189.490 1446.110 190.670 ;
        RECT 1444.930 11.090 1446.110 12.270 ;
        RECT 1444.930 9.490 1446.110 10.670 ;
        RECT 1444.930 -2.910 1446.110 -1.730 ;
        RECT 1444.930 -4.510 1446.110 -3.330 ;
        RECT 1624.930 3523.010 1626.110 3524.190 ;
        RECT 1624.930 3521.410 1626.110 3522.590 ;
        RECT 1624.930 3431.090 1626.110 3432.270 ;
        RECT 1624.930 3429.490 1626.110 3430.670 ;
        RECT 1624.930 3251.090 1626.110 3252.270 ;
        RECT 1624.930 3249.490 1626.110 3250.670 ;
        RECT 1624.930 3071.090 1626.110 3072.270 ;
        RECT 1624.930 3069.490 1626.110 3070.670 ;
        RECT 1624.930 2891.090 1626.110 2892.270 ;
        RECT 1624.930 2889.490 1626.110 2890.670 ;
        RECT 1624.930 2711.090 1626.110 2712.270 ;
        RECT 1624.930 2709.490 1626.110 2710.670 ;
        RECT 1624.930 2531.090 1626.110 2532.270 ;
        RECT 1624.930 2529.490 1626.110 2530.670 ;
        RECT 1624.930 2351.090 1626.110 2352.270 ;
        RECT 1624.930 2349.490 1626.110 2350.670 ;
        RECT 1624.930 2171.090 1626.110 2172.270 ;
        RECT 1624.930 2169.490 1626.110 2170.670 ;
        RECT 1624.930 1991.090 1626.110 1992.270 ;
        RECT 1624.930 1989.490 1626.110 1990.670 ;
        RECT 1624.930 1811.090 1626.110 1812.270 ;
        RECT 1624.930 1809.490 1626.110 1810.670 ;
        RECT 1624.930 1631.090 1626.110 1632.270 ;
        RECT 1624.930 1629.490 1626.110 1630.670 ;
        RECT 1624.930 1451.090 1626.110 1452.270 ;
        RECT 1624.930 1449.490 1626.110 1450.670 ;
        RECT 1624.930 1271.090 1626.110 1272.270 ;
        RECT 1624.930 1269.490 1626.110 1270.670 ;
        RECT 1624.930 1091.090 1626.110 1092.270 ;
        RECT 1624.930 1089.490 1626.110 1090.670 ;
        RECT 1624.930 911.090 1626.110 912.270 ;
        RECT 1624.930 909.490 1626.110 910.670 ;
        RECT 1624.930 731.090 1626.110 732.270 ;
        RECT 1624.930 729.490 1626.110 730.670 ;
        RECT 1624.930 551.090 1626.110 552.270 ;
        RECT 1624.930 549.490 1626.110 550.670 ;
        RECT 1624.930 371.090 1626.110 372.270 ;
        RECT 1624.930 369.490 1626.110 370.670 ;
        RECT 1624.930 191.090 1626.110 192.270 ;
        RECT 1624.930 189.490 1626.110 190.670 ;
        RECT 1624.930 11.090 1626.110 12.270 ;
        RECT 1624.930 9.490 1626.110 10.670 ;
        RECT 1624.930 -2.910 1626.110 -1.730 ;
        RECT 1624.930 -4.510 1626.110 -3.330 ;
        RECT 1804.930 3523.010 1806.110 3524.190 ;
        RECT 1804.930 3521.410 1806.110 3522.590 ;
        RECT 1804.930 3431.090 1806.110 3432.270 ;
        RECT 1804.930 3429.490 1806.110 3430.670 ;
        RECT 1804.930 3251.090 1806.110 3252.270 ;
        RECT 1804.930 3249.490 1806.110 3250.670 ;
        RECT 1804.930 3071.090 1806.110 3072.270 ;
        RECT 1804.930 3069.490 1806.110 3070.670 ;
        RECT 1804.930 2891.090 1806.110 2892.270 ;
        RECT 1804.930 2889.490 1806.110 2890.670 ;
        RECT 1804.930 2711.090 1806.110 2712.270 ;
        RECT 1804.930 2709.490 1806.110 2710.670 ;
        RECT 1804.930 2531.090 1806.110 2532.270 ;
        RECT 1804.930 2529.490 1806.110 2530.670 ;
        RECT 1804.930 2351.090 1806.110 2352.270 ;
        RECT 1804.930 2349.490 1806.110 2350.670 ;
        RECT 1804.930 2171.090 1806.110 2172.270 ;
        RECT 1804.930 2169.490 1806.110 2170.670 ;
        RECT 1804.930 1991.090 1806.110 1992.270 ;
        RECT 1804.930 1989.490 1806.110 1990.670 ;
        RECT 1804.930 1811.090 1806.110 1812.270 ;
        RECT 1804.930 1809.490 1806.110 1810.670 ;
        RECT 1804.930 1631.090 1806.110 1632.270 ;
        RECT 1804.930 1629.490 1806.110 1630.670 ;
        RECT 1804.930 1451.090 1806.110 1452.270 ;
        RECT 1804.930 1449.490 1806.110 1450.670 ;
        RECT 1804.930 1271.090 1806.110 1272.270 ;
        RECT 1804.930 1269.490 1806.110 1270.670 ;
        RECT 1804.930 1091.090 1806.110 1092.270 ;
        RECT 1804.930 1089.490 1806.110 1090.670 ;
        RECT 1804.930 911.090 1806.110 912.270 ;
        RECT 1804.930 909.490 1806.110 910.670 ;
        RECT 1804.930 731.090 1806.110 732.270 ;
        RECT 1804.930 729.490 1806.110 730.670 ;
        RECT 1804.930 551.090 1806.110 552.270 ;
        RECT 1804.930 549.490 1806.110 550.670 ;
        RECT 1804.930 371.090 1806.110 372.270 ;
        RECT 1804.930 369.490 1806.110 370.670 ;
        RECT 1804.930 191.090 1806.110 192.270 ;
        RECT 1804.930 189.490 1806.110 190.670 ;
        RECT 1804.930 11.090 1806.110 12.270 ;
        RECT 1804.930 9.490 1806.110 10.670 ;
        RECT 1804.930 -2.910 1806.110 -1.730 ;
        RECT 1804.930 -4.510 1806.110 -3.330 ;
        RECT 1984.930 3523.010 1986.110 3524.190 ;
        RECT 1984.930 3521.410 1986.110 3522.590 ;
        RECT 1984.930 3431.090 1986.110 3432.270 ;
        RECT 1984.930 3429.490 1986.110 3430.670 ;
        RECT 1984.930 3251.090 1986.110 3252.270 ;
        RECT 1984.930 3249.490 1986.110 3250.670 ;
        RECT 1984.930 3071.090 1986.110 3072.270 ;
        RECT 1984.930 3069.490 1986.110 3070.670 ;
        RECT 1984.930 2891.090 1986.110 2892.270 ;
        RECT 1984.930 2889.490 1986.110 2890.670 ;
        RECT 1984.930 2711.090 1986.110 2712.270 ;
        RECT 1984.930 2709.490 1986.110 2710.670 ;
        RECT 1984.930 2531.090 1986.110 2532.270 ;
        RECT 1984.930 2529.490 1986.110 2530.670 ;
        RECT 1984.930 2351.090 1986.110 2352.270 ;
        RECT 1984.930 2349.490 1986.110 2350.670 ;
        RECT 1984.930 2171.090 1986.110 2172.270 ;
        RECT 1984.930 2169.490 1986.110 2170.670 ;
        RECT 1984.930 1991.090 1986.110 1992.270 ;
        RECT 1984.930 1989.490 1986.110 1990.670 ;
        RECT 1984.930 1811.090 1986.110 1812.270 ;
        RECT 1984.930 1809.490 1986.110 1810.670 ;
        RECT 1984.930 1631.090 1986.110 1632.270 ;
        RECT 1984.930 1629.490 1986.110 1630.670 ;
        RECT 1984.930 1451.090 1986.110 1452.270 ;
        RECT 1984.930 1449.490 1986.110 1450.670 ;
        RECT 1984.930 1271.090 1986.110 1272.270 ;
        RECT 1984.930 1269.490 1986.110 1270.670 ;
        RECT 1984.930 1091.090 1986.110 1092.270 ;
        RECT 1984.930 1089.490 1986.110 1090.670 ;
        RECT 1984.930 911.090 1986.110 912.270 ;
        RECT 1984.930 909.490 1986.110 910.670 ;
        RECT 1984.930 731.090 1986.110 732.270 ;
        RECT 1984.930 729.490 1986.110 730.670 ;
        RECT 1984.930 551.090 1986.110 552.270 ;
        RECT 1984.930 549.490 1986.110 550.670 ;
        RECT 1984.930 371.090 1986.110 372.270 ;
        RECT 1984.930 369.490 1986.110 370.670 ;
        RECT 1984.930 191.090 1986.110 192.270 ;
        RECT 1984.930 189.490 1986.110 190.670 ;
        RECT 1984.930 11.090 1986.110 12.270 ;
        RECT 1984.930 9.490 1986.110 10.670 ;
        RECT 1984.930 -2.910 1986.110 -1.730 ;
        RECT 1984.930 -4.510 1986.110 -3.330 ;
        RECT 2164.930 3523.010 2166.110 3524.190 ;
        RECT 2164.930 3521.410 2166.110 3522.590 ;
        RECT 2164.930 3431.090 2166.110 3432.270 ;
        RECT 2164.930 3429.490 2166.110 3430.670 ;
        RECT 2164.930 3251.090 2166.110 3252.270 ;
        RECT 2164.930 3249.490 2166.110 3250.670 ;
        RECT 2164.930 3071.090 2166.110 3072.270 ;
        RECT 2164.930 3069.490 2166.110 3070.670 ;
        RECT 2164.930 2891.090 2166.110 2892.270 ;
        RECT 2164.930 2889.490 2166.110 2890.670 ;
        RECT 2164.930 2711.090 2166.110 2712.270 ;
        RECT 2164.930 2709.490 2166.110 2710.670 ;
        RECT 2164.930 2531.090 2166.110 2532.270 ;
        RECT 2164.930 2529.490 2166.110 2530.670 ;
        RECT 2164.930 2351.090 2166.110 2352.270 ;
        RECT 2164.930 2349.490 2166.110 2350.670 ;
        RECT 2164.930 2171.090 2166.110 2172.270 ;
        RECT 2164.930 2169.490 2166.110 2170.670 ;
        RECT 2164.930 1991.090 2166.110 1992.270 ;
        RECT 2164.930 1989.490 2166.110 1990.670 ;
        RECT 2164.930 1811.090 2166.110 1812.270 ;
        RECT 2164.930 1809.490 2166.110 1810.670 ;
        RECT 2164.930 1631.090 2166.110 1632.270 ;
        RECT 2164.930 1629.490 2166.110 1630.670 ;
        RECT 2164.930 1451.090 2166.110 1452.270 ;
        RECT 2164.930 1449.490 2166.110 1450.670 ;
        RECT 2164.930 1271.090 2166.110 1272.270 ;
        RECT 2164.930 1269.490 2166.110 1270.670 ;
        RECT 2164.930 1091.090 2166.110 1092.270 ;
        RECT 2164.930 1089.490 2166.110 1090.670 ;
        RECT 2164.930 911.090 2166.110 912.270 ;
        RECT 2164.930 909.490 2166.110 910.670 ;
        RECT 2164.930 731.090 2166.110 732.270 ;
        RECT 2164.930 729.490 2166.110 730.670 ;
        RECT 2164.930 551.090 2166.110 552.270 ;
        RECT 2164.930 549.490 2166.110 550.670 ;
        RECT 2164.930 371.090 2166.110 372.270 ;
        RECT 2164.930 369.490 2166.110 370.670 ;
        RECT 2164.930 191.090 2166.110 192.270 ;
        RECT 2164.930 189.490 2166.110 190.670 ;
        RECT 2164.930 11.090 2166.110 12.270 ;
        RECT 2164.930 9.490 2166.110 10.670 ;
        RECT 2164.930 -2.910 2166.110 -1.730 ;
        RECT 2164.930 -4.510 2166.110 -3.330 ;
        RECT 2344.930 3523.010 2346.110 3524.190 ;
        RECT 2344.930 3521.410 2346.110 3522.590 ;
        RECT 2344.930 3431.090 2346.110 3432.270 ;
        RECT 2344.930 3429.490 2346.110 3430.670 ;
        RECT 2344.930 3251.090 2346.110 3252.270 ;
        RECT 2344.930 3249.490 2346.110 3250.670 ;
        RECT 2344.930 3071.090 2346.110 3072.270 ;
        RECT 2344.930 3069.490 2346.110 3070.670 ;
        RECT 2344.930 2891.090 2346.110 2892.270 ;
        RECT 2344.930 2889.490 2346.110 2890.670 ;
        RECT 2344.930 2711.090 2346.110 2712.270 ;
        RECT 2344.930 2709.490 2346.110 2710.670 ;
        RECT 2344.930 2531.090 2346.110 2532.270 ;
        RECT 2344.930 2529.490 2346.110 2530.670 ;
        RECT 2344.930 2351.090 2346.110 2352.270 ;
        RECT 2344.930 2349.490 2346.110 2350.670 ;
        RECT 2344.930 2171.090 2346.110 2172.270 ;
        RECT 2344.930 2169.490 2346.110 2170.670 ;
        RECT 2344.930 1991.090 2346.110 1992.270 ;
        RECT 2344.930 1989.490 2346.110 1990.670 ;
        RECT 2344.930 1811.090 2346.110 1812.270 ;
        RECT 2344.930 1809.490 2346.110 1810.670 ;
        RECT 2344.930 1631.090 2346.110 1632.270 ;
        RECT 2344.930 1629.490 2346.110 1630.670 ;
        RECT 2344.930 1451.090 2346.110 1452.270 ;
        RECT 2344.930 1449.490 2346.110 1450.670 ;
        RECT 2344.930 1271.090 2346.110 1272.270 ;
        RECT 2344.930 1269.490 2346.110 1270.670 ;
        RECT 2344.930 1091.090 2346.110 1092.270 ;
        RECT 2344.930 1089.490 2346.110 1090.670 ;
        RECT 2344.930 911.090 2346.110 912.270 ;
        RECT 2344.930 909.490 2346.110 910.670 ;
        RECT 2344.930 731.090 2346.110 732.270 ;
        RECT 2344.930 729.490 2346.110 730.670 ;
        RECT 2344.930 551.090 2346.110 552.270 ;
        RECT 2344.930 549.490 2346.110 550.670 ;
        RECT 2344.930 371.090 2346.110 372.270 ;
        RECT 2344.930 369.490 2346.110 370.670 ;
        RECT 2344.930 191.090 2346.110 192.270 ;
        RECT 2344.930 189.490 2346.110 190.670 ;
        RECT 2344.930 11.090 2346.110 12.270 ;
        RECT 2344.930 9.490 2346.110 10.670 ;
        RECT 2344.930 -2.910 2346.110 -1.730 ;
        RECT 2344.930 -4.510 2346.110 -3.330 ;
        RECT 2524.930 3523.010 2526.110 3524.190 ;
        RECT 2524.930 3521.410 2526.110 3522.590 ;
        RECT 2524.930 3431.090 2526.110 3432.270 ;
        RECT 2524.930 3429.490 2526.110 3430.670 ;
        RECT 2524.930 3251.090 2526.110 3252.270 ;
        RECT 2524.930 3249.490 2526.110 3250.670 ;
        RECT 2524.930 3071.090 2526.110 3072.270 ;
        RECT 2524.930 3069.490 2526.110 3070.670 ;
        RECT 2524.930 2891.090 2526.110 2892.270 ;
        RECT 2524.930 2889.490 2526.110 2890.670 ;
        RECT 2524.930 2711.090 2526.110 2712.270 ;
        RECT 2524.930 2709.490 2526.110 2710.670 ;
        RECT 2524.930 2531.090 2526.110 2532.270 ;
        RECT 2524.930 2529.490 2526.110 2530.670 ;
        RECT 2524.930 2351.090 2526.110 2352.270 ;
        RECT 2524.930 2349.490 2526.110 2350.670 ;
        RECT 2524.930 2171.090 2526.110 2172.270 ;
        RECT 2524.930 2169.490 2526.110 2170.670 ;
        RECT 2524.930 1991.090 2526.110 1992.270 ;
        RECT 2524.930 1989.490 2526.110 1990.670 ;
        RECT 2524.930 1811.090 2526.110 1812.270 ;
        RECT 2524.930 1809.490 2526.110 1810.670 ;
        RECT 2524.930 1631.090 2526.110 1632.270 ;
        RECT 2524.930 1629.490 2526.110 1630.670 ;
        RECT 2524.930 1451.090 2526.110 1452.270 ;
        RECT 2524.930 1449.490 2526.110 1450.670 ;
        RECT 2524.930 1271.090 2526.110 1272.270 ;
        RECT 2524.930 1269.490 2526.110 1270.670 ;
        RECT 2524.930 1091.090 2526.110 1092.270 ;
        RECT 2524.930 1089.490 2526.110 1090.670 ;
        RECT 2524.930 911.090 2526.110 912.270 ;
        RECT 2524.930 909.490 2526.110 910.670 ;
        RECT 2524.930 731.090 2526.110 732.270 ;
        RECT 2524.930 729.490 2526.110 730.670 ;
        RECT 2524.930 551.090 2526.110 552.270 ;
        RECT 2524.930 549.490 2526.110 550.670 ;
        RECT 2524.930 371.090 2526.110 372.270 ;
        RECT 2524.930 369.490 2526.110 370.670 ;
        RECT 2524.930 191.090 2526.110 192.270 ;
        RECT 2524.930 189.490 2526.110 190.670 ;
        RECT 2524.930 11.090 2526.110 12.270 ;
        RECT 2524.930 9.490 2526.110 10.670 ;
        RECT 2524.930 -2.910 2526.110 -1.730 ;
        RECT 2524.930 -4.510 2526.110 -3.330 ;
        RECT 2704.930 3523.010 2706.110 3524.190 ;
        RECT 2704.930 3521.410 2706.110 3522.590 ;
        RECT 2704.930 3431.090 2706.110 3432.270 ;
        RECT 2704.930 3429.490 2706.110 3430.670 ;
        RECT 2704.930 3251.090 2706.110 3252.270 ;
        RECT 2704.930 3249.490 2706.110 3250.670 ;
        RECT 2704.930 3071.090 2706.110 3072.270 ;
        RECT 2704.930 3069.490 2706.110 3070.670 ;
        RECT 2704.930 2891.090 2706.110 2892.270 ;
        RECT 2704.930 2889.490 2706.110 2890.670 ;
        RECT 2704.930 2711.090 2706.110 2712.270 ;
        RECT 2704.930 2709.490 2706.110 2710.670 ;
        RECT 2704.930 2531.090 2706.110 2532.270 ;
        RECT 2704.930 2529.490 2706.110 2530.670 ;
        RECT 2704.930 2351.090 2706.110 2352.270 ;
        RECT 2704.930 2349.490 2706.110 2350.670 ;
        RECT 2704.930 2171.090 2706.110 2172.270 ;
        RECT 2704.930 2169.490 2706.110 2170.670 ;
        RECT 2704.930 1991.090 2706.110 1992.270 ;
        RECT 2704.930 1989.490 2706.110 1990.670 ;
        RECT 2704.930 1811.090 2706.110 1812.270 ;
        RECT 2704.930 1809.490 2706.110 1810.670 ;
        RECT 2704.930 1631.090 2706.110 1632.270 ;
        RECT 2704.930 1629.490 2706.110 1630.670 ;
        RECT 2704.930 1451.090 2706.110 1452.270 ;
        RECT 2704.930 1449.490 2706.110 1450.670 ;
        RECT 2704.930 1271.090 2706.110 1272.270 ;
        RECT 2704.930 1269.490 2706.110 1270.670 ;
        RECT 2704.930 1091.090 2706.110 1092.270 ;
        RECT 2704.930 1089.490 2706.110 1090.670 ;
        RECT 2704.930 911.090 2706.110 912.270 ;
        RECT 2704.930 909.490 2706.110 910.670 ;
        RECT 2704.930 731.090 2706.110 732.270 ;
        RECT 2704.930 729.490 2706.110 730.670 ;
        RECT 2704.930 551.090 2706.110 552.270 ;
        RECT 2704.930 549.490 2706.110 550.670 ;
        RECT 2704.930 371.090 2706.110 372.270 ;
        RECT 2704.930 369.490 2706.110 370.670 ;
        RECT 2704.930 191.090 2706.110 192.270 ;
        RECT 2704.930 189.490 2706.110 190.670 ;
        RECT 2704.930 11.090 2706.110 12.270 ;
        RECT 2704.930 9.490 2706.110 10.670 ;
        RECT 2704.930 -2.910 2706.110 -1.730 ;
        RECT 2704.930 -4.510 2706.110 -3.330 ;
        RECT 2884.930 3523.010 2886.110 3524.190 ;
        RECT 2884.930 3521.410 2886.110 3522.590 ;
        RECT 2884.930 3431.090 2886.110 3432.270 ;
        RECT 2884.930 3429.490 2886.110 3430.670 ;
        RECT 2884.930 3251.090 2886.110 3252.270 ;
        RECT 2884.930 3249.490 2886.110 3250.670 ;
        RECT 2884.930 3071.090 2886.110 3072.270 ;
        RECT 2884.930 3069.490 2886.110 3070.670 ;
        RECT 2884.930 2891.090 2886.110 2892.270 ;
        RECT 2884.930 2889.490 2886.110 2890.670 ;
        RECT 2884.930 2711.090 2886.110 2712.270 ;
        RECT 2884.930 2709.490 2886.110 2710.670 ;
        RECT 2884.930 2531.090 2886.110 2532.270 ;
        RECT 2884.930 2529.490 2886.110 2530.670 ;
        RECT 2884.930 2351.090 2886.110 2352.270 ;
        RECT 2884.930 2349.490 2886.110 2350.670 ;
        RECT 2884.930 2171.090 2886.110 2172.270 ;
        RECT 2884.930 2169.490 2886.110 2170.670 ;
        RECT 2884.930 1991.090 2886.110 1992.270 ;
        RECT 2884.930 1989.490 2886.110 1990.670 ;
        RECT 2884.930 1811.090 2886.110 1812.270 ;
        RECT 2884.930 1809.490 2886.110 1810.670 ;
        RECT 2884.930 1631.090 2886.110 1632.270 ;
        RECT 2884.930 1629.490 2886.110 1630.670 ;
        RECT 2884.930 1451.090 2886.110 1452.270 ;
        RECT 2884.930 1449.490 2886.110 1450.670 ;
        RECT 2884.930 1271.090 2886.110 1272.270 ;
        RECT 2884.930 1269.490 2886.110 1270.670 ;
        RECT 2884.930 1091.090 2886.110 1092.270 ;
        RECT 2884.930 1089.490 2886.110 1090.670 ;
        RECT 2884.930 911.090 2886.110 912.270 ;
        RECT 2884.930 909.490 2886.110 910.670 ;
        RECT 2884.930 731.090 2886.110 732.270 ;
        RECT 2884.930 729.490 2886.110 730.670 ;
        RECT 2884.930 551.090 2886.110 552.270 ;
        RECT 2884.930 549.490 2886.110 550.670 ;
        RECT 2884.930 371.090 2886.110 372.270 ;
        RECT 2884.930 369.490 2886.110 370.670 ;
        RECT 2884.930 191.090 2886.110 192.270 ;
        RECT 2884.930 189.490 2886.110 190.670 ;
        RECT 2884.930 11.090 2886.110 12.270 ;
        RECT 2884.930 9.490 2886.110 10.670 ;
        RECT 2884.930 -2.910 2886.110 -1.730 ;
        RECT 2884.930 -4.510 2886.110 -3.330 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT 2927.510 3431.090 2928.690 3432.270 ;
        RECT 2927.510 3429.490 2928.690 3430.670 ;
        RECT 2927.510 3251.090 2928.690 3252.270 ;
        RECT 2927.510 3249.490 2928.690 3250.670 ;
        RECT 2927.510 3071.090 2928.690 3072.270 ;
        RECT 2927.510 3069.490 2928.690 3070.670 ;
        RECT 2927.510 2891.090 2928.690 2892.270 ;
        RECT 2927.510 2889.490 2928.690 2890.670 ;
        RECT 2927.510 2711.090 2928.690 2712.270 ;
        RECT 2927.510 2709.490 2928.690 2710.670 ;
        RECT 2927.510 2531.090 2928.690 2532.270 ;
        RECT 2927.510 2529.490 2928.690 2530.670 ;
        RECT 2927.510 2351.090 2928.690 2352.270 ;
        RECT 2927.510 2349.490 2928.690 2350.670 ;
        RECT 2927.510 2171.090 2928.690 2172.270 ;
        RECT 2927.510 2169.490 2928.690 2170.670 ;
        RECT 2927.510 1991.090 2928.690 1992.270 ;
        RECT 2927.510 1989.490 2928.690 1990.670 ;
        RECT 2927.510 1811.090 2928.690 1812.270 ;
        RECT 2927.510 1809.490 2928.690 1810.670 ;
        RECT 2927.510 1631.090 2928.690 1632.270 ;
        RECT 2927.510 1629.490 2928.690 1630.670 ;
        RECT 2927.510 1451.090 2928.690 1452.270 ;
        RECT 2927.510 1449.490 2928.690 1450.670 ;
        RECT 2927.510 1271.090 2928.690 1272.270 ;
        RECT 2927.510 1269.490 2928.690 1270.670 ;
        RECT 2927.510 1091.090 2928.690 1092.270 ;
        RECT 2927.510 1089.490 2928.690 1090.670 ;
        RECT 2927.510 911.090 2928.690 912.270 ;
        RECT 2927.510 909.490 2928.690 910.670 ;
        RECT 2927.510 731.090 2928.690 732.270 ;
        RECT 2927.510 729.490 2928.690 730.670 ;
        RECT 2927.510 551.090 2928.690 552.270 ;
        RECT 2927.510 549.490 2928.690 550.670 ;
        RECT 2927.510 371.090 2928.690 372.270 ;
        RECT 2927.510 369.490 2928.690 370.670 ;
        RECT 2927.510 191.090 2928.690 192.270 ;
        RECT 2927.510 189.490 2928.690 190.670 ;
        RECT 2927.510 11.090 2928.690 12.270 ;
        RECT 2927.510 9.490 2928.690 10.670 ;
        RECT 2927.510 -2.910 2928.690 -1.730 ;
        RECT 2927.510 -4.510 2928.690 -3.330 ;
      LAYER met5 ;
        RECT -9.980 3524.300 -6.980 3524.310 ;
        RECT 4.020 3524.300 7.020 3524.310 ;
        RECT 184.020 3524.300 187.020 3524.310 ;
        RECT 364.020 3524.300 367.020 3524.310 ;
        RECT 544.020 3524.300 547.020 3524.310 ;
        RECT 724.020 3524.300 727.020 3524.310 ;
        RECT 904.020 3524.300 907.020 3524.310 ;
        RECT 1084.020 3524.300 1087.020 3524.310 ;
        RECT 1264.020 3524.300 1267.020 3524.310 ;
        RECT 1444.020 3524.300 1447.020 3524.310 ;
        RECT 1624.020 3524.300 1627.020 3524.310 ;
        RECT 1804.020 3524.300 1807.020 3524.310 ;
        RECT 1984.020 3524.300 1987.020 3524.310 ;
        RECT 2164.020 3524.300 2167.020 3524.310 ;
        RECT 2344.020 3524.300 2347.020 3524.310 ;
        RECT 2524.020 3524.300 2527.020 3524.310 ;
        RECT 2704.020 3524.300 2707.020 3524.310 ;
        RECT 2884.020 3524.300 2887.020 3524.310 ;
        RECT 2926.600 3524.300 2929.600 3524.310 ;
        RECT -9.980 3521.300 2929.600 3524.300 ;
        RECT -9.980 3521.290 -6.980 3521.300 ;
        RECT 4.020 3521.290 7.020 3521.300 ;
        RECT 184.020 3521.290 187.020 3521.300 ;
        RECT 364.020 3521.290 367.020 3521.300 ;
        RECT 544.020 3521.290 547.020 3521.300 ;
        RECT 724.020 3521.290 727.020 3521.300 ;
        RECT 904.020 3521.290 907.020 3521.300 ;
        RECT 1084.020 3521.290 1087.020 3521.300 ;
        RECT 1264.020 3521.290 1267.020 3521.300 ;
        RECT 1444.020 3521.290 1447.020 3521.300 ;
        RECT 1624.020 3521.290 1627.020 3521.300 ;
        RECT 1804.020 3521.290 1807.020 3521.300 ;
        RECT 1984.020 3521.290 1987.020 3521.300 ;
        RECT 2164.020 3521.290 2167.020 3521.300 ;
        RECT 2344.020 3521.290 2347.020 3521.300 ;
        RECT 2524.020 3521.290 2527.020 3521.300 ;
        RECT 2704.020 3521.290 2707.020 3521.300 ;
        RECT 2884.020 3521.290 2887.020 3521.300 ;
        RECT 2926.600 3521.290 2929.600 3521.300 ;
        RECT -9.980 3432.380 -6.980 3432.390 ;
        RECT 4.020 3432.380 7.020 3432.390 ;
        RECT 184.020 3432.380 187.020 3432.390 ;
        RECT 364.020 3432.380 367.020 3432.390 ;
        RECT 544.020 3432.380 547.020 3432.390 ;
        RECT 724.020 3432.380 727.020 3432.390 ;
        RECT 904.020 3432.380 907.020 3432.390 ;
        RECT 1084.020 3432.380 1087.020 3432.390 ;
        RECT 1264.020 3432.380 1267.020 3432.390 ;
        RECT 1444.020 3432.380 1447.020 3432.390 ;
        RECT 1624.020 3432.380 1627.020 3432.390 ;
        RECT 1804.020 3432.380 1807.020 3432.390 ;
        RECT 1984.020 3432.380 1987.020 3432.390 ;
        RECT 2164.020 3432.380 2167.020 3432.390 ;
        RECT 2344.020 3432.380 2347.020 3432.390 ;
        RECT 2524.020 3432.380 2527.020 3432.390 ;
        RECT 2704.020 3432.380 2707.020 3432.390 ;
        RECT 2884.020 3432.380 2887.020 3432.390 ;
        RECT 2926.600 3432.380 2929.600 3432.390 ;
        RECT -14.580 3429.380 2934.200 3432.380 ;
        RECT -9.980 3429.370 -6.980 3429.380 ;
        RECT 4.020 3429.370 7.020 3429.380 ;
        RECT 184.020 3429.370 187.020 3429.380 ;
        RECT 364.020 3429.370 367.020 3429.380 ;
        RECT 544.020 3429.370 547.020 3429.380 ;
        RECT 724.020 3429.370 727.020 3429.380 ;
        RECT 904.020 3429.370 907.020 3429.380 ;
        RECT 1084.020 3429.370 1087.020 3429.380 ;
        RECT 1264.020 3429.370 1267.020 3429.380 ;
        RECT 1444.020 3429.370 1447.020 3429.380 ;
        RECT 1624.020 3429.370 1627.020 3429.380 ;
        RECT 1804.020 3429.370 1807.020 3429.380 ;
        RECT 1984.020 3429.370 1987.020 3429.380 ;
        RECT 2164.020 3429.370 2167.020 3429.380 ;
        RECT 2344.020 3429.370 2347.020 3429.380 ;
        RECT 2524.020 3429.370 2527.020 3429.380 ;
        RECT 2704.020 3429.370 2707.020 3429.380 ;
        RECT 2884.020 3429.370 2887.020 3429.380 ;
        RECT 2926.600 3429.370 2929.600 3429.380 ;
        RECT -9.980 3252.380 -6.980 3252.390 ;
        RECT 4.020 3252.380 7.020 3252.390 ;
        RECT 184.020 3252.380 187.020 3252.390 ;
        RECT 364.020 3252.380 367.020 3252.390 ;
        RECT 544.020 3252.380 547.020 3252.390 ;
        RECT 724.020 3252.380 727.020 3252.390 ;
        RECT 904.020 3252.380 907.020 3252.390 ;
        RECT 1084.020 3252.380 1087.020 3252.390 ;
        RECT 1264.020 3252.380 1267.020 3252.390 ;
        RECT 1444.020 3252.380 1447.020 3252.390 ;
        RECT 1624.020 3252.380 1627.020 3252.390 ;
        RECT 1804.020 3252.380 1807.020 3252.390 ;
        RECT 1984.020 3252.380 1987.020 3252.390 ;
        RECT 2164.020 3252.380 2167.020 3252.390 ;
        RECT 2344.020 3252.380 2347.020 3252.390 ;
        RECT 2524.020 3252.380 2527.020 3252.390 ;
        RECT 2704.020 3252.380 2707.020 3252.390 ;
        RECT 2884.020 3252.380 2887.020 3252.390 ;
        RECT 2926.600 3252.380 2929.600 3252.390 ;
        RECT -14.580 3249.380 2934.200 3252.380 ;
        RECT -9.980 3249.370 -6.980 3249.380 ;
        RECT 4.020 3249.370 7.020 3249.380 ;
        RECT 184.020 3249.370 187.020 3249.380 ;
        RECT 364.020 3249.370 367.020 3249.380 ;
        RECT 544.020 3249.370 547.020 3249.380 ;
        RECT 724.020 3249.370 727.020 3249.380 ;
        RECT 904.020 3249.370 907.020 3249.380 ;
        RECT 1084.020 3249.370 1087.020 3249.380 ;
        RECT 1264.020 3249.370 1267.020 3249.380 ;
        RECT 1444.020 3249.370 1447.020 3249.380 ;
        RECT 1624.020 3249.370 1627.020 3249.380 ;
        RECT 1804.020 3249.370 1807.020 3249.380 ;
        RECT 1984.020 3249.370 1987.020 3249.380 ;
        RECT 2164.020 3249.370 2167.020 3249.380 ;
        RECT 2344.020 3249.370 2347.020 3249.380 ;
        RECT 2524.020 3249.370 2527.020 3249.380 ;
        RECT 2704.020 3249.370 2707.020 3249.380 ;
        RECT 2884.020 3249.370 2887.020 3249.380 ;
        RECT 2926.600 3249.370 2929.600 3249.380 ;
        RECT -9.980 3072.380 -6.980 3072.390 ;
        RECT 4.020 3072.380 7.020 3072.390 ;
        RECT 184.020 3072.380 187.020 3072.390 ;
        RECT 364.020 3072.380 367.020 3072.390 ;
        RECT 544.020 3072.380 547.020 3072.390 ;
        RECT 724.020 3072.380 727.020 3072.390 ;
        RECT 904.020 3072.380 907.020 3072.390 ;
        RECT 1084.020 3072.380 1087.020 3072.390 ;
        RECT 1264.020 3072.380 1267.020 3072.390 ;
        RECT 1444.020 3072.380 1447.020 3072.390 ;
        RECT 1624.020 3072.380 1627.020 3072.390 ;
        RECT 1804.020 3072.380 1807.020 3072.390 ;
        RECT 1984.020 3072.380 1987.020 3072.390 ;
        RECT 2164.020 3072.380 2167.020 3072.390 ;
        RECT 2344.020 3072.380 2347.020 3072.390 ;
        RECT 2524.020 3072.380 2527.020 3072.390 ;
        RECT 2704.020 3072.380 2707.020 3072.390 ;
        RECT 2884.020 3072.380 2887.020 3072.390 ;
        RECT 2926.600 3072.380 2929.600 3072.390 ;
        RECT -14.580 3069.380 2934.200 3072.380 ;
        RECT -9.980 3069.370 -6.980 3069.380 ;
        RECT 4.020 3069.370 7.020 3069.380 ;
        RECT 184.020 3069.370 187.020 3069.380 ;
        RECT 364.020 3069.370 367.020 3069.380 ;
        RECT 544.020 3069.370 547.020 3069.380 ;
        RECT 724.020 3069.370 727.020 3069.380 ;
        RECT 904.020 3069.370 907.020 3069.380 ;
        RECT 1084.020 3069.370 1087.020 3069.380 ;
        RECT 1264.020 3069.370 1267.020 3069.380 ;
        RECT 1444.020 3069.370 1447.020 3069.380 ;
        RECT 1624.020 3069.370 1627.020 3069.380 ;
        RECT 1804.020 3069.370 1807.020 3069.380 ;
        RECT 1984.020 3069.370 1987.020 3069.380 ;
        RECT 2164.020 3069.370 2167.020 3069.380 ;
        RECT 2344.020 3069.370 2347.020 3069.380 ;
        RECT 2524.020 3069.370 2527.020 3069.380 ;
        RECT 2704.020 3069.370 2707.020 3069.380 ;
        RECT 2884.020 3069.370 2887.020 3069.380 ;
        RECT 2926.600 3069.370 2929.600 3069.380 ;
        RECT -9.980 2892.380 -6.980 2892.390 ;
        RECT 4.020 2892.380 7.020 2892.390 ;
        RECT 184.020 2892.380 187.020 2892.390 ;
        RECT 364.020 2892.380 367.020 2892.390 ;
        RECT 544.020 2892.380 547.020 2892.390 ;
        RECT 724.020 2892.380 727.020 2892.390 ;
        RECT 904.020 2892.380 907.020 2892.390 ;
        RECT 1084.020 2892.380 1087.020 2892.390 ;
        RECT 1264.020 2892.380 1267.020 2892.390 ;
        RECT 1444.020 2892.380 1447.020 2892.390 ;
        RECT 1624.020 2892.380 1627.020 2892.390 ;
        RECT 1804.020 2892.380 1807.020 2892.390 ;
        RECT 1984.020 2892.380 1987.020 2892.390 ;
        RECT 2164.020 2892.380 2167.020 2892.390 ;
        RECT 2344.020 2892.380 2347.020 2892.390 ;
        RECT 2524.020 2892.380 2527.020 2892.390 ;
        RECT 2704.020 2892.380 2707.020 2892.390 ;
        RECT 2884.020 2892.380 2887.020 2892.390 ;
        RECT 2926.600 2892.380 2929.600 2892.390 ;
        RECT -14.580 2889.380 2934.200 2892.380 ;
        RECT -9.980 2889.370 -6.980 2889.380 ;
        RECT 4.020 2889.370 7.020 2889.380 ;
        RECT 184.020 2889.370 187.020 2889.380 ;
        RECT 364.020 2889.370 367.020 2889.380 ;
        RECT 544.020 2889.370 547.020 2889.380 ;
        RECT 724.020 2889.370 727.020 2889.380 ;
        RECT 904.020 2889.370 907.020 2889.380 ;
        RECT 1084.020 2889.370 1087.020 2889.380 ;
        RECT 1264.020 2889.370 1267.020 2889.380 ;
        RECT 1444.020 2889.370 1447.020 2889.380 ;
        RECT 1624.020 2889.370 1627.020 2889.380 ;
        RECT 1804.020 2889.370 1807.020 2889.380 ;
        RECT 1984.020 2889.370 1987.020 2889.380 ;
        RECT 2164.020 2889.370 2167.020 2889.380 ;
        RECT 2344.020 2889.370 2347.020 2889.380 ;
        RECT 2524.020 2889.370 2527.020 2889.380 ;
        RECT 2704.020 2889.370 2707.020 2889.380 ;
        RECT 2884.020 2889.370 2887.020 2889.380 ;
        RECT 2926.600 2889.370 2929.600 2889.380 ;
        RECT -9.980 2712.380 -6.980 2712.390 ;
        RECT 4.020 2712.380 7.020 2712.390 ;
        RECT 184.020 2712.380 187.020 2712.390 ;
        RECT 364.020 2712.380 367.020 2712.390 ;
        RECT 544.020 2712.380 547.020 2712.390 ;
        RECT 724.020 2712.380 727.020 2712.390 ;
        RECT 904.020 2712.380 907.020 2712.390 ;
        RECT 1084.020 2712.380 1087.020 2712.390 ;
        RECT 1264.020 2712.380 1267.020 2712.390 ;
        RECT 1444.020 2712.380 1447.020 2712.390 ;
        RECT 1624.020 2712.380 1627.020 2712.390 ;
        RECT 1804.020 2712.380 1807.020 2712.390 ;
        RECT 1984.020 2712.380 1987.020 2712.390 ;
        RECT 2164.020 2712.380 2167.020 2712.390 ;
        RECT 2344.020 2712.380 2347.020 2712.390 ;
        RECT 2524.020 2712.380 2527.020 2712.390 ;
        RECT 2704.020 2712.380 2707.020 2712.390 ;
        RECT 2884.020 2712.380 2887.020 2712.390 ;
        RECT 2926.600 2712.380 2929.600 2712.390 ;
        RECT -14.580 2709.380 2934.200 2712.380 ;
        RECT -9.980 2709.370 -6.980 2709.380 ;
        RECT 4.020 2709.370 7.020 2709.380 ;
        RECT 184.020 2709.370 187.020 2709.380 ;
        RECT 364.020 2709.370 367.020 2709.380 ;
        RECT 544.020 2709.370 547.020 2709.380 ;
        RECT 724.020 2709.370 727.020 2709.380 ;
        RECT 904.020 2709.370 907.020 2709.380 ;
        RECT 1084.020 2709.370 1087.020 2709.380 ;
        RECT 1264.020 2709.370 1267.020 2709.380 ;
        RECT 1444.020 2709.370 1447.020 2709.380 ;
        RECT 1624.020 2709.370 1627.020 2709.380 ;
        RECT 1804.020 2709.370 1807.020 2709.380 ;
        RECT 1984.020 2709.370 1987.020 2709.380 ;
        RECT 2164.020 2709.370 2167.020 2709.380 ;
        RECT 2344.020 2709.370 2347.020 2709.380 ;
        RECT 2524.020 2709.370 2527.020 2709.380 ;
        RECT 2704.020 2709.370 2707.020 2709.380 ;
        RECT 2884.020 2709.370 2887.020 2709.380 ;
        RECT 2926.600 2709.370 2929.600 2709.380 ;
        RECT -9.980 2532.380 -6.980 2532.390 ;
        RECT 4.020 2532.380 7.020 2532.390 ;
        RECT 184.020 2532.380 187.020 2532.390 ;
        RECT 364.020 2532.380 367.020 2532.390 ;
        RECT 544.020 2532.380 547.020 2532.390 ;
        RECT 724.020 2532.380 727.020 2532.390 ;
        RECT 904.020 2532.380 907.020 2532.390 ;
        RECT 1084.020 2532.380 1087.020 2532.390 ;
        RECT 1264.020 2532.380 1267.020 2532.390 ;
        RECT 1444.020 2532.380 1447.020 2532.390 ;
        RECT 1624.020 2532.380 1627.020 2532.390 ;
        RECT 1804.020 2532.380 1807.020 2532.390 ;
        RECT 1984.020 2532.380 1987.020 2532.390 ;
        RECT 2164.020 2532.380 2167.020 2532.390 ;
        RECT 2344.020 2532.380 2347.020 2532.390 ;
        RECT 2524.020 2532.380 2527.020 2532.390 ;
        RECT 2704.020 2532.380 2707.020 2532.390 ;
        RECT 2884.020 2532.380 2887.020 2532.390 ;
        RECT 2926.600 2532.380 2929.600 2532.390 ;
        RECT -14.580 2529.380 2934.200 2532.380 ;
        RECT -9.980 2529.370 -6.980 2529.380 ;
        RECT 4.020 2529.370 7.020 2529.380 ;
        RECT 184.020 2529.370 187.020 2529.380 ;
        RECT 364.020 2529.370 367.020 2529.380 ;
        RECT 544.020 2529.370 547.020 2529.380 ;
        RECT 724.020 2529.370 727.020 2529.380 ;
        RECT 904.020 2529.370 907.020 2529.380 ;
        RECT 1084.020 2529.370 1087.020 2529.380 ;
        RECT 1264.020 2529.370 1267.020 2529.380 ;
        RECT 1444.020 2529.370 1447.020 2529.380 ;
        RECT 1624.020 2529.370 1627.020 2529.380 ;
        RECT 1804.020 2529.370 1807.020 2529.380 ;
        RECT 1984.020 2529.370 1987.020 2529.380 ;
        RECT 2164.020 2529.370 2167.020 2529.380 ;
        RECT 2344.020 2529.370 2347.020 2529.380 ;
        RECT 2524.020 2529.370 2527.020 2529.380 ;
        RECT 2704.020 2529.370 2707.020 2529.380 ;
        RECT 2884.020 2529.370 2887.020 2529.380 ;
        RECT 2926.600 2529.370 2929.600 2529.380 ;
        RECT -9.980 2352.380 -6.980 2352.390 ;
        RECT 4.020 2352.380 7.020 2352.390 ;
        RECT 184.020 2352.380 187.020 2352.390 ;
        RECT 364.020 2352.380 367.020 2352.390 ;
        RECT 544.020 2352.380 547.020 2352.390 ;
        RECT 724.020 2352.380 727.020 2352.390 ;
        RECT 904.020 2352.380 907.020 2352.390 ;
        RECT 1084.020 2352.380 1087.020 2352.390 ;
        RECT 1264.020 2352.380 1267.020 2352.390 ;
        RECT 1444.020 2352.380 1447.020 2352.390 ;
        RECT 1624.020 2352.380 1627.020 2352.390 ;
        RECT 1804.020 2352.380 1807.020 2352.390 ;
        RECT 1984.020 2352.380 1987.020 2352.390 ;
        RECT 2164.020 2352.380 2167.020 2352.390 ;
        RECT 2344.020 2352.380 2347.020 2352.390 ;
        RECT 2524.020 2352.380 2527.020 2352.390 ;
        RECT 2704.020 2352.380 2707.020 2352.390 ;
        RECT 2884.020 2352.380 2887.020 2352.390 ;
        RECT 2926.600 2352.380 2929.600 2352.390 ;
        RECT -14.580 2349.380 2934.200 2352.380 ;
        RECT -9.980 2349.370 -6.980 2349.380 ;
        RECT 4.020 2349.370 7.020 2349.380 ;
        RECT 184.020 2349.370 187.020 2349.380 ;
        RECT 364.020 2349.370 367.020 2349.380 ;
        RECT 544.020 2349.370 547.020 2349.380 ;
        RECT 724.020 2349.370 727.020 2349.380 ;
        RECT 904.020 2349.370 907.020 2349.380 ;
        RECT 1084.020 2349.370 1087.020 2349.380 ;
        RECT 1264.020 2349.370 1267.020 2349.380 ;
        RECT 1444.020 2349.370 1447.020 2349.380 ;
        RECT 1624.020 2349.370 1627.020 2349.380 ;
        RECT 1804.020 2349.370 1807.020 2349.380 ;
        RECT 1984.020 2349.370 1987.020 2349.380 ;
        RECT 2164.020 2349.370 2167.020 2349.380 ;
        RECT 2344.020 2349.370 2347.020 2349.380 ;
        RECT 2524.020 2349.370 2527.020 2349.380 ;
        RECT 2704.020 2349.370 2707.020 2349.380 ;
        RECT 2884.020 2349.370 2887.020 2349.380 ;
        RECT 2926.600 2349.370 2929.600 2349.380 ;
        RECT -9.980 2172.380 -6.980 2172.390 ;
        RECT 4.020 2172.380 7.020 2172.390 ;
        RECT 184.020 2172.380 187.020 2172.390 ;
        RECT 364.020 2172.380 367.020 2172.390 ;
        RECT 544.020 2172.380 547.020 2172.390 ;
        RECT 724.020 2172.380 727.020 2172.390 ;
        RECT 904.020 2172.380 907.020 2172.390 ;
        RECT 1084.020 2172.380 1087.020 2172.390 ;
        RECT 1264.020 2172.380 1267.020 2172.390 ;
        RECT 1444.020 2172.380 1447.020 2172.390 ;
        RECT 1624.020 2172.380 1627.020 2172.390 ;
        RECT 1804.020 2172.380 1807.020 2172.390 ;
        RECT 1984.020 2172.380 1987.020 2172.390 ;
        RECT 2164.020 2172.380 2167.020 2172.390 ;
        RECT 2344.020 2172.380 2347.020 2172.390 ;
        RECT 2524.020 2172.380 2527.020 2172.390 ;
        RECT 2704.020 2172.380 2707.020 2172.390 ;
        RECT 2884.020 2172.380 2887.020 2172.390 ;
        RECT 2926.600 2172.380 2929.600 2172.390 ;
        RECT -14.580 2169.380 2934.200 2172.380 ;
        RECT -9.980 2169.370 -6.980 2169.380 ;
        RECT 4.020 2169.370 7.020 2169.380 ;
        RECT 184.020 2169.370 187.020 2169.380 ;
        RECT 364.020 2169.370 367.020 2169.380 ;
        RECT 544.020 2169.370 547.020 2169.380 ;
        RECT 724.020 2169.370 727.020 2169.380 ;
        RECT 904.020 2169.370 907.020 2169.380 ;
        RECT 1084.020 2169.370 1087.020 2169.380 ;
        RECT 1264.020 2169.370 1267.020 2169.380 ;
        RECT 1444.020 2169.370 1447.020 2169.380 ;
        RECT 1624.020 2169.370 1627.020 2169.380 ;
        RECT 1804.020 2169.370 1807.020 2169.380 ;
        RECT 1984.020 2169.370 1987.020 2169.380 ;
        RECT 2164.020 2169.370 2167.020 2169.380 ;
        RECT 2344.020 2169.370 2347.020 2169.380 ;
        RECT 2524.020 2169.370 2527.020 2169.380 ;
        RECT 2704.020 2169.370 2707.020 2169.380 ;
        RECT 2884.020 2169.370 2887.020 2169.380 ;
        RECT 2926.600 2169.370 2929.600 2169.380 ;
        RECT -9.980 1992.380 -6.980 1992.390 ;
        RECT 4.020 1992.380 7.020 1992.390 ;
        RECT 184.020 1992.380 187.020 1992.390 ;
        RECT 364.020 1992.380 367.020 1992.390 ;
        RECT 544.020 1992.380 547.020 1992.390 ;
        RECT 724.020 1992.380 727.020 1992.390 ;
        RECT 904.020 1992.380 907.020 1992.390 ;
        RECT 1084.020 1992.380 1087.020 1992.390 ;
        RECT 1264.020 1992.380 1267.020 1992.390 ;
        RECT 1444.020 1992.380 1447.020 1992.390 ;
        RECT 1624.020 1992.380 1627.020 1992.390 ;
        RECT 1804.020 1992.380 1807.020 1992.390 ;
        RECT 1984.020 1992.380 1987.020 1992.390 ;
        RECT 2164.020 1992.380 2167.020 1992.390 ;
        RECT 2344.020 1992.380 2347.020 1992.390 ;
        RECT 2524.020 1992.380 2527.020 1992.390 ;
        RECT 2704.020 1992.380 2707.020 1992.390 ;
        RECT 2884.020 1992.380 2887.020 1992.390 ;
        RECT 2926.600 1992.380 2929.600 1992.390 ;
        RECT -14.580 1989.380 2934.200 1992.380 ;
        RECT -9.980 1989.370 -6.980 1989.380 ;
        RECT 4.020 1989.370 7.020 1989.380 ;
        RECT 184.020 1989.370 187.020 1989.380 ;
        RECT 364.020 1989.370 367.020 1989.380 ;
        RECT 544.020 1989.370 547.020 1989.380 ;
        RECT 724.020 1989.370 727.020 1989.380 ;
        RECT 904.020 1989.370 907.020 1989.380 ;
        RECT 1084.020 1989.370 1087.020 1989.380 ;
        RECT 1264.020 1989.370 1267.020 1989.380 ;
        RECT 1444.020 1989.370 1447.020 1989.380 ;
        RECT 1624.020 1989.370 1627.020 1989.380 ;
        RECT 1804.020 1989.370 1807.020 1989.380 ;
        RECT 1984.020 1989.370 1987.020 1989.380 ;
        RECT 2164.020 1989.370 2167.020 1989.380 ;
        RECT 2344.020 1989.370 2347.020 1989.380 ;
        RECT 2524.020 1989.370 2527.020 1989.380 ;
        RECT 2704.020 1989.370 2707.020 1989.380 ;
        RECT 2884.020 1989.370 2887.020 1989.380 ;
        RECT 2926.600 1989.370 2929.600 1989.380 ;
        RECT -9.980 1812.380 -6.980 1812.390 ;
        RECT 4.020 1812.380 7.020 1812.390 ;
        RECT 184.020 1812.380 187.020 1812.390 ;
        RECT 364.020 1812.380 367.020 1812.390 ;
        RECT 544.020 1812.380 547.020 1812.390 ;
        RECT 724.020 1812.380 727.020 1812.390 ;
        RECT 904.020 1812.380 907.020 1812.390 ;
        RECT 1084.020 1812.380 1087.020 1812.390 ;
        RECT 1264.020 1812.380 1267.020 1812.390 ;
        RECT 1444.020 1812.380 1447.020 1812.390 ;
        RECT 1624.020 1812.380 1627.020 1812.390 ;
        RECT 1804.020 1812.380 1807.020 1812.390 ;
        RECT 1984.020 1812.380 1987.020 1812.390 ;
        RECT 2164.020 1812.380 2167.020 1812.390 ;
        RECT 2344.020 1812.380 2347.020 1812.390 ;
        RECT 2524.020 1812.380 2527.020 1812.390 ;
        RECT 2704.020 1812.380 2707.020 1812.390 ;
        RECT 2884.020 1812.380 2887.020 1812.390 ;
        RECT 2926.600 1812.380 2929.600 1812.390 ;
        RECT -14.580 1809.380 2934.200 1812.380 ;
        RECT -9.980 1809.370 -6.980 1809.380 ;
        RECT 4.020 1809.370 7.020 1809.380 ;
        RECT 184.020 1809.370 187.020 1809.380 ;
        RECT 364.020 1809.370 367.020 1809.380 ;
        RECT 544.020 1809.370 547.020 1809.380 ;
        RECT 724.020 1809.370 727.020 1809.380 ;
        RECT 904.020 1809.370 907.020 1809.380 ;
        RECT 1084.020 1809.370 1087.020 1809.380 ;
        RECT 1264.020 1809.370 1267.020 1809.380 ;
        RECT 1444.020 1809.370 1447.020 1809.380 ;
        RECT 1624.020 1809.370 1627.020 1809.380 ;
        RECT 1804.020 1809.370 1807.020 1809.380 ;
        RECT 1984.020 1809.370 1987.020 1809.380 ;
        RECT 2164.020 1809.370 2167.020 1809.380 ;
        RECT 2344.020 1809.370 2347.020 1809.380 ;
        RECT 2524.020 1809.370 2527.020 1809.380 ;
        RECT 2704.020 1809.370 2707.020 1809.380 ;
        RECT 2884.020 1809.370 2887.020 1809.380 ;
        RECT 2926.600 1809.370 2929.600 1809.380 ;
        RECT -9.980 1632.380 -6.980 1632.390 ;
        RECT 4.020 1632.380 7.020 1632.390 ;
        RECT 184.020 1632.380 187.020 1632.390 ;
        RECT 364.020 1632.380 367.020 1632.390 ;
        RECT 544.020 1632.380 547.020 1632.390 ;
        RECT 724.020 1632.380 727.020 1632.390 ;
        RECT 904.020 1632.380 907.020 1632.390 ;
        RECT 1084.020 1632.380 1087.020 1632.390 ;
        RECT 1264.020 1632.380 1267.020 1632.390 ;
        RECT 1444.020 1632.380 1447.020 1632.390 ;
        RECT 1624.020 1632.380 1627.020 1632.390 ;
        RECT 1804.020 1632.380 1807.020 1632.390 ;
        RECT 1984.020 1632.380 1987.020 1632.390 ;
        RECT 2164.020 1632.380 2167.020 1632.390 ;
        RECT 2344.020 1632.380 2347.020 1632.390 ;
        RECT 2524.020 1632.380 2527.020 1632.390 ;
        RECT 2704.020 1632.380 2707.020 1632.390 ;
        RECT 2884.020 1632.380 2887.020 1632.390 ;
        RECT 2926.600 1632.380 2929.600 1632.390 ;
        RECT -14.580 1629.380 2934.200 1632.380 ;
        RECT -9.980 1629.370 -6.980 1629.380 ;
        RECT 4.020 1629.370 7.020 1629.380 ;
        RECT 184.020 1629.370 187.020 1629.380 ;
        RECT 364.020 1629.370 367.020 1629.380 ;
        RECT 544.020 1629.370 547.020 1629.380 ;
        RECT 724.020 1629.370 727.020 1629.380 ;
        RECT 904.020 1629.370 907.020 1629.380 ;
        RECT 1084.020 1629.370 1087.020 1629.380 ;
        RECT 1264.020 1629.370 1267.020 1629.380 ;
        RECT 1444.020 1629.370 1447.020 1629.380 ;
        RECT 1624.020 1629.370 1627.020 1629.380 ;
        RECT 1804.020 1629.370 1807.020 1629.380 ;
        RECT 1984.020 1629.370 1987.020 1629.380 ;
        RECT 2164.020 1629.370 2167.020 1629.380 ;
        RECT 2344.020 1629.370 2347.020 1629.380 ;
        RECT 2524.020 1629.370 2527.020 1629.380 ;
        RECT 2704.020 1629.370 2707.020 1629.380 ;
        RECT 2884.020 1629.370 2887.020 1629.380 ;
        RECT 2926.600 1629.370 2929.600 1629.380 ;
        RECT -9.980 1452.380 -6.980 1452.390 ;
        RECT 4.020 1452.380 7.020 1452.390 ;
        RECT 184.020 1452.380 187.020 1452.390 ;
        RECT 364.020 1452.380 367.020 1452.390 ;
        RECT 544.020 1452.380 547.020 1452.390 ;
        RECT 724.020 1452.380 727.020 1452.390 ;
        RECT 904.020 1452.380 907.020 1452.390 ;
        RECT 1084.020 1452.380 1087.020 1452.390 ;
        RECT 1264.020 1452.380 1267.020 1452.390 ;
        RECT 1444.020 1452.380 1447.020 1452.390 ;
        RECT 1624.020 1452.380 1627.020 1452.390 ;
        RECT 1804.020 1452.380 1807.020 1452.390 ;
        RECT 1984.020 1452.380 1987.020 1452.390 ;
        RECT 2164.020 1452.380 2167.020 1452.390 ;
        RECT 2344.020 1452.380 2347.020 1452.390 ;
        RECT 2524.020 1452.380 2527.020 1452.390 ;
        RECT 2704.020 1452.380 2707.020 1452.390 ;
        RECT 2884.020 1452.380 2887.020 1452.390 ;
        RECT 2926.600 1452.380 2929.600 1452.390 ;
        RECT -14.580 1449.380 2934.200 1452.380 ;
        RECT -9.980 1449.370 -6.980 1449.380 ;
        RECT 4.020 1449.370 7.020 1449.380 ;
        RECT 184.020 1449.370 187.020 1449.380 ;
        RECT 364.020 1449.370 367.020 1449.380 ;
        RECT 544.020 1449.370 547.020 1449.380 ;
        RECT 724.020 1449.370 727.020 1449.380 ;
        RECT 904.020 1449.370 907.020 1449.380 ;
        RECT 1084.020 1449.370 1087.020 1449.380 ;
        RECT 1264.020 1449.370 1267.020 1449.380 ;
        RECT 1444.020 1449.370 1447.020 1449.380 ;
        RECT 1624.020 1449.370 1627.020 1449.380 ;
        RECT 1804.020 1449.370 1807.020 1449.380 ;
        RECT 1984.020 1449.370 1987.020 1449.380 ;
        RECT 2164.020 1449.370 2167.020 1449.380 ;
        RECT 2344.020 1449.370 2347.020 1449.380 ;
        RECT 2524.020 1449.370 2527.020 1449.380 ;
        RECT 2704.020 1449.370 2707.020 1449.380 ;
        RECT 2884.020 1449.370 2887.020 1449.380 ;
        RECT 2926.600 1449.370 2929.600 1449.380 ;
        RECT -9.980 1272.380 -6.980 1272.390 ;
        RECT 4.020 1272.380 7.020 1272.390 ;
        RECT 184.020 1272.380 187.020 1272.390 ;
        RECT 364.020 1272.380 367.020 1272.390 ;
        RECT 544.020 1272.380 547.020 1272.390 ;
        RECT 724.020 1272.380 727.020 1272.390 ;
        RECT 904.020 1272.380 907.020 1272.390 ;
        RECT 1084.020 1272.380 1087.020 1272.390 ;
        RECT 1264.020 1272.380 1267.020 1272.390 ;
        RECT 1444.020 1272.380 1447.020 1272.390 ;
        RECT 1624.020 1272.380 1627.020 1272.390 ;
        RECT 1804.020 1272.380 1807.020 1272.390 ;
        RECT 1984.020 1272.380 1987.020 1272.390 ;
        RECT 2164.020 1272.380 2167.020 1272.390 ;
        RECT 2344.020 1272.380 2347.020 1272.390 ;
        RECT 2524.020 1272.380 2527.020 1272.390 ;
        RECT 2704.020 1272.380 2707.020 1272.390 ;
        RECT 2884.020 1272.380 2887.020 1272.390 ;
        RECT 2926.600 1272.380 2929.600 1272.390 ;
        RECT -14.580 1269.380 2934.200 1272.380 ;
        RECT -9.980 1269.370 -6.980 1269.380 ;
        RECT 4.020 1269.370 7.020 1269.380 ;
        RECT 184.020 1269.370 187.020 1269.380 ;
        RECT 364.020 1269.370 367.020 1269.380 ;
        RECT 544.020 1269.370 547.020 1269.380 ;
        RECT 724.020 1269.370 727.020 1269.380 ;
        RECT 904.020 1269.370 907.020 1269.380 ;
        RECT 1084.020 1269.370 1087.020 1269.380 ;
        RECT 1264.020 1269.370 1267.020 1269.380 ;
        RECT 1444.020 1269.370 1447.020 1269.380 ;
        RECT 1624.020 1269.370 1627.020 1269.380 ;
        RECT 1804.020 1269.370 1807.020 1269.380 ;
        RECT 1984.020 1269.370 1987.020 1269.380 ;
        RECT 2164.020 1269.370 2167.020 1269.380 ;
        RECT 2344.020 1269.370 2347.020 1269.380 ;
        RECT 2524.020 1269.370 2527.020 1269.380 ;
        RECT 2704.020 1269.370 2707.020 1269.380 ;
        RECT 2884.020 1269.370 2887.020 1269.380 ;
        RECT 2926.600 1269.370 2929.600 1269.380 ;
        RECT -9.980 1092.380 -6.980 1092.390 ;
        RECT 4.020 1092.380 7.020 1092.390 ;
        RECT 184.020 1092.380 187.020 1092.390 ;
        RECT 364.020 1092.380 367.020 1092.390 ;
        RECT 544.020 1092.380 547.020 1092.390 ;
        RECT 724.020 1092.380 727.020 1092.390 ;
        RECT 904.020 1092.380 907.020 1092.390 ;
        RECT 1084.020 1092.380 1087.020 1092.390 ;
        RECT 1264.020 1092.380 1267.020 1092.390 ;
        RECT 1444.020 1092.380 1447.020 1092.390 ;
        RECT 1624.020 1092.380 1627.020 1092.390 ;
        RECT 1804.020 1092.380 1807.020 1092.390 ;
        RECT 1984.020 1092.380 1987.020 1092.390 ;
        RECT 2164.020 1092.380 2167.020 1092.390 ;
        RECT 2344.020 1092.380 2347.020 1092.390 ;
        RECT 2524.020 1092.380 2527.020 1092.390 ;
        RECT 2704.020 1092.380 2707.020 1092.390 ;
        RECT 2884.020 1092.380 2887.020 1092.390 ;
        RECT 2926.600 1092.380 2929.600 1092.390 ;
        RECT -14.580 1089.380 2934.200 1092.380 ;
        RECT -9.980 1089.370 -6.980 1089.380 ;
        RECT 4.020 1089.370 7.020 1089.380 ;
        RECT 184.020 1089.370 187.020 1089.380 ;
        RECT 364.020 1089.370 367.020 1089.380 ;
        RECT 544.020 1089.370 547.020 1089.380 ;
        RECT 724.020 1089.370 727.020 1089.380 ;
        RECT 904.020 1089.370 907.020 1089.380 ;
        RECT 1084.020 1089.370 1087.020 1089.380 ;
        RECT 1264.020 1089.370 1267.020 1089.380 ;
        RECT 1444.020 1089.370 1447.020 1089.380 ;
        RECT 1624.020 1089.370 1627.020 1089.380 ;
        RECT 1804.020 1089.370 1807.020 1089.380 ;
        RECT 1984.020 1089.370 1987.020 1089.380 ;
        RECT 2164.020 1089.370 2167.020 1089.380 ;
        RECT 2344.020 1089.370 2347.020 1089.380 ;
        RECT 2524.020 1089.370 2527.020 1089.380 ;
        RECT 2704.020 1089.370 2707.020 1089.380 ;
        RECT 2884.020 1089.370 2887.020 1089.380 ;
        RECT 2926.600 1089.370 2929.600 1089.380 ;
        RECT -9.980 912.380 -6.980 912.390 ;
        RECT 4.020 912.380 7.020 912.390 ;
        RECT 184.020 912.380 187.020 912.390 ;
        RECT 364.020 912.380 367.020 912.390 ;
        RECT 544.020 912.380 547.020 912.390 ;
        RECT 724.020 912.380 727.020 912.390 ;
        RECT 904.020 912.380 907.020 912.390 ;
        RECT 1084.020 912.380 1087.020 912.390 ;
        RECT 1264.020 912.380 1267.020 912.390 ;
        RECT 1444.020 912.380 1447.020 912.390 ;
        RECT 1624.020 912.380 1627.020 912.390 ;
        RECT 1804.020 912.380 1807.020 912.390 ;
        RECT 1984.020 912.380 1987.020 912.390 ;
        RECT 2164.020 912.380 2167.020 912.390 ;
        RECT 2344.020 912.380 2347.020 912.390 ;
        RECT 2524.020 912.380 2527.020 912.390 ;
        RECT 2704.020 912.380 2707.020 912.390 ;
        RECT 2884.020 912.380 2887.020 912.390 ;
        RECT 2926.600 912.380 2929.600 912.390 ;
        RECT -14.580 909.380 2934.200 912.380 ;
        RECT -9.980 909.370 -6.980 909.380 ;
        RECT 4.020 909.370 7.020 909.380 ;
        RECT 184.020 909.370 187.020 909.380 ;
        RECT 364.020 909.370 367.020 909.380 ;
        RECT 544.020 909.370 547.020 909.380 ;
        RECT 724.020 909.370 727.020 909.380 ;
        RECT 904.020 909.370 907.020 909.380 ;
        RECT 1084.020 909.370 1087.020 909.380 ;
        RECT 1264.020 909.370 1267.020 909.380 ;
        RECT 1444.020 909.370 1447.020 909.380 ;
        RECT 1624.020 909.370 1627.020 909.380 ;
        RECT 1804.020 909.370 1807.020 909.380 ;
        RECT 1984.020 909.370 1987.020 909.380 ;
        RECT 2164.020 909.370 2167.020 909.380 ;
        RECT 2344.020 909.370 2347.020 909.380 ;
        RECT 2524.020 909.370 2527.020 909.380 ;
        RECT 2704.020 909.370 2707.020 909.380 ;
        RECT 2884.020 909.370 2887.020 909.380 ;
        RECT 2926.600 909.370 2929.600 909.380 ;
        RECT -9.980 732.380 -6.980 732.390 ;
        RECT 4.020 732.380 7.020 732.390 ;
        RECT 184.020 732.380 187.020 732.390 ;
        RECT 364.020 732.380 367.020 732.390 ;
        RECT 544.020 732.380 547.020 732.390 ;
        RECT 724.020 732.380 727.020 732.390 ;
        RECT 904.020 732.380 907.020 732.390 ;
        RECT 1084.020 732.380 1087.020 732.390 ;
        RECT 1264.020 732.380 1267.020 732.390 ;
        RECT 1444.020 732.380 1447.020 732.390 ;
        RECT 1624.020 732.380 1627.020 732.390 ;
        RECT 1804.020 732.380 1807.020 732.390 ;
        RECT 1984.020 732.380 1987.020 732.390 ;
        RECT 2164.020 732.380 2167.020 732.390 ;
        RECT 2344.020 732.380 2347.020 732.390 ;
        RECT 2524.020 732.380 2527.020 732.390 ;
        RECT 2704.020 732.380 2707.020 732.390 ;
        RECT 2884.020 732.380 2887.020 732.390 ;
        RECT 2926.600 732.380 2929.600 732.390 ;
        RECT -14.580 729.380 2934.200 732.380 ;
        RECT -9.980 729.370 -6.980 729.380 ;
        RECT 4.020 729.370 7.020 729.380 ;
        RECT 184.020 729.370 187.020 729.380 ;
        RECT 364.020 729.370 367.020 729.380 ;
        RECT 544.020 729.370 547.020 729.380 ;
        RECT 724.020 729.370 727.020 729.380 ;
        RECT 904.020 729.370 907.020 729.380 ;
        RECT 1084.020 729.370 1087.020 729.380 ;
        RECT 1264.020 729.370 1267.020 729.380 ;
        RECT 1444.020 729.370 1447.020 729.380 ;
        RECT 1624.020 729.370 1627.020 729.380 ;
        RECT 1804.020 729.370 1807.020 729.380 ;
        RECT 1984.020 729.370 1987.020 729.380 ;
        RECT 2164.020 729.370 2167.020 729.380 ;
        RECT 2344.020 729.370 2347.020 729.380 ;
        RECT 2524.020 729.370 2527.020 729.380 ;
        RECT 2704.020 729.370 2707.020 729.380 ;
        RECT 2884.020 729.370 2887.020 729.380 ;
        RECT 2926.600 729.370 2929.600 729.380 ;
        RECT -9.980 552.380 -6.980 552.390 ;
        RECT 4.020 552.380 7.020 552.390 ;
        RECT 184.020 552.380 187.020 552.390 ;
        RECT 364.020 552.380 367.020 552.390 ;
        RECT 544.020 552.380 547.020 552.390 ;
        RECT 724.020 552.380 727.020 552.390 ;
        RECT 904.020 552.380 907.020 552.390 ;
        RECT 1084.020 552.380 1087.020 552.390 ;
        RECT 1264.020 552.380 1267.020 552.390 ;
        RECT 1444.020 552.380 1447.020 552.390 ;
        RECT 1624.020 552.380 1627.020 552.390 ;
        RECT 1804.020 552.380 1807.020 552.390 ;
        RECT 1984.020 552.380 1987.020 552.390 ;
        RECT 2164.020 552.380 2167.020 552.390 ;
        RECT 2344.020 552.380 2347.020 552.390 ;
        RECT 2524.020 552.380 2527.020 552.390 ;
        RECT 2704.020 552.380 2707.020 552.390 ;
        RECT 2884.020 552.380 2887.020 552.390 ;
        RECT 2926.600 552.380 2929.600 552.390 ;
        RECT -14.580 549.380 2934.200 552.380 ;
        RECT -9.980 549.370 -6.980 549.380 ;
        RECT 4.020 549.370 7.020 549.380 ;
        RECT 184.020 549.370 187.020 549.380 ;
        RECT 364.020 549.370 367.020 549.380 ;
        RECT 544.020 549.370 547.020 549.380 ;
        RECT 724.020 549.370 727.020 549.380 ;
        RECT 904.020 549.370 907.020 549.380 ;
        RECT 1084.020 549.370 1087.020 549.380 ;
        RECT 1264.020 549.370 1267.020 549.380 ;
        RECT 1444.020 549.370 1447.020 549.380 ;
        RECT 1624.020 549.370 1627.020 549.380 ;
        RECT 1804.020 549.370 1807.020 549.380 ;
        RECT 1984.020 549.370 1987.020 549.380 ;
        RECT 2164.020 549.370 2167.020 549.380 ;
        RECT 2344.020 549.370 2347.020 549.380 ;
        RECT 2524.020 549.370 2527.020 549.380 ;
        RECT 2704.020 549.370 2707.020 549.380 ;
        RECT 2884.020 549.370 2887.020 549.380 ;
        RECT 2926.600 549.370 2929.600 549.380 ;
        RECT -9.980 372.380 -6.980 372.390 ;
        RECT 4.020 372.380 7.020 372.390 ;
        RECT 184.020 372.380 187.020 372.390 ;
        RECT 364.020 372.380 367.020 372.390 ;
        RECT 544.020 372.380 547.020 372.390 ;
        RECT 724.020 372.380 727.020 372.390 ;
        RECT 904.020 372.380 907.020 372.390 ;
        RECT 1084.020 372.380 1087.020 372.390 ;
        RECT 1264.020 372.380 1267.020 372.390 ;
        RECT 1444.020 372.380 1447.020 372.390 ;
        RECT 1624.020 372.380 1627.020 372.390 ;
        RECT 1804.020 372.380 1807.020 372.390 ;
        RECT 1984.020 372.380 1987.020 372.390 ;
        RECT 2164.020 372.380 2167.020 372.390 ;
        RECT 2344.020 372.380 2347.020 372.390 ;
        RECT 2524.020 372.380 2527.020 372.390 ;
        RECT 2704.020 372.380 2707.020 372.390 ;
        RECT 2884.020 372.380 2887.020 372.390 ;
        RECT 2926.600 372.380 2929.600 372.390 ;
        RECT -14.580 369.380 2934.200 372.380 ;
        RECT -9.980 369.370 -6.980 369.380 ;
        RECT 4.020 369.370 7.020 369.380 ;
        RECT 184.020 369.370 187.020 369.380 ;
        RECT 364.020 369.370 367.020 369.380 ;
        RECT 544.020 369.370 547.020 369.380 ;
        RECT 724.020 369.370 727.020 369.380 ;
        RECT 904.020 369.370 907.020 369.380 ;
        RECT 1084.020 369.370 1087.020 369.380 ;
        RECT 1264.020 369.370 1267.020 369.380 ;
        RECT 1444.020 369.370 1447.020 369.380 ;
        RECT 1624.020 369.370 1627.020 369.380 ;
        RECT 1804.020 369.370 1807.020 369.380 ;
        RECT 1984.020 369.370 1987.020 369.380 ;
        RECT 2164.020 369.370 2167.020 369.380 ;
        RECT 2344.020 369.370 2347.020 369.380 ;
        RECT 2524.020 369.370 2527.020 369.380 ;
        RECT 2704.020 369.370 2707.020 369.380 ;
        RECT 2884.020 369.370 2887.020 369.380 ;
        RECT 2926.600 369.370 2929.600 369.380 ;
        RECT -9.980 192.380 -6.980 192.390 ;
        RECT 4.020 192.380 7.020 192.390 ;
        RECT 184.020 192.380 187.020 192.390 ;
        RECT 364.020 192.380 367.020 192.390 ;
        RECT 544.020 192.380 547.020 192.390 ;
        RECT 724.020 192.380 727.020 192.390 ;
        RECT 904.020 192.380 907.020 192.390 ;
        RECT 1084.020 192.380 1087.020 192.390 ;
        RECT 1264.020 192.380 1267.020 192.390 ;
        RECT 1444.020 192.380 1447.020 192.390 ;
        RECT 1624.020 192.380 1627.020 192.390 ;
        RECT 1804.020 192.380 1807.020 192.390 ;
        RECT 1984.020 192.380 1987.020 192.390 ;
        RECT 2164.020 192.380 2167.020 192.390 ;
        RECT 2344.020 192.380 2347.020 192.390 ;
        RECT 2524.020 192.380 2527.020 192.390 ;
        RECT 2704.020 192.380 2707.020 192.390 ;
        RECT 2884.020 192.380 2887.020 192.390 ;
        RECT 2926.600 192.380 2929.600 192.390 ;
        RECT -14.580 189.380 2934.200 192.380 ;
        RECT -9.980 189.370 -6.980 189.380 ;
        RECT 4.020 189.370 7.020 189.380 ;
        RECT 184.020 189.370 187.020 189.380 ;
        RECT 364.020 189.370 367.020 189.380 ;
        RECT 544.020 189.370 547.020 189.380 ;
        RECT 724.020 189.370 727.020 189.380 ;
        RECT 904.020 189.370 907.020 189.380 ;
        RECT 1084.020 189.370 1087.020 189.380 ;
        RECT 1264.020 189.370 1267.020 189.380 ;
        RECT 1444.020 189.370 1447.020 189.380 ;
        RECT 1624.020 189.370 1627.020 189.380 ;
        RECT 1804.020 189.370 1807.020 189.380 ;
        RECT 1984.020 189.370 1987.020 189.380 ;
        RECT 2164.020 189.370 2167.020 189.380 ;
        RECT 2344.020 189.370 2347.020 189.380 ;
        RECT 2524.020 189.370 2527.020 189.380 ;
        RECT 2704.020 189.370 2707.020 189.380 ;
        RECT 2884.020 189.370 2887.020 189.380 ;
        RECT 2926.600 189.370 2929.600 189.380 ;
        RECT -9.980 12.380 -6.980 12.390 ;
        RECT 4.020 12.380 7.020 12.390 ;
        RECT 184.020 12.380 187.020 12.390 ;
        RECT 364.020 12.380 367.020 12.390 ;
        RECT 544.020 12.380 547.020 12.390 ;
        RECT 724.020 12.380 727.020 12.390 ;
        RECT 904.020 12.380 907.020 12.390 ;
        RECT 1084.020 12.380 1087.020 12.390 ;
        RECT 1264.020 12.380 1267.020 12.390 ;
        RECT 1444.020 12.380 1447.020 12.390 ;
        RECT 1624.020 12.380 1627.020 12.390 ;
        RECT 1804.020 12.380 1807.020 12.390 ;
        RECT 1984.020 12.380 1987.020 12.390 ;
        RECT 2164.020 12.380 2167.020 12.390 ;
        RECT 2344.020 12.380 2347.020 12.390 ;
        RECT 2524.020 12.380 2527.020 12.390 ;
        RECT 2704.020 12.380 2707.020 12.390 ;
        RECT 2884.020 12.380 2887.020 12.390 ;
        RECT 2926.600 12.380 2929.600 12.390 ;
        RECT -14.580 9.380 2934.200 12.380 ;
        RECT -9.980 9.370 -6.980 9.380 ;
        RECT 4.020 9.370 7.020 9.380 ;
        RECT 184.020 9.370 187.020 9.380 ;
        RECT 364.020 9.370 367.020 9.380 ;
        RECT 544.020 9.370 547.020 9.380 ;
        RECT 724.020 9.370 727.020 9.380 ;
        RECT 904.020 9.370 907.020 9.380 ;
        RECT 1084.020 9.370 1087.020 9.380 ;
        RECT 1264.020 9.370 1267.020 9.380 ;
        RECT 1444.020 9.370 1447.020 9.380 ;
        RECT 1624.020 9.370 1627.020 9.380 ;
        RECT 1804.020 9.370 1807.020 9.380 ;
        RECT 1984.020 9.370 1987.020 9.380 ;
        RECT 2164.020 9.370 2167.020 9.380 ;
        RECT 2344.020 9.370 2347.020 9.380 ;
        RECT 2524.020 9.370 2527.020 9.380 ;
        RECT 2704.020 9.370 2707.020 9.380 ;
        RECT 2884.020 9.370 2887.020 9.380 ;
        RECT 2926.600 9.370 2929.600 9.380 ;
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 4.020 -1.620 7.020 -1.610 ;
        RECT 184.020 -1.620 187.020 -1.610 ;
        RECT 364.020 -1.620 367.020 -1.610 ;
        RECT 544.020 -1.620 547.020 -1.610 ;
        RECT 724.020 -1.620 727.020 -1.610 ;
        RECT 904.020 -1.620 907.020 -1.610 ;
        RECT 1084.020 -1.620 1087.020 -1.610 ;
        RECT 1264.020 -1.620 1267.020 -1.610 ;
        RECT 1444.020 -1.620 1447.020 -1.610 ;
        RECT 1624.020 -1.620 1627.020 -1.610 ;
        RECT 1804.020 -1.620 1807.020 -1.610 ;
        RECT 1984.020 -1.620 1987.020 -1.610 ;
        RECT 2164.020 -1.620 2167.020 -1.610 ;
        RECT 2344.020 -1.620 2347.020 -1.610 ;
        RECT 2524.020 -1.620 2527.020 -1.610 ;
        RECT 2704.020 -1.620 2707.020 -1.610 ;
        RECT 2884.020 -1.620 2887.020 -1.610 ;
        RECT 2926.600 -1.620 2929.600 -1.610 ;
        RECT -9.980 -4.620 2929.600 -1.620 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 4.020 -4.630 7.020 -4.620 ;
        RECT 184.020 -4.630 187.020 -4.620 ;
        RECT 364.020 -4.630 367.020 -4.620 ;
        RECT 544.020 -4.630 547.020 -4.620 ;
        RECT 724.020 -4.630 727.020 -4.620 ;
        RECT 904.020 -4.630 907.020 -4.620 ;
        RECT 1084.020 -4.630 1087.020 -4.620 ;
        RECT 1264.020 -4.630 1267.020 -4.620 ;
        RECT 1444.020 -4.630 1447.020 -4.620 ;
        RECT 1624.020 -4.630 1627.020 -4.620 ;
        RECT 1804.020 -4.630 1807.020 -4.620 ;
        RECT 1984.020 -4.630 1987.020 -4.620 ;
        RECT 2164.020 -4.630 2167.020 -4.620 ;
        RECT 2344.020 -4.630 2347.020 -4.620 ;
        RECT 2524.020 -4.630 2527.020 -4.620 ;
        RECT 2704.020 -4.630 2707.020 -4.620 ;
        RECT 2884.020 -4.630 2887.020 -4.620 ;
        RECT 2926.600 -4.630 2929.600 -4.620 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -14.580 -9.220 -11.580 3528.900 ;
        RECT 94.020 -9.220 97.020 3528.900 ;
        RECT 274.020 -9.220 277.020 3528.900 ;
        RECT 454.020 -9.220 457.020 3528.900 ;
        RECT 634.020 -9.220 637.020 3528.900 ;
        RECT 814.020 -9.220 817.020 3528.900 ;
        RECT 994.020 -9.220 997.020 3528.900 ;
        RECT 1174.020 -9.220 1177.020 3528.900 ;
        RECT 1354.020 -9.220 1357.020 3528.900 ;
        RECT 1534.020 -9.220 1537.020 3528.900 ;
        RECT 1714.020 -9.220 1717.020 3528.900 ;
        RECT 1894.020 -9.220 1897.020 3528.900 ;
        RECT 2074.020 -9.220 2077.020 3528.900 ;
        RECT 2254.020 -9.220 2257.020 3528.900 ;
        RECT 2434.020 -9.220 2437.020 3528.900 ;
        RECT 2614.020 -9.220 2617.020 3528.900 ;
        RECT 2794.020 -9.220 2797.020 3528.900 ;
        RECT 2931.200 -9.220 2934.200 3528.900 ;
      LAYER via4 ;
        RECT -13.670 3527.610 -12.490 3528.790 ;
        RECT -13.670 3526.010 -12.490 3527.190 ;
        RECT -13.670 3341.090 -12.490 3342.270 ;
        RECT -13.670 3339.490 -12.490 3340.670 ;
        RECT -13.670 3161.090 -12.490 3162.270 ;
        RECT -13.670 3159.490 -12.490 3160.670 ;
        RECT -13.670 2981.090 -12.490 2982.270 ;
        RECT -13.670 2979.490 -12.490 2980.670 ;
        RECT -13.670 2801.090 -12.490 2802.270 ;
        RECT -13.670 2799.490 -12.490 2800.670 ;
        RECT -13.670 2621.090 -12.490 2622.270 ;
        RECT -13.670 2619.490 -12.490 2620.670 ;
        RECT -13.670 2441.090 -12.490 2442.270 ;
        RECT -13.670 2439.490 -12.490 2440.670 ;
        RECT -13.670 2261.090 -12.490 2262.270 ;
        RECT -13.670 2259.490 -12.490 2260.670 ;
        RECT -13.670 2081.090 -12.490 2082.270 ;
        RECT -13.670 2079.490 -12.490 2080.670 ;
        RECT -13.670 1901.090 -12.490 1902.270 ;
        RECT -13.670 1899.490 -12.490 1900.670 ;
        RECT -13.670 1721.090 -12.490 1722.270 ;
        RECT -13.670 1719.490 -12.490 1720.670 ;
        RECT -13.670 1541.090 -12.490 1542.270 ;
        RECT -13.670 1539.490 -12.490 1540.670 ;
        RECT -13.670 1361.090 -12.490 1362.270 ;
        RECT -13.670 1359.490 -12.490 1360.670 ;
        RECT -13.670 1181.090 -12.490 1182.270 ;
        RECT -13.670 1179.490 -12.490 1180.670 ;
        RECT -13.670 1001.090 -12.490 1002.270 ;
        RECT -13.670 999.490 -12.490 1000.670 ;
        RECT -13.670 821.090 -12.490 822.270 ;
        RECT -13.670 819.490 -12.490 820.670 ;
        RECT -13.670 641.090 -12.490 642.270 ;
        RECT -13.670 639.490 -12.490 640.670 ;
        RECT -13.670 461.090 -12.490 462.270 ;
        RECT -13.670 459.490 -12.490 460.670 ;
        RECT -13.670 281.090 -12.490 282.270 ;
        RECT -13.670 279.490 -12.490 280.670 ;
        RECT -13.670 101.090 -12.490 102.270 ;
        RECT -13.670 99.490 -12.490 100.670 ;
        RECT -13.670 -7.510 -12.490 -6.330 ;
        RECT -13.670 -9.110 -12.490 -7.930 ;
        RECT 94.930 3527.610 96.110 3528.790 ;
        RECT 94.930 3526.010 96.110 3527.190 ;
        RECT 94.930 3341.090 96.110 3342.270 ;
        RECT 94.930 3339.490 96.110 3340.670 ;
        RECT 94.930 3161.090 96.110 3162.270 ;
        RECT 94.930 3159.490 96.110 3160.670 ;
        RECT 94.930 2981.090 96.110 2982.270 ;
        RECT 94.930 2979.490 96.110 2980.670 ;
        RECT 94.930 2801.090 96.110 2802.270 ;
        RECT 94.930 2799.490 96.110 2800.670 ;
        RECT 94.930 2621.090 96.110 2622.270 ;
        RECT 94.930 2619.490 96.110 2620.670 ;
        RECT 94.930 2441.090 96.110 2442.270 ;
        RECT 94.930 2439.490 96.110 2440.670 ;
        RECT 94.930 2261.090 96.110 2262.270 ;
        RECT 94.930 2259.490 96.110 2260.670 ;
        RECT 94.930 2081.090 96.110 2082.270 ;
        RECT 94.930 2079.490 96.110 2080.670 ;
        RECT 94.930 1901.090 96.110 1902.270 ;
        RECT 94.930 1899.490 96.110 1900.670 ;
        RECT 94.930 1721.090 96.110 1722.270 ;
        RECT 94.930 1719.490 96.110 1720.670 ;
        RECT 94.930 1541.090 96.110 1542.270 ;
        RECT 94.930 1539.490 96.110 1540.670 ;
        RECT 94.930 1361.090 96.110 1362.270 ;
        RECT 94.930 1359.490 96.110 1360.670 ;
        RECT 94.930 1181.090 96.110 1182.270 ;
        RECT 94.930 1179.490 96.110 1180.670 ;
        RECT 94.930 1001.090 96.110 1002.270 ;
        RECT 94.930 999.490 96.110 1000.670 ;
        RECT 94.930 821.090 96.110 822.270 ;
        RECT 94.930 819.490 96.110 820.670 ;
        RECT 94.930 641.090 96.110 642.270 ;
        RECT 94.930 639.490 96.110 640.670 ;
        RECT 94.930 461.090 96.110 462.270 ;
        RECT 94.930 459.490 96.110 460.670 ;
        RECT 94.930 281.090 96.110 282.270 ;
        RECT 94.930 279.490 96.110 280.670 ;
        RECT 94.930 101.090 96.110 102.270 ;
        RECT 94.930 99.490 96.110 100.670 ;
        RECT 94.930 -7.510 96.110 -6.330 ;
        RECT 94.930 -9.110 96.110 -7.930 ;
        RECT 274.930 3527.610 276.110 3528.790 ;
        RECT 274.930 3526.010 276.110 3527.190 ;
        RECT 274.930 3341.090 276.110 3342.270 ;
        RECT 274.930 3339.490 276.110 3340.670 ;
        RECT 274.930 3161.090 276.110 3162.270 ;
        RECT 274.930 3159.490 276.110 3160.670 ;
        RECT 274.930 2981.090 276.110 2982.270 ;
        RECT 274.930 2979.490 276.110 2980.670 ;
        RECT 274.930 2801.090 276.110 2802.270 ;
        RECT 274.930 2799.490 276.110 2800.670 ;
        RECT 274.930 2621.090 276.110 2622.270 ;
        RECT 274.930 2619.490 276.110 2620.670 ;
        RECT 274.930 2441.090 276.110 2442.270 ;
        RECT 274.930 2439.490 276.110 2440.670 ;
        RECT 274.930 2261.090 276.110 2262.270 ;
        RECT 274.930 2259.490 276.110 2260.670 ;
        RECT 274.930 2081.090 276.110 2082.270 ;
        RECT 274.930 2079.490 276.110 2080.670 ;
        RECT 274.930 1901.090 276.110 1902.270 ;
        RECT 274.930 1899.490 276.110 1900.670 ;
        RECT 274.930 1721.090 276.110 1722.270 ;
        RECT 274.930 1719.490 276.110 1720.670 ;
        RECT 274.930 1541.090 276.110 1542.270 ;
        RECT 274.930 1539.490 276.110 1540.670 ;
        RECT 274.930 1361.090 276.110 1362.270 ;
        RECT 274.930 1359.490 276.110 1360.670 ;
        RECT 274.930 1181.090 276.110 1182.270 ;
        RECT 274.930 1179.490 276.110 1180.670 ;
        RECT 274.930 1001.090 276.110 1002.270 ;
        RECT 274.930 999.490 276.110 1000.670 ;
        RECT 274.930 821.090 276.110 822.270 ;
        RECT 274.930 819.490 276.110 820.670 ;
        RECT 274.930 641.090 276.110 642.270 ;
        RECT 274.930 639.490 276.110 640.670 ;
        RECT 274.930 461.090 276.110 462.270 ;
        RECT 274.930 459.490 276.110 460.670 ;
        RECT 274.930 281.090 276.110 282.270 ;
        RECT 274.930 279.490 276.110 280.670 ;
        RECT 274.930 101.090 276.110 102.270 ;
        RECT 274.930 99.490 276.110 100.670 ;
        RECT 274.930 -7.510 276.110 -6.330 ;
        RECT 274.930 -9.110 276.110 -7.930 ;
        RECT 454.930 3527.610 456.110 3528.790 ;
        RECT 454.930 3526.010 456.110 3527.190 ;
        RECT 454.930 3341.090 456.110 3342.270 ;
        RECT 454.930 3339.490 456.110 3340.670 ;
        RECT 454.930 3161.090 456.110 3162.270 ;
        RECT 454.930 3159.490 456.110 3160.670 ;
        RECT 454.930 2981.090 456.110 2982.270 ;
        RECT 454.930 2979.490 456.110 2980.670 ;
        RECT 454.930 2801.090 456.110 2802.270 ;
        RECT 454.930 2799.490 456.110 2800.670 ;
        RECT 454.930 2621.090 456.110 2622.270 ;
        RECT 454.930 2619.490 456.110 2620.670 ;
        RECT 454.930 2441.090 456.110 2442.270 ;
        RECT 454.930 2439.490 456.110 2440.670 ;
        RECT 454.930 2261.090 456.110 2262.270 ;
        RECT 454.930 2259.490 456.110 2260.670 ;
        RECT 454.930 2081.090 456.110 2082.270 ;
        RECT 454.930 2079.490 456.110 2080.670 ;
        RECT 454.930 1901.090 456.110 1902.270 ;
        RECT 454.930 1899.490 456.110 1900.670 ;
        RECT 454.930 1721.090 456.110 1722.270 ;
        RECT 454.930 1719.490 456.110 1720.670 ;
        RECT 454.930 1541.090 456.110 1542.270 ;
        RECT 454.930 1539.490 456.110 1540.670 ;
        RECT 454.930 1361.090 456.110 1362.270 ;
        RECT 454.930 1359.490 456.110 1360.670 ;
        RECT 454.930 1181.090 456.110 1182.270 ;
        RECT 454.930 1179.490 456.110 1180.670 ;
        RECT 454.930 1001.090 456.110 1002.270 ;
        RECT 454.930 999.490 456.110 1000.670 ;
        RECT 454.930 821.090 456.110 822.270 ;
        RECT 454.930 819.490 456.110 820.670 ;
        RECT 454.930 641.090 456.110 642.270 ;
        RECT 454.930 639.490 456.110 640.670 ;
        RECT 454.930 461.090 456.110 462.270 ;
        RECT 454.930 459.490 456.110 460.670 ;
        RECT 454.930 281.090 456.110 282.270 ;
        RECT 454.930 279.490 456.110 280.670 ;
        RECT 454.930 101.090 456.110 102.270 ;
        RECT 454.930 99.490 456.110 100.670 ;
        RECT 454.930 -7.510 456.110 -6.330 ;
        RECT 454.930 -9.110 456.110 -7.930 ;
        RECT 634.930 3527.610 636.110 3528.790 ;
        RECT 634.930 3526.010 636.110 3527.190 ;
        RECT 634.930 3341.090 636.110 3342.270 ;
        RECT 634.930 3339.490 636.110 3340.670 ;
        RECT 634.930 3161.090 636.110 3162.270 ;
        RECT 634.930 3159.490 636.110 3160.670 ;
        RECT 634.930 2981.090 636.110 2982.270 ;
        RECT 634.930 2979.490 636.110 2980.670 ;
        RECT 634.930 2801.090 636.110 2802.270 ;
        RECT 634.930 2799.490 636.110 2800.670 ;
        RECT 634.930 2621.090 636.110 2622.270 ;
        RECT 634.930 2619.490 636.110 2620.670 ;
        RECT 634.930 2441.090 636.110 2442.270 ;
        RECT 634.930 2439.490 636.110 2440.670 ;
        RECT 634.930 2261.090 636.110 2262.270 ;
        RECT 634.930 2259.490 636.110 2260.670 ;
        RECT 634.930 2081.090 636.110 2082.270 ;
        RECT 634.930 2079.490 636.110 2080.670 ;
        RECT 634.930 1901.090 636.110 1902.270 ;
        RECT 634.930 1899.490 636.110 1900.670 ;
        RECT 634.930 1721.090 636.110 1722.270 ;
        RECT 634.930 1719.490 636.110 1720.670 ;
        RECT 634.930 1541.090 636.110 1542.270 ;
        RECT 634.930 1539.490 636.110 1540.670 ;
        RECT 634.930 1361.090 636.110 1362.270 ;
        RECT 634.930 1359.490 636.110 1360.670 ;
        RECT 634.930 1181.090 636.110 1182.270 ;
        RECT 634.930 1179.490 636.110 1180.670 ;
        RECT 634.930 1001.090 636.110 1002.270 ;
        RECT 634.930 999.490 636.110 1000.670 ;
        RECT 634.930 821.090 636.110 822.270 ;
        RECT 634.930 819.490 636.110 820.670 ;
        RECT 634.930 641.090 636.110 642.270 ;
        RECT 634.930 639.490 636.110 640.670 ;
        RECT 634.930 461.090 636.110 462.270 ;
        RECT 634.930 459.490 636.110 460.670 ;
        RECT 634.930 281.090 636.110 282.270 ;
        RECT 634.930 279.490 636.110 280.670 ;
        RECT 634.930 101.090 636.110 102.270 ;
        RECT 634.930 99.490 636.110 100.670 ;
        RECT 634.930 -7.510 636.110 -6.330 ;
        RECT 634.930 -9.110 636.110 -7.930 ;
        RECT 814.930 3527.610 816.110 3528.790 ;
        RECT 814.930 3526.010 816.110 3527.190 ;
        RECT 814.930 3341.090 816.110 3342.270 ;
        RECT 814.930 3339.490 816.110 3340.670 ;
        RECT 814.930 3161.090 816.110 3162.270 ;
        RECT 814.930 3159.490 816.110 3160.670 ;
        RECT 814.930 2981.090 816.110 2982.270 ;
        RECT 814.930 2979.490 816.110 2980.670 ;
        RECT 814.930 2801.090 816.110 2802.270 ;
        RECT 814.930 2799.490 816.110 2800.670 ;
        RECT 814.930 2621.090 816.110 2622.270 ;
        RECT 814.930 2619.490 816.110 2620.670 ;
        RECT 814.930 2441.090 816.110 2442.270 ;
        RECT 814.930 2439.490 816.110 2440.670 ;
        RECT 814.930 2261.090 816.110 2262.270 ;
        RECT 814.930 2259.490 816.110 2260.670 ;
        RECT 814.930 2081.090 816.110 2082.270 ;
        RECT 814.930 2079.490 816.110 2080.670 ;
        RECT 814.930 1901.090 816.110 1902.270 ;
        RECT 814.930 1899.490 816.110 1900.670 ;
        RECT 814.930 1721.090 816.110 1722.270 ;
        RECT 814.930 1719.490 816.110 1720.670 ;
        RECT 814.930 1541.090 816.110 1542.270 ;
        RECT 814.930 1539.490 816.110 1540.670 ;
        RECT 814.930 1361.090 816.110 1362.270 ;
        RECT 814.930 1359.490 816.110 1360.670 ;
        RECT 814.930 1181.090 816.110 1182.270 ;
        RECT 814.930 1179.490 816.110 1180.670 ;
        RECT 814.930 1001.090 816.110 1002.270 ;
        RECT 814.930 999.490 816.110 1000.670 ;
        RECT 814.930 821.090 816.110 822.270 ;
        RECT 814.930 819.490 816.110 820.670 ;
        RECT 814.930 641.090 816.110 642.270 ;
        RECT 814.930 639.490 816.110 640.670 ;
        RECT 814.930 461.090 816.110 462.270 ;
        RECT 814.930 459.490 816.110 460.670 ;
        RECT 814.930 281.090 816.110 282.270 ;
        RECT 814.930 279.490 816.110 280.670 ;
        RECT 814.930 101.090 816.110 102.270 ;
        RECT 814.930 99.490 816.110 100.670 ;
        RECT 814.930 -7.510 816.110 -6.330 ;
        RECT 814.930 -9.110 816.110 -7.930 ;
        RECT 994.930 3527.610 996.110 3528.790 ;
        RECT 994.930 3526.010 996.110 3527.190 ;
        RECT 994.930 3341.090 996.110 3342.270 ;
        RECT 994.930 3339.490 996.110 3340.670 ;
        RECT 994.930 3161.090 996.110 3162.270 ;
        RECT 994.930 3159.490 996.110 3160.670 ;
        RECT 994.930 2981.090 996.110 2982.270 ;
        RECT 994.930 2979.490 996.110 2980.670 ;
        RECT 994.930 2801.090 996.110 2802.270 ;
        RECT 994.930 2799.490 996.110 2800.670 ;
        RECT 994.930 2621.090 996.110 2622.270 ;
        RECT 994.930 2619.490 996.110 2620.670 ;
        RECT 994.930 2441.090 996.110 2442.270 ;
        RECT 994.930 2439.490 996.110 2440.670 ;
        RECT 994.930 2261.090 996.110 2262.270 ;
        RECT 994.930 2259.490 996.110 2260.670 ;
        RECT 994.930 2081.090 996.110 2082.270 ;
        RECT 994.930 2079.490 996.110 2080.670 ;
        RECT 994.930 1901.090 996.110 1902.270 ;
        RECT 994.930 1899.490 996.110 1900.670 ;
        RECT 994.930 1721.090 996.110 1722.270 ;
        RECT 994.930 1719.490 996.110 1720.670 ;
        RECT 994.930 1541.090 996.110 1542.270 ;
        RECT 994.930 1539.490 996.110 1540.670 ;
        RECT 994.930 1361.090 996.110 1362.270 ;
        RECT 994.930 1359.490 996.110 1360.670 ;
        RECT 994.930 1181.090 996.110 1182.270 ;
        RECT 994.930 1179.490 996.110 1180.670 ;
        RECT 994.930 1001.090 996.110 1002.270 ;
        RECT 994.930 999.490 996.110 1000.670 ;
        RECT 994.930 821.090 996.110 822.270 ;
        RECT 994.930 819.490 996.110 820.670 ;
        RECT 994.930 641.090 996.110 642.270 ;
        RECT 994.930 639.490 996.110 640.670 ;
        RECT 994.930 461.090 996.110 462.270 ;
        RECT 994.930 459.490 996.110 460.670 ;
        RECT 994.930 281.090 996.110 282.270 ;
        RECT 994.930 279.490 996.110 280.670 ;
        RECT 994.930 101.090 996.110 102.270 ;
        RECT 994.930 99.490 996.110 100.670 ;
        RECT 994.930 -7.510 996.110 -6.330 ;
        RECT 994.930 -9.110 996.110 -7.930 ;
        RECT 1174.930 3527.610 1176.110 3528.790 ;
        RECT 1174.930 3526.010 1176.110 3527.190 ;
        RECT 1174.930 3341.090 1176.110 3342.270 ;
        RECT 1174.930 3339.490 1176.110 3340.670 ;
        RECT 1174.930 3161.090 1176.110 3162.270 ;
        RECT 1174.930 3159.490 1176.110 3160.670 ;
        RECT 1174.930 2981.090 1176.110 2982.270 ;
        RECT 1174.930 2979.490 1176.110 2980.670 ;
        RECT 1174.930 2801.090 1176.110 2802.270 ;
        RECT 1174.930 2799.490 1176.110 2800.670 ;
        RECT 1174.930 2621.090 1176.110 2622.270 ;
        RECT 1174.930 2619.490 1176.110 2620.670 ;
        RECT 1174.930 2441.090 1176.110 2442.270 ;
        RECT 1174.930 2439.490 1176.110 2440.670 ;
        RECT 1174.930 2261.090 1176.110 2262.270 ;
        RECT 1174.930 2259.490 1176.110 2260.670 ;
        RECT 1174.930 2081.090 1176.110 2082.270 ;
        RECT 1174.930 2079.490 1176.110 2080.670 ;
        RECT 1174.930 1901.090 1176.110 1902.270 ;
        RECT 1174.930 1899.490 1176.110 1900.670 ;
        RECT 1174.930 1721.090 1176.110 1722.270 ;
        RECT 1174.930 1719.490 1176.110 1720.670 ;
        RECT 1174.930 1541.090 1176.110 1542.270 ;
        RECT 1174.930 1539.490 1176.110 1540.670 ;
        RECT 1174.930 1361.090 1176.110 1362.270 ;
        RECT 1174.930 1359.490 1176.110 1360.670 ;
        RECT 1174.930 1181.090 1176.110 1182.270 ;
        RECT 1174.930 1179.490 1176.110 1180.670 ;
        RECT 1174.930 1001.090 1176.110 1002.270 ;
        RECT 1174.930 999.490 1176.110 1000.670 ;
        RECT 1174.930 821.090 1176.110 822.270 ;
        RECT 1174.930 819.490 1176.110 820.670 ;
        RECT 1174.930 641.090 1176.110 642.270 ;
        RECT 1174.930 639.490 1176.110 640.670 ;
        RECT 1174.930 461.090 1176.110 462.270 ;
        RECT 1174.930 459.490 1176.110 460.670 ;
        RECT 1174.930 281.090 1176.110 282.270 ;
        RECT 1174.930 279.490 1176.110 280.670 ;
        RECT 1174.930 101.090 1176.110 102.270 ;
        RECT 1174.930 99.490 1176.110 100.670 ;
        RECT 1174.930 -7.510 1176.110 -6.330 ;
        RECT 1174.930 -9.110 1176.110 -7.930 ;
        RECT 1354.930 3527.610 1356.110 3528.790 ;
        RECT 1354.930 3526.010 1356.110 3527.190 ;
        RECT 1354.930 3341.090 1356.110 3342.270 ;
        RECT 1354.930 3339.490 1356.110 3340.670 ;
        RECT 1354.930 3161.090 1356.110 3162.270 ;
        RECT 1354.930 3159.490 1356.110 3160.670 ;
        RECT 1354.930 2981.090 1356.110 2982.270 ;
        RECT 1354.930 2979.490 1356.110 2980.670 ;
        RECT 1354.930 2801.090 1356.110 2802.270 ;
        RECT 1354.930 2799.490 1356.110 2800.670 ;
        RECT 1354.930 2621.090 1356.110 2622.270 ;
        RECT 1354.930 2619.490 1356.110 2620.670 ;
        RECT 1354.930 2441.090 1356.110 2442.270 ;
        RECT 1354.930 2439.490 1356.110 2440.670 ;
        RECT 1354.930 2261.090 1356.110 2262.270 ;
        RECT 1354.930 2259.490 1356.110 2260.670 ;
        RECT 1354.930 2081.090 1356.110 2082.270 ;
        RECT 1354.930 2079.490 1356.110 2080.670 ;
        RECT 1354.930 1901.090 1356.110 1902.270 ;
        RECT 1354.930 1899.490 1356.110 1900.670 ;
        RECT 1354.930 1721.090 1356.110 1722.270 ;
        RECT 1354.930 1719.490 1356.110 1720.670 ;
        RECT 1354.930 1541.090 1356.110 1542.270 ;
        RECT 1354.930 1539.490 1356.110 1540.670 ;
        RECT 1354.930 1361.090 1356.110 1362.270 ;
        RECT 1354.930 1359.490 1356.110 1360.670 ;
        RECT 1354.930 1181.090 1356.110 1182.270 ;
        RECT 1354.930 1179.490 1356.110 1180.670 ;
        RECT 1354.930 1001.090 1356.110 1002.270 ;
        RECT 1354.930 999.490 1356.110 1000.670 ;
        RECT 1354.930 821.090 1356.110 822.270 ;
        RECT 1354.930 819.490 1356.110 820.670 ;
        RECT 1354.930 641.090 1356.110 642.270 ;
        RECT 1354.930 639.490 1356.110 640.670 ;
        RECT 1354.930 461.090 1356.110 462.270 ;
        RECT 1354.930 459.490 1356.110 460.670 ;
        RECT 1354.930 281.090 1356.110 282.270 ;
        RECT 1354.930 279.490 1356.110 280.670 ;
        RECT 1354.930 101.090 1356.110 102.270 ;
        RECT 1354.930 99.490 1356.110 100.670 ;
        RECT 1354.930 -7.510 1356.110 -6.330 ;
        RECT 1354.930 -9.110 1356.110 -7.930 ;
        RECT 1534.930 3527.610 1536.110 3528.790 ;
        RECT 1534.930 3526.010 1536.110 3527.190 ;
        RECT 1534.930 3341.090 1536.110 3342.270 ;
        RECT 1534.930 3339.490 1536.110 3340.670 ;
        RECT 1534.930 3161.090 1536.110 3162.270 ;
        RECT 1534.930 3159.490 1536.110 3160.670 ;
        RECT 1534.930 2981.090 1536.110 2982.270 ;
        RECT 1534.930 2979.490 1536.110 2980.670 ;
        RECT 1534.930 2801.090 1536.110 2802.270 ;
        RECT 1534.930 2799.490 1536.110 2800.670 ;
        RECT 1534.930 2621.090 1536.110 2622.270 ;
        RECT 1534.930 2619.490 1536.110 2620.670 ;
        RECT 1534.930 2441.090 1536.110 2442.270 ;
        RECT 1534.930 2439.490 1536.110 2440.670 ;
        RECT 1534.930 2261.090 1536.110 2262.270 ;
        RECT 1534.930 2259.490 1536.110 2260.670 ;
        RECT 1534.930 2081.090 1536.110 2082.270 ;
        RECT 1534.930 2079.490 1536.110 2080.670 ;
        RECT 1534.930 1901.090 1536.110 1902.270 ;
        RECT 1534.930 1899.490 1536.110 1900.670 ;
        RECT 1534.930 1721.090 1536.110 1722.270 ;
        RECT 1534.930 1719.490 1536.110 1720.670 ;
        RECT 1534.930 1541.090 1536.110 1542.270 ;
        RECT 1534.930 1539.490 1536.110 1540.670 ;
        RECT 1534.930 1361.090 1536.110 1362.270 ;
        RECT 1534.930 1359.490 1536.110 1360.670 ;
        RECT 1534.930 1181.090 1536.110 1182.270 ;
        RECT 1534.930 1179.490 1536.110 1180.670 ;
        RECT 1534.930 1001.090 1536.110 1002.270 ;
        RECT 1534.930 999.490 1536.110 1000.670 ;
        RECT 1534.930 821.090 1536.110 822.270 ;
        RECT 1534.930 819.490 1536.110 820.670 ;
        RECT 1534.930 641.090 1536.110 642.270 ;
        RECT 1534.930 639.490 1536.110 640.670 ;
        RECT 1534.930 461.090 1536.110 462.270 ;
        RECT 1534.930 459.490 1536.110 460.670 ;
        RECT 1534.930 281.090 1536.110 282.270 ;
        RECT 1534.930 279.490 1536.110 280.670 ;
        RECT 1534.930 101.090 1536.110 102.270 ;
        RECT 1534.930 99.490 1536.110 100.670 ;
        RECT 1534.930 -7.510 1536.110 -6.330 ;
        RECT 1534.930 -9.110 1536.110 -7.930 ;
        RECT 1714.930 3527.610 1716.110 3528.790 ;
        RECT 1714.930 3526.010 1716.110 3527.190 ;
        RECT 1714.930 3341.090 1716.110 3342.270 ;
        RECT 1714.930 3339.490 1716.110 3340.670 ;
        RECT 1714.930 3161.090 1716.110 3162.270 ;
        RECT 1714.930 3159.490 1716.110 3160.670 ;
        RECT 1714.930 2981.090 1716.110 2982.270 ;
        RECT 1714.930 2979.490 1716.110 2980.670 ;
        RECT 1714.930 2801.090 1716.110 2802.270 ;
        RECT 1714.930 2799.490 1716.110 2800.670 ;
        RECT 1714.930 2621.090 1716.110 2622.270 ;
        RECT 1714.930 2619.490 1716.110 2620.670 ;
        RECT 1714.930 2441.090 1716.110 2442.270 ;
        RECT 1714.930 2439.490 1716.110 2440.670 ;
        RECT 1714.930 2261.090 1716.110 2262.270 ;
        RECT 1714.930 2259.490 1716.110 2260.670 ;
        RECT 1714.930 2081.090 1716.110 2082.270 ;
        RECT 1714.930 2079.490 1716.110 2080.670 ;
        RECT 1714.930 1901.090 1716.110 1902.270 ;
        RECT 1714.930 1899.490 1716.110 1900.670 ;
        RECT 1714.930 1721.090 1716.110 1722.270 ;
        RECT 1714.930 1719.490 1716.110 1720.670 ;
        RECT 1714.930 1541.090 1716.110 1542.270 ;
        RECT 1714.930 1539.490 1716.110 1540.670 ;
        RECT 1714.930 1361.090 1716.110 1362.270 ;
        RECT 1714.930 1359.490 1716.110 1360.670 ;
        RECT 1714.930 1181.090 1716.110 1182.270 ;
        RECT 1714.930 1179.490 1716.110 1180.670 ;
        RECT 1714.930 1001.090 1716.110 1002.270 ;
        RECT 1714.930 999.490 1716.110 1000.670 ;
        RECT 1714.930 821.090 1716.110 822.270 ;
        RECT 1714.930 819.490 1716.110 820.670 ;
        RECT 1714.930 641.090 1716.110 642.270 ;
        RECT 1714.930 639.490 1716.110 640.670 ;
        RECT 1714.930 461.090 1716.110 462.270 ;
        RECT 1714.930 459.490 1716.110 460.670 ;
        RECT 1714.930 281.090 1716.110 282.270 ;
        RECT 1714.930 279.490 1716.110 280.670 ;
        RECT 1714.930 101.090 1716.110 102.270 ;
        RECT 1714.930 99.490 1716.110 100.670 ;
        RECT 1714.930 -7.510 1716.110 -6.330 ;
        RECT 1714.930 -9.110 1716.110 -7.930 ;
        RECT 1894.930 3527.610 1896.110 3528.790 ;
        RECT 1894.930 3526.010 1896.110 3527.190 ;
        RECT 1894.930 3341.090 1896.110 3342.270 ;
        RECT 1894.930 3339.490 1896.110 3340.670 ;
        RECT 1894.930 3161.090 1896.110 3162.270 ;
        RECT 1894.930 3159.490 1896.110 3160.670 ;
        RECT 1894.930 2981.090 1896.110 2982.270 ;
        RECT 1894.930 2979.490 1896.110 2980.670 ;
        RECT 1894.930 2801.090 1896.110 2802.270 ;
        RECT 1894.930 2799.490 1896.110 2800.670 ;
        RECT 1894.930 2621.090 1896.110 2622.270 ;
        RECT 1894.930 2619.490 1896.110 2620.670 ;
        RECT 1894.930 2441.090 1896.110 2442.270 ;
        RECT 1894.930 2439.490 1896.110 2440.670 ;
        RECT 1894.930 2261.090 1896.110 2262.270 ;
        RECT 1894.930 2259.490 1896.110 2260.670 ;
        RECT 1894.930 2081.090 1896.110 2082.270 ;
        RECT 1894.930 2079.490 1896.110 2080.670 ;
        RECT 1894.930 1901.090 1896.110 1902.270 ;
        RECT 1894.930 1899.490 1896.110 1900.670 ;
        RECT 1894.930 1721.090 1896.110 1722.270 ;
        RECT 1894.930 1719.490 1896.110 1720.670 ;
        RECT 1894.930 1541.090 1896.110 1542.270 ;
        RECT 1894.930 1539.490 1896.110 1540.670 ;
        RECT 1894.930 1361.090 1896.110 1362.270 ;
        RECT 1894.930 1359.490 1896.110 1360.670 ;
        RECT 1894.930 1181.090 1896.110 1182.270 ;
        RECT 1894.930 1179.490 1896.110 1180.670 ;
        RECT 1894.930 1001.090 1896.110 1002.270 ;
        RECT 1894.930 999.490 1896.110 1000.670 ;
        RECT 1894.930 821.090 1896.110 822.270 ;
        RECT 1894.930 819.490 1896.110 820.670 ;
        RECT 1894.930 641.090 1896.110 642.270 ;
        RECT 1894.930 639.490 1896.110 640.670 ;
        RECT 1894.930 461.090 1896.110 462.270 ;
        RECT 1894.930 459.490 1896.110 460.670 ;
        RECT 1894.930 281.090 1896.110 282.270 ;
        RECT 1894.930 279.490 1896.110 280.670 ;
        RECT 1894.930 101.090 1896.110 102.270 ;
        RECT 1894.930 99.490 1896.110 100.670 ;
        RECT 1894.930 -7.510 1896.110 -6.330 ;
        RECT 1894.930 -9.110 1896.110 -7.930 ;
        RECT 2074.930 3527.610 2076.110 3528.790 ;
        RECT 2074.930 3526.010 2076.110 3527.190 ;
        RECT 2074.930 3341.090 2076.110 3342.270 ;
        RECT 2074.930 3339.490 2076.110 3340.670 ;
        RECT 2074.930 3161.090 2076.110 3162.270 ;
        RECT 2074.930 3159.490 2076.110 3160.670 ;
        RECT 2074.930 2981.090 2076.110 2982.270 ;
        RECT 2074.930 2979.490 2076.110 2980.670 ;
        RECT 2074.930 2801.090 2076.110 2802.270 ;
        RECT 2074.930 2799.490 2076.110 2800.670 ;
        RECT 2074.930 2621.090 2076.110 2622.270 ;
        RECT 2074.930 2619.490 2076.110 2620.670 ;
        RECT 2074.930 2441.090 2076.110 2442.270 ;
        RECT 2074.930 2439.490 2076.110 2440.670 ;
        RECT 2074.930 2261.090 2076.110 2262.270 ;
        RECT 2074.930 2259.490 2076.110 2260.670 ;
        RECT 2074.930 2081.090 2076.110 2082.270 ;
        RECT 2074.930 2079.490 2076.110 2080.670 ;
        RECT 2074.930 1901.090 2076.110 1902.270 ;
        RECT 2074.930 1899.490 2076.110 1900.670 ;
        RECT 2074.930 1721.090 2076.110 1722.270 ;
        RECT 2074.930 1719.490 2076.110 1720.670 ;
        RECT 2074.930 1541.090 2076.110 1542.270 ;
        RECT 2074.930 1539.490 2076.110 1540.670 ;
        RECT 2074.930 1361.090 2076.110 1362.270 ;
        RECT 2074.930 1359.490 2076.110 1360.670 ;
        RECT 2074.930 1181.090 2076.110 1182.270 ;
        RECT 2074.930 1179.490 2076.110 1180.670 ;
        RECT 2074.930 1001.090 2076.110 1002.270 ;
        RECT 2074.930 999.490 2076.110 1000.670 ;
        RECT 2074.930 821.090 2076.110 822.270 ;
        RECT 2074.930 819.490 2076.110 820.670 ;
        RECT 2074.930 641.090 2076.110 642.270 ;
        RECT 2074.930 639.490 2076.110 640.670 ;
        RECT 2074.930 461.090 2076.110 462.270 ;
        RECT 2074.930 459.490 2076.110 460.670 ;
        RECT 2074.930 281.090 2076.110 282.270 ;
        RECT 2074.930 279.490 2076.110 280.670 ;
        RECT 2074.930 101.090 2076.110 102.270 ;
        RECT 2074.930 99.490 2076.110 100.670 ;
        RECT 2074.930 -7.510 2076.110 -6.330 ;
        RECT 2074.930 -9.110 2076.110 -7.930 ;
        RECT 2254.930 3527.610 2256.110 3528.790 ;
        RECT 2254.930 3526.010 2256.110 3527.190 ;
        RECT 2254.930 3341.090 2256.110 3342.270 ;
        RECT 2254.930 3339.490 2256.110 3340.670 ;
        RECT 2254.930 3161.090 2256.110 3162.270 ;
        RECT 2254.930 3159.490 2256.110 3160.670 ;
        RECT 2254.930 2981.090 2256.110 2982.270 ;
        RECT 2254.930 2979.490 2256.110 2980.670 ;
        RECT 2254.930 2801.090 2256.110 2802.270 ;
        RECT 2254.930 2799.490 2256.110 2800.670 ;
        RECT 2254.930 2621.090 2256.110 2622.270 ;
        RECT 2254.930 2619.490 2256.110 2620.670 ;
        RECT 2254.930 2441.090 2256.110 2442.270 ;
        RECT 2254.930 2439.490 2256.110 2440.670 ;
        RECT 2254.930 2261.090 2256.110 2262.270 ;
        RECT 2254.930 2259.490 2256.110 2260.670 ;
        RECT 2254.930 2081.090 2256.110 2082.270 ;
        RECT 2254.930 2079.490 2256.110 2080.670 ;
        RECT 2254.930 1901.090 2256.110 1902.270 ;
        RECT 2254.930 1899.490 2256.110 1900.670 ;
        RECT 2254.930 1721.090 2256.110 1722.270 ;
        RECT 2254.930 1719.490 2256.110 1720.670 ;
        RECT 2254.930 1541.090 2256.110 1542.270 ;
        RECT 2254.930 1539.490 2256.110 1540.670 ;
        RECT 2254.930 1361.090 2256.110 1362.270 ;
        RECT 2254.930 1359.490 2256.110 1360.670 ;
        RECT 2254.930 1181.090 2256.110 1182.270 ;
        RECT 2254.930 1179.490 2256.110 1180.670 ;
        RECT 2254.930 1001.090 2256.110 1002.270 ;
        RECT 2254.930 999.490 2256.110 1000.670 ;
        RECT 2254.930 821.090 2256.110 822.270 ;
        RECT 2254.930 819.490 2256.110 820.670 ;
        RECT 2254.930 641.090 2256.110 642.270 ;
        RECT 2254.930 639.490 2256.110 640.670 ;
        RECT 2254.930 461.090 2256.110 462.270 ;
        RECT 2254.930 459.490 2256.110 460.670 ;
        RECT 2254.930 281.090 2256.110 282.270 ;
        RECT 2254.930 279.490 2256.110 280.670 ;
        RECT 2254.930 101.090 2256.110 102.270 ;
        RECT 2254.930 99.490 2256.110 100.670 ;
        RECT 2254.930 -7.510 2256.110 -6.330 ;
        RECT 2254.930 -9.110 2256.110 -7.930 ;
        RECT 2434.930 3527.610 2436.110 3528.790 ;
        RECT 2434.930 3526.010 2436.110 3527.190 ;
        RECT 2434.930 3341.090 2436.110 3342.270 ;
        RECT 2434.930 3339.490 2436.110 3340.670 ;
        RECT 2434.930 3161.090 2436.110 3162.270 ;
        RECT 2434.930 3159.490 2436.110 3160.670 ;
        RECT 2434.930 2981.090 2436.110 2982.270 ;
        RECT 2434.930 2979.490 2436.110 2980.670 ;
        RECT 2434.930 2801.090 2436.110 2802.270 ;
        RECT 2434.930 2799.490 2436.110 2800.670 ;
        RECT 2434.930 2621.090 2436.110 2622.270 ;
        RECT 2434.930 2619.490 2436.110 2620.670 ;
        RECT 2434.930 2441.090 2436.110 2442.270 ;
        RECT 2434.930 2439.490 2436.110 2440.670 ;
        RECT 2434.930 2261.090 2436.110 2262.270 ;
        RECT 2434.930 2259.490 2436.110 2260.670 ;
        RECT 2434.930 2081.090 2436.110 2082.270 ;
        RECT 2434.930 2079.490 2436.110 2080.670 ;
        RECT 2434.930 1901.090 2436.110 1902.270 ;
        RECT 2434.930 1899.490 2436.110 1900.670 ;
        RECT 2434.930 1721.090 2436.110 1722.270 ;
        RECT 2434.930 1719.490 2436.110 1720.670 ;
        RECT 2434.930 1541.090 2436.110 1542.270 ;
        RECT 2434.930 1539.490 2436.110 1540.670 ;
        RECT 2434.930 1361.090 2436.110 1362.270 ;
        RECT 2434.930 1359.490 2436.110 1360.670 ;
        RECT 2434.930 1181.090 2436.110 1182.270 ;
        RECT 2434.930 1179.490 2436.110 1180.670 ;
        RECT 2434.930 1001.090 2436.110 1002.270 ;
        RECT 2434.930 999.490 2436.110 1000.670 ;
        RECT 2434.930 821.090 2436.110 822.270 ;
        RECT 2434.930 819.490 2436.110 820.670 ;
        RECT 2434.930 641.090 2436.110 642.270 ;
        RECT 2434.930 639.490 2436.110 640.670 ;
        RECT 2434.930 461.090 2436.110 462.270 ;
        RECT 2434.930 459.490 2436.110 460.670 ;
        RECT 2434.930 281.090 2436.110 282.270 ;
        RECT 2434.930 279.490 2436.110 280.670 ;
        RECT 2434.930 101.090 2436.110 102.270 ;
        RECT 2434.930 99.490 2436.110 100.670 ;
        RECT 2434.930 -7.510 2436.110 -6.330 ;
        RECT 2434.930 -9.110 2436.110 -7.930 ;
        RECT 2614.930 3527.610 2616.110 3528.790 ;
        RECT 2614.930 3526.010 2616.110 3527.190 ;
        RECT 2614.930 3341.090 2616.110 3342.270 ;
        RECT 2614.930 3339.490 2616.110 3340.670 ;
        RECT 2614.930 3161.090 2616.110 3162.270 ;
        RECT 2614.930 3159.490 2616.110 3160.670 ;
        RECT 2614.930 2981.090 2616.110 2982.270 ;
        RECT 2614.930 2979.490 2616.110 2980.670 ;
        RECT 2614.930 2801.090 2616.110 2802.270 ;
        RECT 2614.930 2799.490 2616.110 2800.670 ;
        RECT 2614.930 2621.090 2616.110 2622.270 ;
        RECT 2614.930 2619.490 2616.110 2620.670 ;
        RECT 2614.930 2441.090 2616.110 2442.270 ;
        RECT 2614.930 2439.490 2616.110 2440.670 ;
        RECT 2614.930 2261.090 2616.110 2262.270 ;
        RECT 2614.930 2259.490 2616.110 2260.670 ;
        RECT 2614.930 2081.090 2616.110 2082.270 ;
        RECT 2614.930 2079.490 2616.110 2080.670 ;
        RECT 2614.930 1901.090 2616.110 1902.270 ;
        RECT 2614.930 1899.490 2616.110 1900.670 ;
        RECT 2614.930 1721.090 2616.110 1722.270 ;
        RECT 2614.930 1719.490 2616.110 1720.670 ;
        RECT 2614.930 1541.090 2616.110 1542.270 ;
        RECT 2614.930 1539.490 2616.110 1540.670 ;
        RECT 2614.930 1361.090 2616.110 1362.270 ;
        RECT 2614.930 1359.490 2616.110 1360.670 ;
        RECT 2614.930 1181.090 2616.110 1182.270 ;
        RECT 2614.930 1179.490 2616.110 1180.670 ;
        RECT 2614.930 1001.090 2616.110 1002.270 ;
        RECT 2614.930 999.490 2616.110 1000.670 ;
        RECT 2614.930 821.090 2616.110 822.270 ;
        RECT 2614.930 819.490 2616.110 820.670 ;
        RECT 2614.930 641.090 2616.110 642.270 ;
        RECT 2614.930 639.490 2616.110 640.670 ;
        RECT 2614.930 461.090 2616.110 462.270 ;
        RECT 2614.930 459.490 2616.110 460.670 ;
        RECT 2614.930 281.090 2616.110 282.270 ;
        RECT 2614.930 279.490 2616.110 280.670 ;
        RECT 2614.930 101.090 2616.110 102.270 ;
        RECT 2614.930 99.490 2616.110 100.670 ;
        RECT 2614.930 -7.510 2616.110 -6.330 ;
        RECT 2614.930 -9.110 2616.110 -7.930 ;
        RECT 2794.930 3527.610 2796.110 3528.790 ;
        RECT 2794.930 3526.010 2796.110 3527.190 ;
        RECT 2794.930 3341.090 2796.110 3342.270 ;
        RECT 2794.930 3339.490 2796.110 3340.670 ;
        RECT 2794.930 3161.090 2796.110 3162.270 ;
        RECT 2794.930 3159.490 2796.110 3160.670 ;
        RECT 2794.930 2981.090 2796.110 2982.270 ;
        RECT 2794.930 2979.490 2796.110 2980.670 ;
        RECT 2794.930 2801.090 2796.110 2802.270 ;
        RECT 2794.930 2799.490 2796.110 2800.670 ;
        RECT 2794.930 2621.090 2796.110 2622.270 ;
        RECT 2794.930 2619.490 2796.110 2620.670 ;
        RECT 2794.930 2441.090 2796.110 2442.270 ;
        RECT 2794.930 2439.490 2796.110 2440.670 ;
        RECT 2794.930 2261.090 2796.110 2262.270 ;
        RECT 2794.930 2259.490 2796.110 2260.670 ;
        RECT 2794.930 2081.090 2796.110 2082.270 ;
        RECT 2794.930 2079.490 2796.110 2080.670 ;
        RECT 2794.930 1901.090 2796.110 1902.270 ;
        RECT 2794.930 1899.490 2796.110 1900.670 ;
        RECT 2794.930 1721.090 2796.110 1722.270 ;
        RECT 2794.930 1719.490 2796.110 1720.670 ;
        RECT 2794.930 1541.090 2796.110 1542.270 ;
        RECT 2794.930 1539.490 2796.110 1540.670 ;
        RECT 2794.930 1361.090 2796.110 1362.270 ;
        RECT 2794.930 1359.490 2796.110 1360.670 ;
        RECT 2794.930 1181.090 2796.110 1182.270 ;
        RECT 2794.930 1179.490 2796.110 1180.670 ;
        RECT 2794.930 1001.090 2796.110 1002.270 ;
        RECT 2794.930 999.490 2796.110 1000.670 ;
        RECT 2794.930 821.090 2796.110 822.270 ;
        RECT 2794.930 819.490 2796.110 820.670 ;
        RECT 2794.930 641.090 2796.110 642.270 ;
        RECT 2794.930 639.490 2796.110 640.670 ;
        RECT 2794.930 461.090 2796.110 462.270 ;
        RECT 2794.930 459.490 2796.110 460.670 ;
        RECT 2794.930 281.090 2796.110 282.270 ;
        RECT 2794.930 279.490 2796.110 280.670 ;
        RECT 2794.930 101.090 2796.110 102.270 ;
        RECT 2794.930 99.490 2796.110 100.670 ;
        RECT 2794.930 -7.510 2796.110 -6.330 ;
        RECT 2794.930 -9.110 2796.110 -7.930 ;
        RECT 2932.110 3527.610 2933.290 3528.790 ;
        RECT 2932.110 3526.010 2933.290 3527.190 ;
        RECT 2932.110 3341.090 2933.290 3342.270 ;
        RECT 2932.110 3339.490 2933.290 3340.670 ;
        RECT 2932.110 3161.090 2933.290 3162.270 ;
        RECT 2932.110 3159.490 2933.290 3160.670 ;
        RECT 2932.110 2981.090 2933.290 2982.270 ;
        RECT 2932.110 2979.490 2933.290 2980.670 ;
        RECT 2932.110 2801.090 2933.290 2802.270 ;
        RECT 2932.110 2799.490 2933.290 2800.670 ;
        RECT 2932.110 2621.090 2933.290 2622.270 ;
        RECT 2932.110 2619.490 2933.290 2620.670 ;
        RECT 2932.110 2441.090 2933.290 2442.270 ;
        RECT 2932.110 2439.490 2933.290 2440.670 ;
        RECT 2932.110 2261.090 2933.290 2262.270 ;
        RECT 2932.110 2259.490 2933.290 2260.670 ;
        RECT 2932.110 2081.090 2933.290 2082.270 ;
        RECT 2932.110 2079.490 2933.290 2080.670 ;
        RECT 2932.110 1901.090 2933.290 1902.270 ;
        RECT 2932.110 1899.490 2933.290 1900.670 ;
        RECT 2932.110 1721.090 2933.290 1722.270 ;
        RECT 2932.110 1719.490 2933.290 1720.670 ;
        RECT 2932.110 1541.090 2933.290 1542.270 ;
        RECT 2932.110 1539.490 2933.290 1540.670 ;
        RECT 2932.110 1361.090 2933.290 1362.270 ;
        RECT 2932.110 1359.490 2933.290 1360.670 ;
        RECT 2932.110 1181.090 2933.290 1182.270 ;
        RECT 2932.110 1179.490 2933.290 1180.670 ;
        RECT 2932.110 1001.090 2933.290 1002.270 ;
        RECT 2932.110 999.490 2933.290 1000.670 ;
        RECT 2932.110 821.090 2933.290 822.270 ;
        RECT 2932.110 819.490 2933.290 820.670 ;
        RECT 2932.110 641.090 2933.290 642.270 ;
        RECT 2932.110 639.490 2933.290 640.670 ;
        RECT 2932.110 461.090 2933.290 462.270 ;
        RECT 2932.110 459.490 2933.290 460.670 ;
        RECT 2932.110 281.090 2933.290 282.270 ;
        RECT 2932.110 279.490 2933.290 280.670 ;
        RECT 2932.110 101.090 2933.290 102.270 ;
        RECT 2932.110 99.490 2933.290 100.670 ;
        RECT 2932.110 -7.510 2933.290 -6.330 ;
        RECT 2932.110 -9.110 2933.290 -7.930 ;
      LAYER met5 ;
        RECT -14.580 3528.900 -11.580 3528.910 ;
        RECT 94.020 3528.900 97.020 3528.910 ;
        RECT 274.020 3528.900 277.020 3528.910 ;
        RECT 454.020 3528.900 457.020 3528.910 ;
        RECT 634.020 3528.900 637.020 3528.910 ;
        RECT 814.020 3528.900 817.020 3528.910 ;
        RECT 994.020 3528.900 997.020 3528.910 ;
        RECT 1174.020 3528.900 1177.020 3528.910 ;
        RECT 1354.020 3528.900 1357.020 3528.910 ;
        RECT 1534.020 3528.900 1537.020 3528.910 ;
        RECT 1714.020 3528.900 1717.020 3528.910 ;
        RECT 1894.020 3528.900 1897.020 3528.910 ;
        RECT 2074.020 3528.900 2077.020 3528.910 ;
        RECT 2254.020 3528.900 2257.020 3528.910 ;
        RECT 2434.020 3528.900 2437.020 3528.910 ;
        RECT 2614.020 3528.900 2617.020 3528.910 ;
        RECT 2794.020 3528.900 2797.020 3528.910 ;
        RECT 2931.200 3528.900 2934.200 3528.910 ;
        RECT -14.580 3525.900 2934.200 3528.900 ;
        RECT -14.580 3525.890 -11.580 3525.900 ;
        RECT 94.020 3525.890 97.020 3525.900 ;
        RECT 274.020 3525.890 277.020 3525.900 ;
        RECT 454.020 3525.890 457.020 3525.900 ;
        RECT 634.020 3525.890 637.020 3525.900 ;
        RECT 814.020 3525.890 817.020 3525.900 ;
        RECT 994.020 3525.890 997.020 3525.900 ;
        RECT 1174.020 3525.890 1177.020 3525.900 ;
        RECT 1354.020 3525.890 1357.020 3525.900 ;
        RECT 1534.020 3525.890 1537.020 3525.900 ;
        RECT 1714.020 3525.890 1717.020 3525.900 ;
        RECT 1894.020 3525.890 1897.020 3525.900 ;
        RECT 2074.020 3525.890 2077.020 3525.900 ;
        RECT 2254.020 3525.890 2257.020 3525.900 ;
        RECT 2434.020 3525.890 2437.020 3525.900 ;
        RECT 2614.020 3525.890 2617.020 3525.900 ;
        RECT 2794.020 3525.890 2797.020 3525.900 ;
        RECT 2931.200 3525.890 2934.200 3525.900 ;
        RECT -14.580 3342.380 -11.580 3342.390 ;
        RECT 94.020 3342.380 97.020 3342.390 ;
        RECT 274.020 3342.380 277.020 3342.390 ;
        RECT 454.020 3342.380 457.020 3342.390 ;
        RECT 634.020 3342.380 637.020 3342.390 ;
        RECT 814.020 3342.380 817.020 3342.390 ;
        RECT 994.020 3342.380 997.020 3342.390 ;
        RECT 1174.020 3342.380 1177.020 3342.390 ;
        RECT 1354.020 3342.380 1357.020 3342.390 ;
        RECT 1534.020 3342.380 1537.020 3342.390 ;
        RECT 1714.020 3342.380 1717.020 3342.390 ;
        RECT 1894.020 3342.380 1897.020 3342.390 ;
        RECT 2074.020 3342.380 2077.020 3342.390 ;
        RECT 2254.020 3342.380 2257.020 3342.390 ;
        RECT 2434.020 3342.380 2437.020 3342.390 ;
        RECT 2614.020 3342.380 2617.020 3342.390 ;
        RECT 2794.020 3342.380 2797.020 3342.390 ;
        RECT 2931.200 3342.380 2934.200 3342.390 ;
        RECT -14.580 3339.380 2934.200 3342.380 ;
        RECT -14.580 3339.370 -11.580 3339.380 ;
        RECT 94.020 3339.370 97.020 3339.380 ;
        RECT 274.020 3339.370 277.020 3339.380 ;
        RECT 454.020 3339.370 457.020 3339.380 ;
        RECT 634.020 3339.370 637.020 3339.380 ;
        RECT 814.020 3339.370 817.020 3339.380 ;
        RECT 994.020 3339.370 997.020 3339.380 ;
        RECT 1174.020 3339.370 1177.020 3339.380 ;
        RECT 1354.020 3339.370 1357.020 3339.380 ;
        RECT 1534.020 3339.370 1537.020 3339.380 ;
        RECT 1714.020 3339.370 1717.020 3339.380 ;
        RECT 1894.020 3339.370 1897.020 3339.380 ;
        RECT 2074.020 3339.370 2077.020 3339.380 ;
        RECT 2254.020 3339.370 2257.020 3339.380 ;
        RECT 2434.020 3339.370 2437.020 3339.380 ;
        RECT 2614.020 3339.370 2617.020 3339.380 ;
        RECT 2794.020 3339.370 2797.020 3339.380 ;
        RECT 2931.200 3339.370 2934.200 3339.380 ;
        RECT -14.580 3162.380 -11.580 3162.390 ;
        RECT 94.020 3162.380 97.020 3162.390 ;
        RECT 274.020 3162.380 277.020 3162.390 ;
        RECT 454.020 3162.380 457.020 3162.390 ;
        RECT 634.020 3162.380 637.020 3162.390 ;
        RECT 814.020 3162.380 817.020 3162.390 ;
        RECT 994.020 3162.380 997.020 3162.390 ;
        RECT 1174.020 3162.380 1177.020 3162.390 ;
        RECT 1354.020 3162.380 1357.020 3162.390 ;
        RECT 1534.020 3162.380 1537.020 3162.390 ;
        RECT 1714.020 3162.380 1717.020 3162.390 ;
        RECT 1894.020 3162.380 1897.020 3162.390 ;
        RECT 2074.020 3162.380 2077.020 3162.390 ;
        RECT 2254.020 3162.380 2257.020 3162.390 ;
        RECT 2434.020 3162.380 2437.020 3162.390 ;
        RECT 2614.020 3162.380 2617.020 3162.390 ;
        RECT 2794.020 3162.380 2797.020 3162.390 ;
        RECT 2931.200 3162.380 2934.200 3162.390 ;
        RECT -14.580 3159.380 2934.200 3162.380 ;
        RECT -14.580 3159.370 -11.580 3159.380 ;
        RECT 94.020 3159.370 97.020 3159.380 ;
        RECT 274.020 3159.370 277.020 3159.380 ;
        RECT 454.020 3159.370 457.020 3159.380 ;
        RECT 634.020 3159.370 637.020 3159.380 ;
        RECT 814.020 3159.370 817.020 3159.380 ;
        RECT 994.020 3159.370 997.020 3159.380 ;
        RECT 1174.020 3159.370 1177.020 3159.380 ;
        RECT 1354.020 3159.370 1357.020 3159.380 ;
        RECT 1534.020 3159.370 1537.020 3159.380 ;
        RECT 1714.020 3159.370 1717.020 3159.380 ;
        RECT 1894.020 3159.370 1897.020 3159.380 ;
        RECT 2074.020 3159.370 2077.020 3159.380 ;
        RECT 2254.020 3159.370 2257.020 3159.380 ;
        RECT 2434.020 3159.370 2437.020 3159.380 ;
        RECT 2614.020 3159.370 2617.020 3159.380 ;
        RECT 2794.020 3159.370 2797.020 3159.380 ;
        RECT 2931.200 3159.370 2934.200 3159.380 ;
        RECT -14.580 2982.380 -11.580 2982.390 ;
        RECT 94.020 2982.380 97.020 2982.390 ;
        RECT 274.020 2982.380 277.020 2982.390 ;
        RECT 454.020 2982.380 457.020 2982.390 ;
        RECT 634.020 2982.380 637.020 2982.390 ;
        RECT 814.020 2982.380 817.020 2982.390 ;
        RECT 994.020 2982.380 997.020 2982.390 ;
        RECT 1174.020 2982.380 1177.020 2982.390 ;
        RECT 1354.020 2982.380 1357.020 2982.390 ;
        RECT 1534.020 2982.380 1537.020 2982.390 ;
        RECT 1714.020 2982.380 1717.020 2982.390 ;
        RECT 1894.020 2982.380 1897.020 2982.390 ;
        RECT 2074.020 2982.380 2077.020 2982.390 ;
        RECT 2254.020 2982.380 2257.020 2982.390 ;
        RECT 2434.020 2982.380 2437.020 2982.390 ;
        RECT 2614.020 2982.380 2617.020 2982.390 ;
        RECT 2794.020 2982.380 2797.020 2982.390 ;
        RECT 2931.200 2982.380 2934.200 2982.390 ;
        RECT -14.580 2979.380 2934.200 2982.380 ;
        RECT -14.580 2979.370 -11.580 2979.380 ;
        RECT 94.020 2979.370 97.020 2979.380 ;
        RECT 274.020 2979.370 277.020 2979.380 ;
        RECT 454.020 2979.370 457.020 2979.380 ;
        RECT 634.020 2979.370 637.020 2979.380 ;
        RECT 814.020 2979.370 817.020 2979.380 ;
        RECT 994.020 2979.370 997.020 2979.380 ;
        RECT 1174.020 2979.370 1177.020 2979.380 ;
        RECT 1354.020 2979.370 1357.020 2979.380 ;
        RECT 1534.020 2979.370 1537.020 2979.380 ;
        RECT 1714.020 2979.370 1717.020 2979.380 ;
        RECT 1894.020 2979.370 1897.020 2979.380 ;
        RECT 2074.020 2979.370 2077.020 2979.380 ;
        RECT 2254.020 2979.370 2257.020 2979.380 ;
        RECT 2434.020 2979.370 2437.020 2979.380 ;
        RECT 2614.020 2979.370 2617.020 2979.380 ;
        RECT 2794.020 2979.370 2797.020 2979.380 ;
        RECT 2931.200 2979.370 2934.200 2979.380 ;
        RECT -14.580 2802.380 -11.580 2802.390 ;
        RECT 94.020 2802.380 97.020 2802.390 ;
        RECT 274.020 2802.380 277.020 2802.390 ;
        RECT 454.020 2802.380 457.020 2802.390 ;
        RECT 634.020 2802.380 637.020 2802.390 ;
        RECT 814.020 2802.380 817.020 2802.390 ;
        RECT 994.020 2802.380 997.020 2802.390 ;
        RECT 1174.020 2802.380 1177.020 2802.390 ;
        RECT 1354.020 2802.380 1357.020 2802.390 ;
        RECT 1534.020 2802.380 1537.020 2802.390 ;
        RECT 1714.020 2802.380 1717.020 2802.390 ;
        RECT 1894.020 2802.380 1897.020 2802.390 ;
        RECT 2074.020 2802.380 2077.020 2802.390 ;
        RECT 2254.020 2802.380 2257.020 2802.390 ;
        RECT 2434.020 2802.380 2437.020 2802.390 ;
        RECT 2614.020 2802.380 2617.020 2802.390 ;
        RECT 2794.020 2802.380 2797.020 2802.390 ;
        RECT 2931.200 2802.380 2934.200 2802.390 ;
        RECT -14.580 2799.380 2934.200 2802.380 ;
        RECT -14.580 2799.370 -11.580 2799.380 ;
        RECT 94.020 2799.370 97.020 2799.380 ;
        RECT 274.020 2799.370 277.020 2799.380 ;
        RECT 454.020 2799.370 457.020 2799.380 ;
        RECT 634.020 2799.370 637.020 2799.380 ;
        RECT 814.020 2799.370 817.020 2799.380 ;
        RECT 994.020 2799.370 997.020 2799.380 ;
        RECT 1174.020 2799.370 1177.020 2799.380 ;
        RECT 1354.020 2799.370 1357.020 2799.380 ;
        RECT 1534.020 2799.370 1537.020 2799.380 ;
        RECT 1714.020 2799.370 1717.020 2799.380 ;
        RECT 1894.020 2799.370 1897.020 2799.380 ;
        RECT 2074.020 2799.370 2077.020 2799.380 ;
        RECT 2254.020 2799.370 2257.020 2799.380 ;
        RECT 2434.020 2799.370 2437.020 2799.380 ;
        RECT 2614.020 2799.370 2617.020 2799.380 ;
        RECT 2794.020 2799.370 2797.020 2799.380 ;
        RECT 2931.200 2799.370 2934.200 2799.380 ;
        RECT -14.580 2622.380 -11.580 2622.390 ;
        RECT 94.020 2622.380 97.020 2622.390 ;
        RECT 274.020 2622.380 277.020 2622.390 ;
        RECT 454.020 2622.380 457.020 2622.390 ;
        RECT 634.020 2622.380 637.020 2622.390 ;
        RECT 814.020 2622.380 817.020 2622.390 ;
        RECT 994.020 2622.380 997.020 2622.390 ;
        RECT 1174.020 2622.380 1177.020 2622.390 ;
        RECT 1354.020 2622.380 1357.020 2622.390 ;
        RECT 1534.020 2622.380 1537.020 2622.390 ;
        RECT 1714.020 2622.380 1717.020 2622.390 ;
        RECT 1894.020 2622.380 1897.020 2622.390 ;
        RECT 2074.020 2622.380 2077.020 2622.390 ;
        RECT 2254.020 2622.380 2257.020 2622.390 ;
        RECT 2434.020 2622.380 2437.020 2622.390 ;
        RECT 2614.020 2622.380 2617.020 2622.390 ;
        RECT 2794.020 2622.380 2797.020 2622.390 ;
        RECT 2931.200 2622.380 2934.200 2622.390 ;
        RECT -14.580 2619.380 2934.200 2622.380 ;
        RECT -14.580 2619.370 -11.580 2619.380 ;
        RECT 94.020 2619.370 97.020 2619.380 ;
        RECT 274.020 2619.370 277.020 2619.380 ;
        RECT 454.020 2619.370 457.020 2619.380 ;
        RECT 634.020 2619.370 637.020 2619.380 ;
        RECT 814.020 2619.370 817.020 2619.380 ;
        RECT 994.020 2619.370 997.020 2619.380 ;
        RECT 1174.020 2619.370 1177.020 2619.380 ;
        RECT 1354.020 2619.370 1357.020 2619.380 ;
        RECT 1534.020 2619.370 1537.020 2619.380 ;
        RECT 1714.020 2619.370 1717.020 2619.380 ;
        RECT 1894.020 2619.370 1897.020 2619.380 ;
        RECT 2074.020 2619.370 2077.020 2619.380 ;
        RECT 2254.020 2619.370 2257.020 2619.380 ;
        RECT 2434.020 2619.370 2437.020 2619.380 ;
        RECT 2614.020 2619.370 2617.020 2619.380 ;
        RECT 2794.020 2619.370 2797.020 2619.380 ;
        RECT 2931.200 2619.370 2934.200 2619.380 ;
        RECT -14.580 2442.380 -11.580 2442.390 ;
        RECT 94.020 2442.380 97.020 2442.390 ;
        RECT 274.020 2442.380 277.020 2442.390 ;
        RECT 454.020 2442.380 457.020 2442.390 ;
        RECT 634.020 2442.380 637.020 2442.390 ;
        RECT 814.020 2442.380 817.020 2442.390 ;
        RECT 994.020 2442.380 997.020 2442.390 ;
        RECT 1174.020 2442.380 1177.020 2442.390 ;
        RECT 1354.020 2442.380 1357.020 2442.390 ;
        RECT 1534.020 2442.380 1537.020 2442.390 ;
        RECT 1714.020 2442.380 1717.020 2442.390 ;
        RECT 1894.020 2442.380 1897.020 2442.390 ;
        RECT 2074.020 2442.380 2077.020 2442.390 ;
        RECT 2254.020 2442.380 2257.020 2442.390 ;
        RECT 2434.020 2442.380 2437.020 2442.390 ;
        RECT 2614.020 2442.380 2617.020 2442.390 ;
        RECT 2794.020 2442.380 2797.020 2442.390 ;
        RECT 2931.200 2442.380 2934.200 2442.390 ;
        RECT -14.580 2439.380 2934.200 2442.380 ;
        RECT -14.580 2439.370 -11.580 2439.380 ;
        RECT 94.020 2439.370 97.020 2439.380 ;
        RECT 274.020 2439.370 277.020 2439.380 ;
        RECT 454.020 2439.370 457.020 2439.380 ;
        RECT 634.020 2439.370 637.020 2439.380 ;
        RECT 814.020 2439.370 817.020 2439.380 ;
        RECT 994.020 2439.370 997.020 2439.380 ;
        RECT 1174.020 2439.370 1177.020 2439.380 ;
        RECT 1354.020 2439.370 1357.020 2439.380 ;
        RECT 1534.020 2439.370 1537.020 2439.380 ;
        RECT 1714.020 2439.370 1717.020 2439.380 ;
        RECT 1894.020 2439.370 1897.020 2439.380 ;
        RECT 2074.020 2439.370 2077.020 2439.380 ;
        RECT 2254.020 2439.370 2257.020 2439.380 ;
        RECT 2434.020 2439.370 2437.020 2439.380 ;
        RECT 2614.020 2439.370 2617.020 2439.380 ;
        RECT 2794.020 2439.370 2797.020 2439.380 ;
        RECT 2931.200 2439.370 2934.200 2439.380 ;
        RECT -14.580 2262.380 -11.580 2262.390 ;
        RECT 94.020 2262.380 97.020 2262.390 ;
        RECT 274.020 2262.380 277.020 2262.390 ;
        RECT 454.020 2262.380 457.020 2262.390 ;
        RECT 634.020 2262.380 637.020 2262.390 ;
        RECT 814.020 2262.380 817.020 2262.390 ;
        RECT 994.020 2262.380 997.020 2262.390 ;
        RECT 1174.020 2262.380 1177.020 2262.390 ;
        RECT 1354.020 2262.380 1357.020 2262.390 ;
        RECT 1534.020 2262.380 1537.020 2262.390 ;
        RECT 1714.020 2262.380 1717.020 2262.390 ;
        RECT 1894.020 2262.380 1897.020 2262.390 ;
        RECT 2074.020 2262.380 2077.020 2262.390 ;
        RECT 2254.020 2262.380 2257.020 2262.390 ;
        RECT 2434.020 2262.380 2437.020 2262.390 ;
        RECT 2614.020 2262.380 2617.020 2262.390 ;
        RECT 2794.020 2262.380 2797.020 2262.390 ;
        RECT 2931.200 2262.380 2934.200 2262.390 ;
        RECT -14.580 2259.380 2934.200 2262.380 ;
        RECT -14.580 2259.370 -11.580 2259.380 ;
        RECT 94.020 2259.370 97.020 2259.380 ;
        RECT 274.020 2259.370 277.020 2259.380 ;
        RECT 454.020 2259.370 457.020 2259.380 ;
        RECT 634.020 2259.370 637.020 2259.380 ;
        RECT 814.020 2259.370 817.020 2259.380 ;
        RECT 994.020 2259.370 997.020 2259.380 ;
        RECT 1174.020 2259.370 1177.020 2259.380 ;
        RECT 1354.020 2259.370 1357.020 2259.380 ;
        RECT 1534.020 2259.370 1537.020 2259.380 ;
        RECT 1714.020 2259.370 1717.020 2259.380 ;
        RECT 1894.020 2259.370 1897.020 2259.380 ;
        RECT 2074.020 2259.370 2077.020 2259.380 ;
        RECT 2254.020 2259.370 2257.020 2259.380 ;
        RECT 2434.020 2259.370 2437.020 2259.380 ;
        RECT 2614.020 2259.370 2617.020 2259.380 ;
        RECT 2794.020 2259.370 2797.020 2259.380 ;
        RECT 2931.200 2259.370 2934.200 2259.380 ;
        RECT -14.580 2082.380 -11.580 2082.390 ;
        RECT 94.020 2082.380 97.020 2082.390 ;
        RECT 274.020 2082.380 277.020 2082.390 ;
        RECT 454.020 2082.380 457.020 2082.390 ;
        RECT 634.020 2082.380 637.020 2082.390 ;
        RECT 814.020 2082.380 817.020 2082.390 ;
        RECT 994.020 2082.380 997.020 2082.390 ;
        RECT 1174.020 2082.380 1177.020 2082.390 ;
        RECT 1354.020 2082.380 1357.020 2082.390 ;
        RECT 1534.020 2082.380 1537.020 2082.390 ;
        RECT 1714.020 2082.380 1717.020 2082.390 ;
        RECT 1894.020 2082.380 1897.020 2082.390 ;
        RECT 2074.020 2082.380 2077.020 2082.390 ;
        RECT 2254.020 2082.380 2257.020 2082.390 ;
        RECT 2434.020 2082.380 2437.020 2082.390 ;
        RECT 2614.020 2082.380 2617.020 2082.390 ;
        RECT 2794.020 2082.380 2797.020 2082.390 ;
        RECT 2931.200 2082.380 2934.200 2082.390 ;
        RECT -14.580 2079.380 2934.200 2082.380 ;
        RECT -14.580 2079.370 -11.580 2079.380 ;
        RECT 94.020 2079.370 97.020 2079.380 ;
        RECT 274.020 2079.370 277.020 2079.380 ;
        RECT 454.020 2079.370 457.020 2079.380 ;
        RECT 634.020 2079.370 637.020 2079.380 ;
        RECT 814.020 2079.370 817.020 2079.380 ;
        RECT 994.020 2079.370 997.020 2079.380 ;
        RECT 1174.020 2079.370 1177.020 2079.380 ;
        RECT 1354.020 2079.370 1357.020 2079.380 ;
        RECT 1534.020 2079.370 1537.020 2079.380 ;
        RECT 1714.020 2079.370 1717.020 2079.380 ;
        RECT 1894.020 2079.370 1897.020 2079.380 ;
        RECT 2074.020 2079.370 2077.020 2079.380 ;
        RECT 2254.020 2079.370 2257.020 2079.380 ;
        RECT 2434.020 2079.370 2437.020 2079.380 ;
        RECT 2614.020 2079.370 2617.020 2079.380 ;
        RECT 2794.020 2079.370 2797.020 2079.380 ;
        RECT 2931.200 2079.370 2934.200 2079.380 ;
        RECT -14.580 1902.380 -11.580 1902.390 ;
        RECT 94.020 1902.380 97.020 1902.390 ;
        RECT 274.020 1902.380 277.020 1902.390 ;
        RECT 454.020 1902.380 457.020 1902.390 ;
        RECT 634.020 1902.380 637.020 1902.390 ;
        RECT 814.020 1902.380 817.020 1902.390 ;
        RECT 994.020 1902.380 997.020 1902.390 ;
        RECT 1174.020 1902.380 1177.020 1902.390 ;
        RECT 1354.020 1902.380 1357.020 1902.390 ;
        RECT 1534.020 1902.380 1537.020 1902.390 ;
        RECT 1714.020 1902.380 1717.020 1902.390 ;
        RECT 1894.020 1902.380 1897.020 1902.390 ;
        RECT 2074.020 1902.380 2077.020 1902.390 ;
        RECT 2254.020 1902.380 2257.020 1902.390 ;
        RECT 2434.020 1902.380 2437.020 1902.390 ;
        RECT 2614.020 1902.380 2617.020 1902.390 ;
        RECT 2794.020 1902.380 2797.020 1902.390 ;
        RECT 2931.200 1902.380 2934.200 1902.390 ;
        RECT -14.580 1899.380 2934.200 1902.380 ;
        RECT -14.580 1899.370 -11.580 1899.380 ;
        RECT 94.020 1899.370 97.020 1899.380 ;
        RECT 274.020 1899.370 277.020 1899.380 ;
        RECT 454.020 1899.370 457.020 1899.380 ;
        RECT 634.020 1899.370 637.020 1899.380 ;
        RECT 814.020 1899.370 817.020 1899.380 ;
        RECT 994.020 1899.370 997.020 1899.380 ;
        RECT 1174.020 1899.370 1177.020 1899.380 ;
        RECT 1354.020 1899.370 1357.020 1899.380 ;
        RECT 1534.020 1899.370 1537.020 1899.380 ;
        RECT 1714.020 1899.370 1717.020 1899.380 ;
        RECT 1894.020 1899.370 1897.020 1899.380 ;
        RECT 2074.020 1899.370 2077.020 1899.380 ;
        RECT 2254.020 1899.370 2257.020 1899.380 ;
        RECT 2434.020 1899.370 2437.020 1899.380 ;
        RECT 2614.020 1899.370 2617.020 1899.380 ;
        RECT 2794.020 1899.370 2797.020 1899.380 ;
        RECT 2931.200 1899.370 2934.200 1899.380 ;
        RECT -14.580 1722.380 -11.580 1722.390 ;
        RECT 94.020 1722.380 97.020 1722.390 ;
        RECT 274.020 1722.380 277.020 1722.390 ;
        RECT 454.020 1722.380 457.020 1722.390 ;
        RECT 634.020 1722.380 637.020 1722.390 ;
        RECT 814.020 1722.380 817.020 1722.390 ;
        RECT 994.020 1722.380 997.020 1722.390 ;
        RECT 1174.020 1722.380 1177.020 1722.390 ;
        RECT 1354.020 1722.380 1357.020 1722.390 ;
        RECT 1534.020 1722.380 1537.020 1722.390 ;
        RECT 1714.020 1722.380 1717.020 1722.390 ;
        RECT 1894.020 1722.380 1897.020 1722.390 ;
        RECT 2074.020 1722.380 2077.020 1722.390 ;
        RECT 2254.020 1722.380 2257.020 1722.390 ;
        RECT 2434.020 1722.380 2437.020 1722.390 ;
        RECT 2614.020 1722.380 2617.020 1722.390 ;
        RECT 2794.020 1722.380 2797.020 1722.390 ;
        RECT 2931.200 1722.380 2934.200 1722.390 ;
        RECT -14.580 1719.380 2934.200 1722.380 ;
        RECT -14.580 1719.370 -11.580 1719.380 ;
        RECT 94.020 1719.370 97.020 1719.380 ;
        RECT 274.020 1719.370 277.020 1719.380 ;
        RECT 454.020 1719.370 457.020 1719.380 ;
        RECT 634.020 1719.370 637.020 1719.380 ;
        RECT 814.020 1719.370 817.020 1719.380 ;
        RECT 994.020 1719.370 997.020 1719.380 ;
        RECT 1174.020 1719.370 1177.020 1719.380 ;
        RECT 1354.020 1719.370 1357.020 1719.380 ;
        RECT 1534.020 1719.370 1537.020 1719.380 ;
        RECT 1714.020 1719.370 1717.020 1719.380 ;
        RECT 1894.020 1719.370 1897.020 1719.380 ;
        RECT 2074.020 1719.370 2077.020 1719.380 ;
        RECT 2254.020 1719.370 2257.020 1719.380 ;
        RECT 2434.020 1719.370 2437.020 1719.380 ;
        RECT 2614.020 1719.370 2617.020 1719.380 ;
        RECT 2794.020 1719.370 2797.020 1719.380 ;
        RECT 2931.200 1719.370 2934.200 1719.380 ;
        RECT -14.580 1542.380 -11.580 1542.390 ;
        RECT 94.020 1542.380 97.020 1542.390 ;
        RECT 274.020 1542.380 277.020 1542.390 ;
        RECT 454.020 1542.380 457.020 1542.390 ;
        RECT 634.020 1542.380 637.020 1542.390 ;
        RECT 814.020 1542.380 817.020 1542.390 ;
        RECT 994.020 1542.380 997.020 1542.390 ;
        RECT 1174.020 1542.380 1177.020 1542.390 ;
        RECT 1354.020 1542.380 1357.020 1542.390 ;
        RECT 1534.020 1542.380 1537.020 1542.390 ;
        RECT 1714.020 1542.380 1717.020 1542.390 ;
        RECT 1894.020 1542.380 1897.020 1542.390 ;
        RECT 2074.020 1542.380 2077.020 1542.390 ;
        RECT 2254.020 1542.380 2257.020 1542.390 ;
        RECT 2434.020 1542.380 2437.020 1542.390 ;
        RECT 2614.020 1542.380 2617.020 1542.390 ;
        RECT 2794.020 1542.380 2797.020 1542.390 ;
        RECT 2931.200 1542.380 2934.200 1542.390 ;
        RECT -14.580 1539.380 2934.200 1542.380 ;
        RECT -14.580 1539.370 -11.580 1539.380 ;
        RECT 94.020 1539.370 97.020 1539.380 ;
        RECT 274.020 1539.370 277.020 1539.380 ;
        RECT 454.020 1539.370 457.020 1539.380 ;
        RECT 634.020 1539.370 637.020 1539.380 ;
        RECT 814.020 1539.370 817.020 1539.380 ;
        RECT 994.020 1539.370 997.020 1539.380 ;
        RECT 1174.020 1539.370 1177.020 1539.380 ;
        RECT 1354.020 1539.370 1357.020 1539.380 ;
        RECT 1534.020 1539.370 1537.020 1539.380 ;
        RECT 1714.020 1539.370 1717.020 1539.380 ;
        RECT 1894.020 1539.370 1897.020 1539.380 ;
        RECT 2074.020 1539.370 2077.020 1539.380 ;
        RECT 2254.020 1539.370 2257.020 1539.380 ;
        RECT 2434.020 1539.370 2437.020 1539.380 ;
        RECT 2614.020 1539.370 2617.020 1539.380 ;
        RECT 2794.020 1539.370 2797.020 1539.380 ;
        RECT 2931.200 1539.370 2934.200 1539.380 ;
        RECT -14.580 1362.380 -11.580 1362.390 ;
        RECT 94.020 1362.380 97.020 1362.390 ;
        RECT 274.020 1362.380 277.020 1362.390 ;
        RECT 454.020 1362.380 457.020 1362.390 ;
        RECT 634.020 1362.380 637.020 1362.390 ;
        RECT 814.020 1362.380 817.020 1362.390 ;
        RECT 994.020 1362.380 997.020 1362.390 ;
        RECT 1174.020 1362.380 1177.020 1362.390 ;
        RECT 1354.020 1362.380 1357.020 1362.390 ;
        RECT 1534.020 1362.380 1537.020 1362.390 ;
        RECT 1714.020 1362.380 1717.020 1362.390 ;
        RECT 1894.020 1362.380 1897.020 1362.390 ;
        RECT 2074.020 1362.380 2077.020 1362.390 ;
        RECT 2254.020 1362.380 2257.020 1362.390 ;
        RECT 2434.020 1362.380 2437.020 1362.390 ;
        RECT 2614.020 1362.380 2617.020 1362.390 ;
        RECT 2794.020 1362.380 2797.020 1362.390 ;
        RECT 2931.200 1362.380 2934.200 1362.390 ;
        RECT -14.580 1359.380 2934.200 1362.380 ;
        RECT -14.580 1359.370 -11.580 1359.380 ;
        RECT 94.020 1359.370 97.020 1359.380 ;
        RECT 274.020 1359.370 277.020 1359.380 ;
        RECT 454.020 1359.370 457.020 1359.380 ;
        RECT 634.020 1359.370 637.020 1359.380 ;
        RECT 814.020 1359.370 817.020 1359.380 ;
        RECT 994.020 1359.370 997.020 1359.380 ;
        RECT 1174.020 1359.370 1177.020 1359.380 ;
        RECT 1354.020 1359.370 1357.020 1359.380 ;
        RECT 1534.020 1359.370 1537.020 1359.380 ;
        RECT 1714.020 1359.370 1717.020 1359.380 ;
        RECT 1894.020 1359.370 1897.020 1359.380 ;
        RECT 2074.020 1359.370 2077.020 1359.380 ;
        RECT 2254.020 1359.370 2257.020 1359.380 ;
        RECT 2434.020 1359.370 2437.020 1359.380 ;
        RECT 2614.020 1359.370 2617.020 1359.380 ;
        RECT 2794.020 1359.370 2797.020 1359.380 ;
        RECT 2931.200 1359.370 2934.200 1359.380 ;
        RECT -14.580 1182.380 -11.580 1182.390 ;
        RECT 94.020 1182.380 97.020 1182.390 ;
        RECT 274.020 1182.380 277.020 1182.390 ;
        RECT 454.020 1182.380 457.020 1182.390 ;
        RECT 634.020 1182.380 637.020 1182.390 ;
        RECT 814.020 1182.380 817.020 1182.390 ;
        RECT 994.020 1182.380 997.020 1182.390 ;
        RECT 1174.020 1182.380 1177.020 1182.390 ;
        RECT 1354.020 1182.380 1357.020 1182.390 ;
        RECT 1534.020 1182.380 1537.020 1182.390 ;
        RECT 1714.020 1182.380 1717.020 1182.390 ;
        RECT 1894.020 1182.380 1897.020 1182.390 ;
        RECT 2074.020 1182.380 2077.020 1182.390 ;
        RECT 2254.020 1182.380 2257.020 1182.390 ;
        RECT 2434.020 1182.380 2437.020 1182.390 ;
        RECT 2614.020 1182.380 2617.020 1182.390 ;
        RECT 2794.020 1182.380 2797.020 1182.390 ;
        RECT 2931.200 1182.380 2934.200 1182.390 ;
        RECT -14.580 1179.380 2934.200 1182.380 ;
        RECT -14.580 1179.370 -11.580 1179.380 ;
        RECT 94.020 1179.370 97.020 1179.380 ;
        RECT 274.020 1179.370 277.020 1179.380 ;
        RECT 454.020 1179.370 457.020 1179.380 ;
        RECT 634.020 1179.370 637.020 1179.380 ;
        RECT 814.020 1179.370 817.020 1179.380 ;
        RECT 994.020 1179.370 997.020 1179.380 ;
        RECT 1174.020 1179.370 1177.020 1179.380 ;
        RECT 1354.020 1179.370 1357.020 1179.380 ;
        RECT 1534.020 1179.370 1537.020 1179.380 ;
        RECT 1714.020 1179.370 1717.020 1179.380 ;
        RECT 1894.020 1179.370 1897.020 1179.380 ;
        RECT 2074.020 1179.370 2077.020 1179.380 ;
        RECT 2254.020 1179.370 2257.020 1179.380 ;
        RECT 2434.020 1179.370 2437.020 1179.380 ;
        RECT 2614.020 1179.370 2617.020 1179.380 ;
        RECT 2794.020 1179.370 2797.020 1179.380 ;
        RECT 2931.200 1179.370 2934.200 1179.380 ;
        RECT -14.580 1002.380 -11.580 1002.390 ;
        RECT 94.020 1002.380 97.020 1002.390 ;
        RECT 274.020 1002.380 277.020 1002.390 ;
        RECT 454.020 1002.380 457.020 1002.390 ;
        RECT 634.020 1002.380 637.020 1002.390 ;
        RECT 814.020 1002.380 817.020 1002.390 ;
        RECT 994.020 1002.380 997.020 1002.390 ;
        RECT 1174.020 1002.380 1177.020 1002.390 ;
        RECT 1354.020 1002.380 1357.020 1002.390 ;
        RECT 1534.020 1002.380 1537.020 1002.390 ;
        RECT 1714.020 1002.380 1717.020 1002.390 ;
        RECT 1894.020 1002.380 1897.020 1002.390 ;
        RECT 2074.020 1002.380 2077.020 1002.390 ;
        RECT 2254.020 1002.380 2257.020 1002.390 ;
        RECT 2434.020 1002.380 2437.020 1002.390 ;
        RECT 2614.020 1002.380 2617.020 1002.390 ;
        RECT 2794.020 1002.380 2797.020 1002.390 ;
        RECT 2931.200 1002.380 2934.200 1002.390 ;
        RECT -14.580 999.380 2934.200 1002.380 ;
        RECT -14.580 999.370 -11.580 999.380 ;
        RECT 94.020 999.370 97.020 999.380 ;
        RECT 274.020 999.370 277.020 999.380 ;
        RECT 454.020 999.370 457.020 999.380 ;
        RECT 634.020 999.370 637.020 999.380 ;
        RECT 814.020 999.370 817.020 999.380 ;
        RECT 994.020 999.370 997.020 999.380 ;
        RECT 1174.020 999.370 1177.020 999.380 ;
        RECT 1354.020 999.370 1357.020 999.380 ;
        RECT 1534.020 999.370 1537.020 999.380 ;
        RECT 1714.020 999.370 1717.020 999.380 ;
        RECT 1894.020 999.370 1897.020 999.380 ;
        RECT 2074.020 999.370 2077.020 999.380 ;
        RECT 2254.020 999.370 2257.020 999.380 ;
        RECT 2434.020 999.370 2437.020 999.380 ;
        RECT 2614.020 999.370 2617.020 999.380 ;
        RECT 2794.020 999.370 2797.020 999.380 ;
        RECT 2931.200 999.370 2934.200 999.380 ;
        RECT -14.580 822.380 -11.580 822.390 ;
        RECT 94.020 822.380 97.020 822.390 ;
        RECT 274.020 822.380 277.020 822.390 ;
        RECT 454.020 822.380 457.020 822.390 ;
        RECT 634.020 822.380 637.020 822.390 ;
        RECT 814.020 822.380 817.020 822.390 ;
        RECT 994.020 822.380 997.020 822.390 ;
        RECT 1174.020 822.380 1177.020 822.390 ;
        RECT 1354.020 822.380 1357.020 822.390 ;
        RECT 1534.020 822.380 1537.020 822.390 ;
        RECT 1714.020 822.380 1717.020 822.390 ;
        RECT 1894.020 822.380 1897.020 822.390 ;
        RECT 2074.020 822.380 2077.020 822.390 ;
        RECT 2254.020 822.380 2257.020 822.390 ;
        RECT 2434.020 822.380 2437.020 822.390 ;
        RECT 2614.020 822.380 2617.020 822.390 ;
        RECT 2794.020 822.380 2797.020 822.390 ;
        RECT 2931.200 822.380 2934.200 822.390 ;
        RECT -14.580 819.380 2934.200 822.380 ;
        RECT -14.580 819.370 -11.580 819.380 ;
        RECT 94.020 819.370 97.020 819.380 ;
        RECT 274.020 819.370 277.020 819.380 ;
        RECT 454.020 819.370 457.020 819.380 ;
        RECT 634.020 819.370 637.020 819.380 ;
        RECT 814.020 819.370 817.020 819.380 ;
        RECT 994.020 819.370 997.020 819.380 ;
        RECT 1174.020 819.370 1177.020 819.380 ;
        RECT 1354.020 819.370 1357.020 819.380 ;
        RECT 1534.020 819.370 1537.020 819.380 ;
        RECT 1714.020 819.370 1717.020 819.380 ;
        RECT 1894.020 819.370 1897.020 819.380 ;
        RECT 2074.020 819.370 2077.020 819.380 ;
        RECT 2254.020 819.370 2257.020 819.380 ;
        RECT 2434.020 819.370 2437.020 819.380 ;
        RECT 2614.020 819.370 2617.020 819.380 ;
        RECT 2794.020 819.370 2797.020 819.380 ;
        RECT 2931.200 819.370 2934.200 819.380 ;
        RECT -14.580 642.380 -11.580 642.390 ;
        RECT 94.020 642.380 97.020 642.390 ;
        RECT 274.020 642.380 277.020 642.390 ;
        RECT 454.020 642.380 457.020 642.390 ;
        RECT 634.020 642.380 637.020 642.390 ;
        RECT 814.020 642.380 817.020 642.390 ;
        RECT 994.020 642.380 997.020 642.390 ;
        RECT 1174.020 642.380 1177.020 642.390 ;
        RECT 1354.020 642.380 1357.020 642.390 ;
        RECT 1534.020 642.380 1537.020 642.390 ;
        RECT 1714.020 642.380 1717.020 642.390 ;
        RECT 1894.020 642.380 1897.020 642.390 ;
        RECT 2074.020 642.380 2077.020 642.390 ;
        RECT 2254.020 642.380 2257.020 642.390 ;
        RECT 2434.020 642.380 2437.020 642.390 ;
        RECT 2614.020 642.380 2617.020 642.390 ;
        RECT 2794.020 642.380 2797.020 642.390 ;
        RECT 2931.200 642.380 2934.200 642.390 ;
        RECT -14.580 639.380 2934.200 642.380 ;
        RECT -14.580 639.370 -11.580 639.380 ;
        RECT 94.020 639.370 97.020 639.380 ;
        RECT 274.020 639.370 277.020 639.380 ;
        RECT 454.020 639.370 457.020 639.380 ;
        RECT 634.020 639.370 637.020 639.380 ;
        RECT 814.020 639.370 817.020 639.380 ;
        RECT 994.020 639.370 997.020 639.380 ;
        RECT 1174.020 639.370 1177.020 639.380 ;
        RECT 1354.020 639.370 1357.020 639.380 ;
        RECT 1534.020 639.370 1537.020 639.380 ;
        RECT 1714.020 639.370 1717.020 639.380 ;
        RECT 1894.020 639.370 1897.020 639.380 ;
        RECT 2074.020 639.370 2077.020 639.380 ;
        RECT 2254.020 639.370 2257.020 639.380 ;
        RECT 2434.020 639.370 2437.020 639.380 ;
        RECT 2614.020 639.370 2617.020 639.380 ;
        RECT 2794.020 639.370 2797.020 639.380 ;
        RECT 2931.200 639.370 2934.200 639.380 ;
        RECT -14.580 462.380 -11.580 462.390 ;
        RECT 94.020 462.380 97.020 462.390 ;
        RECT 274.020 462.380 277.020 462.390 ;
        RECT 454.020 462.380 457.020 462.390 ;
        RECT 634.020 462.380 637.020 462.390 ;
        RECT 814.020 462.380 817.020 462.390 ;
        RECT 994.020 462.380 997.020 462.390 ;
        RECT 1174.020 462.380 1177.020 462.390 ;
        RECT 1354.020 462.380 1357.020 462.390 ;
        RECT 1534.020 462.380 1537.020 462.390 ;
        RECT 1714.020 462.380 1717.020 462.390 ;
        RECT 1894.020 462.380 1897.020 462.390 ;
        RECT 2074.020 462.380 2077.020 462.390 ;
        RECT 2254.020 462.380 2257.020 462.390 ;
        RECT 2434.020 462.380 2437.020 462.390 ;
        RECT 2614.020 462.380 2617.020 462.390 ;
        RECT 2794.020 462.380 2797.020 462.390 ;
        RECT 2931.200 462.380 2934.200 462.390 ;
        RECT -14.580 459.380 2934.200 462.380 ;
        RECT -14.580 459.370 -11.580 459.380 ;
        RECT 94.020 459.370 97.020 459.380 ;
        RECT 274.020 459.370 277.020 459.380 ;
        RECT 454.020 459.370 457.020 459.380 ;
        RECT 634.020 459.370 637.020 459.380 ;
        RECT 814.020 459.370 817.020 459.380 ;
        RECT 994.020 459.370 997.020 459.380 ;
        RECT 1174.020 459.370 1177.020 459.380 ;
        RECT 1354.020 459.370 1357.020 459.380 ;
        RECT 1534.020 459.370 1537.020 459.380 ;
        RECT 1714.020 459.370 1717.020 459.380 ;
        RECT 1894.020 459.370 1897.020 459.380 ;
        RECT 2074.020 459.370 2077.020 459.380 ;
        RECT 2254.020 459.370 2257.020 459.380 ;
        RECT 2434.020 459.370 2437.020 459.380 ;
        RECT 2614.020 459.370 2617.020 459.380 ;
        RECT 2794.020 459.370 2797.020 459.380 ;
        RECT 2931.200 459.370 2934.200 459.380 ;
        RECT -14.580 282.380 -11.580 282.390 ;
        RECT 94.020 282.380 97.020 282.390 ;
        RECT 274.020 282.380 277.020 282.390 ;
        RECT 454.020 282.380 457.020 282.390 ;
        RECT 634.020 282.380 637.020 282.390 ;
        RECT 814.020 282.380 817.020 282.390 ;
        RECT 994.020 282.380 997.020 282.390 ;
        RECT 1174.020 282.380 1177.020 282.390 ;
        RECT 1354.020 282.380 1357.020 282.390 ;
        RECT 1534.020 282.380 1537.020 282.390 ;
        RECT 1714.020 282.380 1717.020 282.390 ;
        RECT 1894.020 282.380 1897.020 282.390 ;
        RECT 2074.020 282.380 2077.020 282.390 ;
        RECT 2254.020 282.380 2257.020 282.390 ;
        RECT 2434.020 282.380 2437.020 282.390 ;
        RECT 2614.020 282.380 2617.020 282.390 ;
        RECT 2794.020 282.380 2797.020 282.390 ;
        RECT 2931.200 282.380 2934.200 282.390 ;
        RECT -14.580 279.380 2934.200 282.380 ;
        RECT -14.580 279.370 -11.580 279.380 ;
        RECT 94.020 279.370 97.020 279.380 ;
        RECT 274.020 279.370 277.020 279.380 ;
        RECT 454.020 279.370 457.020 279.380 ;
        RECT 634.020 279.370 637.020 279.380 ;
        RECT 814.020 279.370 817.020 279.380 ;
        RECT 994.020 279.370 997.020 279.380 ;
        RECT 1174.020 279.370 1177.020 279.380 ;
        RECT 1354.020 279.370 1357.020 279.380 ;
        RECT 1534.020 279.370 1537.020 279.380 ;
        RECT 1714.020 279.370 1717.020 279.380 ;
        RECT 1894.020 279.370 1897.020 279.380 ;
        RECT 2074.020 279.370 2077.020 279.380 ;
        RECT 2254.020 279.370 2257.020 279.380 ;
        RECT 2434.020 279.370 2437.020 279.380 ;
        RECT 2614.020 279.370 2617.020 279.380 ;
        RECT 2794.020 279.370 2797.020 279.380 ;
        RECT 2931.200 279.370 2934.200 279.380 ;
        RECT -14.580 102.380 -11.580 102.390 ;
        RECT 94.020 102.380 97.020 102.390 ;
        RECT 274.020 102.380 277.020 102.390 ;
        RECT 454.020 102.380 457.020 102.390 ;
        RECT 634.020 102.380 637.020 102.390 ;
        RECT 814.020 102.380 817.020 102.390 ;
        RECT 994.020 102.380 997.020 102.390 ;
        RECT 1174.020 102.380 1177.020 102.390 ;
        RECT 1354.020 102.380 1357.020 102.390 ;
        RECT 1534.020 102.380 1537.020 102.390 ;
        RECT 1714.020 102.380 1717.020 102.390 ;
        RECT 1894.020 102.380 1897.020 102.390 ;
        RECT 2074.020 102.380 2077.020 102.390 ;
        RECT 2254.020 102.380 2257.020 102.390 ;
        RECT 2434.020 102.380 2437.020 102.390 ;
        RECT 2614.020 102.380 2617.020 102.390 ;
        RECT 2794.020 102.380 2797.020 102.390 ;
        RECT 2931.200 102.380 2934.200 102.390 ;
        RECT -14.580 99.380 2934.200 102.380 ;
        RECT -14.580 99.370 -11.580 99.380 ;
        RECT 94.020 99.370 97.020 99.380 ;
        RECT 274.020 99.370 277.020 99.380 ;
        RECT 454.020 99.370 457.020 99.380 ;
        RECT 634.020 99.370 637.020 99.380 ;
        RECT 814.020 99.370 817.020 99.380 ;
        RECT 994.020 99.370 997.020 99.380 ;
        RECT 1174.020 99.370 1177.020 99.380 ;
        RECT 1354.020 99.370 1357.020 99.380 ;
        RECT 1534.020 99.370 1537.020 99.380 ;
        RECT 1714.020 99.370 1717.020 99.380 ;
        RECT 1894.020 99.370 1897.020 99.380 ;
        RECT 2074.020 99.370 2077.020 99.380 ;
        RECT 2254.020 99.370 2257.020 99.380 ;
        RECT 2434.020 99.370 2437.020 99.380 ;
        RECT 2614.020 99.370 2617.020 99.380 ;
        RECT 2794.020 99.370 2797.020 99.380 ;
        RECT 2931.200 99.370 2934.200 99.380 ;
        RECT -14.580 -6.220 -11.580 -6.210 ;
        RECT 94.020 -6.220 97.020 -6.210 ;
        RECT 274.020 -6.220 277.020 -6.210 ;
        RECT 454.020 -6.220 457.020 -6.210 ;
        RECT 634.020 -6.220 637.020 -6.210 ;
        RECT 814.020 -6.220 817.020 -6.210 ;
        RECT 994.020 -6.220 997.020 -6.210 ;
        RECT 1174.020 -6.220 1177.020 -6.210 ;
        RECT 1354.020 -6.220 1357.020 -6.210 ;
        RECT 1534.020 -6.220 1537.020 -6.210 ;
        RECT 1714.020 -6.220 1717.020 -6.210 ;
        RECT 1894.020 -6.220 1897.020 -6.210 ;
        RECT 2074.020 -6.220 2077.020 -6.210 ;
        RECT 2254.020 -6.220 2257.020 -6.210 ;
        RECT 2434.020 -6.220 2437.020 -6.210 ;
        RECT 2614.020 -6.220 2617.020 -6.210 ;
        RECT 2794.020 -6.220 2797.020 -6.210 ;
        RECT 2931.200 -6.220 2934.200 -6.210 ;
        RECT -14.580 -9.220 2934.200 -6.220 ;
        RECT -14.580 -9.230 -11.580 -9.220 ;
        RECT 94.020 -9.230 97.020 -9.220 ;
        RECT 274.020 -9.230 277.020 -9.220 ;
        RECT 454.020 -9.230 457.020 -9.220 ;
        RECT 634.020 -9.230 637.020 -9.220 ;
        RECT 814.020 -9.230 817.020 -9.220 ;
        RECT 994.020 -9.230 997.020 -9.220 ;
        RECT 1174.020 -9.230 1177.020 -9.220 ;
        RECT 1354.020 -9.230 1357.020 -9.220 ;
        RECT 1534.020 -9.230 1537.020 -9.220 ;
        RECT 1714.020 -9.230 1717.020 -9.220 ;
        RECT 1894.020 -9.230 1897.020 -9.220 ;
        RECT 2074.020 -9.230 2077.020 -9.220 ;
        RECT 2254.020 -9.230 2257.020 -9.220 ;
        RECT 2434.020 -9.230 2437.020 -9.220 ;
        RECT 2614.020 -9.230 2617.020 -9.220 ;
        RECT 2794.020 -9.230 2797.020 -9.220 ;
        RECT 2931.200 -9.230 2934.200 -9.220 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -19.180 -13.820 -16.180 3533.500 ;
        RECT 22.020 -18.420 25.020 3538.100 ;
        RECT 202.020 -18.420 205.020 3538.100 ;
        RECT 382.020 -18.420 385.020 3538.100 ;
        RECT 562.020 -18.420 565.020 3538.100 ;
        RECT 742.020 -18.420 745.020 3538.100 ;
        RECT 922.020 -18.420 925.020 3538.100 ;
        RECT 1102.020 -18.420 1105.020 3538.100 ;
        RECT 1282.020 -18.420 1285.020 3538.100 ;
        RECT 1462.020 -18.420 1465.020 3538.100 ;
        RECT 1642.020 -18.420 1645.020 3538.100 ;
        RECT 1822.020 -18.420 1825.020 3538.100 ;
        RECT 2002.020 -18.420 2005.020 3538.100 ;
        RECT 2182.020 -18.420 2185.020 3538.100 ;
        RECT 2362.020 -18.420 2365.020 3538.100 ;
        RECT 2542.020 -18.420 2545.020 3538.100 ;
        RECT 2722.020 -18.420 2725.020 3538.100 ;
        RECT 2902.020 -18.420 2905.020 3538.100 ;
        RECT 2935.800 -13.820 2938.800 3533.500 ;
      LAYER via4 ;
        RECT -18.270 3532.210 -17.090 3533.390 ;
        RECT -18.270 3530.610 -17.090 3531.790 ;
        RECT -18.270 3449.090 -17.090 3450.270 ;
        RECT -18.270 3447.490 -17.090 3448.670 ;
        RECT -18.270 3269.090 -17.090 3270.270 ;
        RECT -18.270 3267.490 -17.090 3268.670 ;
        RECT -18.270 3089.090 -17.090 3090.270 ;
        RECT -18.270 3087.490 -17.090 3088.670 ;
        RECT -18.270 2909.090 -17.090 2910.270 ;
        RECT -18.270 2907.490 -17.090 2908.670 ;
        RECT -18.270 2729.090 -17.090 2730.270 ;
        RECT -18.270 2727.490 -17.090 2728.670 ;
        RECT -18.270 2549.090 -17.090 2550.270 ;
        RECT -18.270 2547.490 -17.090 2548.670 ;
        RECT -18.270 2369.090 -17.090 2370.270 ;
        RECT -18.270 2367.490 -17.090 2368.670 ;
        RECT -18.270 2189.090 -17.090 2190.270 ;
        RECT -18.270 2187.490 -17.090 2188.670 ;
        RECT -18.270 2009.090 -17.090 2010.270 ;
        RECT -18.270 2007.490 -17.090 2008.670 ;
        RECT -18.270 1829.090 -17.090 1830.270 ;
        RECT -18.270 1827.490 -17.090 1828.670 ;
        RECT -18.270 1649.090 -17.090 1650.270 ;
        RECT -18.270 1647.490 -17.090 1648.670 ;
        RECT -18.270 1469.090 -17.090 1470.270 ;
        RECT -18.270 1467.490 -17.090 1468.670 ;
        RECT -18.270 1289.090 -17.090 1290.270 ;
        RECT -18.270 1287.490 -17.090 1288.670 ;
        RECT -18.270 1109.090 -17.090 1110.270 ;
        RECT -18.270 1107.490 -17.090 1108.670 ;
        RECT -18.270 929.090 -17.090 930.270 ;
        RECT -18.270 927.490 -17.090 928.670 ;
        RECT -18.270 749.090 -17.090 750.270 ;
        RECT -18.270 747.490 -17.090 748.670 ;
        RECT -18.270 569.090 -17.090 570.270 ;
        RECT -18.270 567.490 -17.090 568.670 ;
        RECT -18.270 389.090 -17.090 390.270 ;
        RECT -18.270 387.490 -17.090 388.670 ;
        RECT -18.270 209.090 -17.090 210.270 ;
        RECT -18.270 207.490 -17.090 208.670 ;
        RECT -18.270 29.090 -17.090 30.270 ;
        RECT -18.270 27.490 -17.090 28.670 ;
        RECT -18.270 -12.110 -17.090 -10.930 ;
        RECT -18.270 -13.710 -17.090 -12.530 ;
        RECT 22.930 3532.210 24.110 3533.390 ;
        RECT 22.930 3530.610 24.110 3531.790 ;
        RECT 22.930 3449.090 24.110 3450.270 ;
        RECT 22.930 3447.490 24.110 3448.670 ;
        RECT 22.930 3269.090 24.110 3270.270 ;
        RECT 22.930 3267.490 24.110 3268.670 ;
        RECT 22.930 3089.090 24.110 3090.270 ;
        RECT 22.930 3087.490 24.110 3088.670 ;
        RECT 22.930 2909.090 24.110 2910.270 ;
        RECT 22.930 2907.490 24.110 2908.670 ;
        RECT 22.930 2729.090 24.110 2730.270 ;
        RECT 22.930 2727.490 24.110 2728.670 ;
        RECT 22.930 2549.090 24.110 2550.270 ;
        RECT 22.930 2547.490 24.110 2548.670 ;
        RECT 22.930 2369.090 24.110 2370.270 ;
        RECT 22.930 2367.490 24.110 2368.670 ;
        RECT 22.930 2189.090 24.110 2190.270 ;
        RECT 22.930 2187.490 24.110 2188.670 ;
        RECT 22.930 2009.090 24.110 2010.270 ;
        RECT 22.930 2007.490 24.110 2008.670 ;
        RECT 22.930 1829.090 24.110 1830.270 ;
        RECT 22.930 1827.490 24.110 1828.670 ;
        RECT 22.930 1649.090 24.110 1650.270 ;
        RECT 22.930 1647.490 24.110 1648.670 ;
        RECT 22.930 1469.090 24.110 1470.270 ;
        RECT 22.930 1467.490 24.110 1468.670 ;
        RECT 22.930 1289.090 24.110 1290.270 ;
        RECT 22.930 1287.490 24.110 1288.670 ;
        RECT 22.930 1109.090 24.110 1110.270 ;
        RECT 22.930 1107.490 24.110 1108.670 ;
        RECT 22.930 929.090 24.110 930.270 ;
        RECT 22.930 927.490 24.110 928.670 ;
        RECT 22.930 749.090 24.110 750.270 ;
        RECT 22.930 747.490 24.110 748.670 ;
        RECT 22.930 569.090 24.110 570.270 ;
        RECT 22.930 567.490 24.110 568.670 ;
        RECT 22.930 389.090 24.110 390.270 ;
        RECT 22.930 387.490 24.110 388.670 ;
        RECT 22.930 209.090 24.110 210.270 ;
        RECT 22.930 207.490 24.110 208.670 ;
        RECT 22.930 29.090 24.110 30.270 ;
        RECT 22.930 27.490 24.110 28.670 ;
        RECT 22.930 -12.110 24.110 -10.930 ;
        RECT 22.930 -13.710 24.110 -12.530 ;
        RECT 202.930 3532.210 204.110 3533.390 ;
        RECT 202.930 3530.610 204.110 3531.790 ;
        RECT 202.930 3449.090 204.110 3450.270 ;
        RECT 202.930 3447.490 204.110 3448.670 ;
        RECT 202.930 3269.090 204.110 3270.270 ;
        RECT 202.930 3267.490 204.110 3268.670 ;
        RECT 202.930 3089.090 204.110 3090.270 ;
        RECT 202.930 3087.490 204.110 3088.670 ;
        RECT 202.930 2909.090 204.110 2910.270 ;
        RECT 202.930 2907.490 204.110 2908.670 ;
        RECT 202.930 2729.090 204.110 2730.270 ;
        RECT 202.930 2727.490 204.110 2728.670 ;
        RECT 202.930 2549.090 204.110 2550.270 ;
        RECT 202.930 2547.490 204.110 2548.670 ;
        RECT 202.930 2369.090 204.110 2370.270 ;
        RECT 202.930 2367.490 204.110 2368.670 ;
        RECT 202.930 2189.090 204.110 2190.270 ;
        RECT 202.930 2187.490 204.110 2188.670 ;
        RECT 202.930 2009.090 204.110 2010.270 ;
        RECT 202.930 2007.490 204.110 2008.670 ;
        RECT 202.930 1829.090 204.110 1830.270 ;
        RECT 202.930 1827.490 204.110 1828.670 ;
        RECT 202.930 1649.090 204.110 1650.270 ;
        RECT 202.930 1647.490 204.110 1648.670 ;
        RECT 202.930 1469.090 204.110 1470.270 ;
        RECT 202.930 1467.490 204.110 1468.670 ;
        RECT 202.930 1289.090 204.110 1290.270 ;
        RECT 202.930 1287.490 204.110 1288.670 ;
        RECT 202.930 1109.090 204.110 1110.270 ;
        RECT 202.930 1107.490 204.110 1108.670 ;
        RECT 202.930 929.090 204.110 930.270 ;
        RECT 202.930 927.490 204.110 928.670 ;
        RECT 202.930 749.090 204.110 750.270 ;
        RECT 202.930 747.490 204.110 748.670 ;
        RECT 202.930 569.090 204.110 570.270 ;
        RECT 202.930 567.490 204.110 568.670 ;
        RECT 202.930 389.090 204.110 390.270 ;
        RECT 202.930 387.490 204.110 388.670 ;
        RECT 202.930 209.090 204.110 210.270 ;
        RECT 202.930 207.490 204.110 208.670 ;
        RECT 202.930 29.090 204.110 30.270 ;
        RECT 202.930 27.490 204.110 28.670 ;
        RECT 202.930 -12.110 204.110 -10.930 ;
        RECT 202.930 -13.710 204.110 -12.530 ;
        RECT 382.930 3532.210 384.110 3533.390 ;
        RECT 382.930 3530.610 384.110 3531.790 ;
        RECT 382.930 3449.090 384.110 3450.270 ;
        RECT 382.930 3447.490 384.110 3448.670 ;
        RECT 382.930 3269.090 384.110 3270.270 ;
        RECT 382.930 3267.490 384.110 3268.670 ;
        RECT 382.930 3089.090 384.110 3090.270 ;
        RECT 382.930 3087.490 384.110 3088.670 ;
        RECT 382.930 2909.090 384.110 2910.270 ;
        RECT 382.930 2907.490 384.110 2908.670 ;
        RECT 382.930 2729.090 384.110 2730.270 ;
        RECT 382.930 2727.490 384.110 2728.670 ;
        RECT 382.930 2549.090 384.110 2550.270 ;
        RECT 382.930 2547.490 384.110 2548.670 ;
        RECT 382.930 2369.090 384.110 2370.270 ;
        RECT 382.930 2367.490 384.110 2368.670 ;
        RECT 382.930 2189.090 384.110 2190.270 ;
        RECT 382.930 2187.490 384.110 2188.670 ;
        RECT 382.930 2009.090 384.110 2010.270 ;
        RECT 382.930 2007.490 384.110 2008.670 ;
        RECT 382.930 1829.090 384.110 1830.270 ;
        RECT 382.930 1827.490 384.110 1828.670 ;
        RECT 382.930 1649.090 384.110 1650.270 ;
        RECT 382.930 1647.490 384.110 1648.670 ;
        RECT 382.930 1469.090 384.110 1470.270 ;
        RECT 382.930 1467.490 384.110 1468.670 ;
        RECT 382.930 1289.090 384.110 1290.270 ;
        RECT 382.930 1287.490 384.110 1288.670 ;
        RECT 382.930 1109.090 384.110 1110.270 ;
        RECT 382.930 1107.490 384.110 1108.670 ;
        RECT 382.930 929.090 384.110 930.270 ;
        RECT 382.930 927.490 384.110 928.670 ;
        RECT 382.930 749.090 384.110 750.270 ;
        RECT 382.930 747.490 384.110 748.670 ;
        RECT 382.930 569.090 384.110 570.270 ;
        RECT 382.930 567.490 384.110 568.670 ;
        RECT 382.930 389.090 384.110 390.270 ;
        RECT 382.930 387.490 384.110 388.670 ;
        RECT 382.930 209.090 384.110 210.270 ;
        RECT 382.930 207.490 384.110 208.670 ;
        RECT 382.930 29.090 384.110 30.270 ;
        RECT 382.930 27.490 384.110 28.670 ;
        RECT 382.930 -12.110 384.110 -10.930 ;
        RECT 382.930 -13.710 384.110 -12.530 ;
        RECT 562.930 3532.210 564.110 3533.390 ;
        RECT 562.930 3530.610 564.110 3531.790 ;
        RECT 562.930 3449.090 564.110 3450.270 ;
        RECT 562.930 3447.490 564.110 3448.670 ;
        RECT 562.930 3269.090 564.110 3270.270 ;
        RECT 562.930 3267.490 564.110 3268.670 ;
        RECT 562.930 3089.090 564.110 3090.270 ;
        RECT 562.930 3087.490 564.110 3088.670 ;
        RECT 562.930 2909.090 564.110 2910.270 ;
        RECT 562.930 2907.490 564.110 2908.670 ;
        RECT 562.930 2729.090 564.110 2730.270 ;
        RECT 562.930 2727.490 564.110 2728.670 ;
        RECT 562.930 2549.090 564.110 2550.270 ;
        RECT 562.930 2547.490 564.110 2548.670 ;
        RECT 562.930 2369.090 564.110 2370.270 ;
        RECT 562.930 2367.490 564.110 2368.670 ;
        RECT 562.930 2189.090 564.110 2190.270 ;
        RECT 562.930 2187.490 564.110 2188.670 ;
        RECT 562.930 2009.090 564.110 2010.270 ;
        RECT 562.930 2007.490 564.110 2008.670 ;
        RECT 562.930 1829.090 564.110 1830.270 ;
        RECT 562.930 1827.490 564.110 1828.670 ;
        RECT 562.930 1649.090 564.110 1650.270 ;
        RECT 562.930 1647.490 564.110 1648.670 ;
        RECT 562.930 1469.090 564.110 1470.270 ;
        RECT 562.930 1467.490 564.110 1468.670 ;
        RECT 562.930 1289.090 564.110 1290.270 ;
        RECT 562.930 1287.490 564.110 1288.670 ;
        RECT 562.930 1109.090 564.110 1110.270 ;
        RECT 562.930 1107.490 564.110 1108.670 ;
        RECT 562.930 929.090 564.110 930.270 ;
        RECT 562.930 927.490 564.110 928.670 ;
        RECT 562.930 749.090 564.110 750.270 ;
        RECT 562.930 747.490 564.110 748.670 ;
        RECT 562.930 569.090 564.110 570.270 ;
        RECT 562.930 567.490 564.110 568.670 ;
        RECT 562.930 389.090 564.110 390.270 ;
        RECT 562.930 387.490 564.110 388.670 ;
        RECT 562.930 209.090 564.110 210.270 ;
        RECT 562.930 207.490 564.110 208.670 ;
        RECT 562.930 29.090 564.110 30.270 ;
        RECT 562.930 27.490 564.110 28.670 ;
        RECT 562.930 -12.110 564.110 -10.930 ;
        RECT 562.930 -13.710 564.110 -12.530 ;
        RECT 742.930 3532.210 744.110 3533.390 ;
        RECT 742.930 3530.610 744.110 3531.790 ;
        RECT 742.930 3449.090 744.110 3450.270 ;
        RECT 742.930 3447.490 744.110 3448.670 ;
        RECT 742.930 3269.090 744.110 3270.270 ;
        RECT 742.930 3267.490 744.110 3268.670 ;
        RECT 742.930 3089.090 744.110 3090.270 ;
        RECT 742.930 3087.490 744.110 3088.670 ;
        RECT 742.930 2909.090 744.110 2910.270 ;
        RECT 742.930 2907.490 744.110 2908.670 ;
        RECT 742.930 2729.090 744.110 2730.270 ;
        RECT 742.930 2727.490 744.110 2728.670 ;
        RECT 742.930 2549.090 744.110 2550.270 ;
        RECT 742.930 2547.490 744.110 2548.670 ;
        RECT 742.930 2369.090 744.110 2370.270 ;
        RECT 742.930 2367.490 744.110 2368.670 ;
        RECT 742.930 2189.090 744.110 2190.270 ;
        RECT 742.930 2187.490 744.110 2188.670 ;
        RECT 742.930 2009.090 744.110 2010.270 ;
        RECT 742.930 2007.490 744.110 2008.670 ;
        RECT 742.930 1829.090 744.110 1830.270 ;
        RECT 742.930 1827.490 744.110 1828.670 ;
        RECT 742.930 1649.090 744.110 1650.270 ;
        RECT 742.930 1647.490 744.110 1648.670 ;
        RECT 742.930 1469.090 744.110 1470.270 ;
        RECT 742.930 1467.490 744.110 1468.670 ;
        RECT 742.930 1289.090 744.110 1290.270 ;
        RECT 742.930 1287.490 744.110 1288.670 ;
        RECT 742.930 1109.090 744.110 1110.270 ;
        RECT 742.930 1107.490 744.110 1108.670 ;
        RECT 742.930 929.090 744.110 930.270 ;
        RECT 742.930 927.490 744.110 928.670 ;
        RECT 742.930 749.090 744.110 750.270 ;
        RECT 742.930 747.490 744.110 748.670 ;
        RECT 742.930 569.090 744.110 570.270 ;
        RECT 742.930 567.490 744.110 568.670 ;
        RECT 742.930 389.090 744.110 390.270 ;
        RECT 742.930 387.490 744.110 388.670 ;
        RECT 742.930 209.090 744.110 210.270 ;
        RECT 742.930 207.490 744.110 208.670 ;
        RECT 742.930 29.090 744.110 30.270 ;
        RECT 742.930 27.490 744.110 28.670 ;
        RECT 742.930 -12.110 744.110 -10.930 ;
        RECT 742.930 -13.710 744.110 -12.530 ;
        RECT 922.930 3532.210 924.110 3533.390 ;
        RECT 922.930 3530.610 924.110 3531.790 ;
        RECT 922.930 3449.090 924.110 3450.270 ;
        RECT 922.930 3447.490 924.110 3448.670 ;
        RECT 922.930 3269.090 924.110 3270.270 ;
        RECT 922.930 3267.490 924.110 3268.670 ;
        RECT 922.930 3089.090 924.110 3090.270 ;
        RECT 922.930 3087.490 924.110 3088.670 ;
        RECT 922.930 2909.090 924.110 2910.270 ;
        RECT 922.930 2907.490 924.110 2908.670 ;
        RECT 922.930 2729.090 924.110 2730.270 ;
        RECT 922.930 2727.490 924.110 2728.670 ;
        RECT 922.930 2549.090 924.110 2550.270 ;
        RECT 922.930 2547.490 924.110 2548.670 ;
        RECT 922.930 2369.090 924.110 2370.270 ;
        RECT 922.930 2367.490 924.110 2368.670 ;
        RECT 922.930 2189.090 924.110 2190.270 ;
        RECT 922.930 2187.490 924.110 2188.670 ;
        RECT 922.930 2009.090 924.110 2010.270 ;
        RECT 922.930 2007.490 924.110 2008.670 ;
        RECT 922.930 1829.090 924.110 1830.270 ;
        RECT 922.930 1827.490 924.110 1828.670 ;
        RECT 922.930 1649.090 924.110 1650.270 ;
        RECT 922.930 1647.490 924.110 1648.670 ;
        RECT 922.930 1469.090 924.110 1470.270 ;
        RECT 922.930 1467.490 924.110 1468.670 ;
        RECT 922.930 1289.090 924.110 1290.270 ;
        RECT 922.930 1287.490 924.110 1288.670 ;
        RECT 922.930 1109.090 924.110 1110.270 ;
        RECT 922.930 1107.490 924.110 1108.670 ;
        RECT 922.930 929.090 924.110 930.270 ;
        RECT 922.930 927.490 924.110 928.670 ;
        RECT 922.930 749.090 924.110 750.270 ;
        RECT 922.930 747.490 924.110 748.670 ;
        RECT 922.930 569.090 924.110 570.270 ;
        RECT 922.930 567.490 924.110 568.670 ;
        RECT 922.930 389.090 924.110 390.270 ;
        RECT 922.930 387.490 924.110 388.670 ;
        RECT 922.930 209.090 924.110 210.270 ;
        RECT 922.930 207.490 924.110 208.670 ;
        RECT 922.930 29.090 924.110 30.270 ;
        RECT 922.930 27.490 924.110 28.670 ;
        RECT 922.930 -12.110 924.110 -10.930 ;
        RECT 922.930 -13.710 924.110 -12.530 ;
        RECT 1102.930 3532.210 1104.110 3533.390 ;
        RECT 1102.930 3530.610 1104.110 3531.790 ;
        RECT 1102.930 3449.090 1104.110 3450.270 ;
        RECT 1102.930 3447.490 1104.110 3448.670 ;
        RECT 1102.930 3269.090 1104.110 3270.270 ;
        RECT 1102.930 3267.490 1104.110 3268.670 ;
        RECT 1102.930 3089.090 1104.110 3090.270 ;
        RECT 1102.930 3087.490 1104.110 3088.670 ;
        RECT 1102.930 2909.090 1104.110 2910.270 ;
        RECT 1102.930 2907.490 1104.110 2908.670 ;
        RECT 1102.930 2729.090 1104.110 2730.270 ;
        RECT 1102.930 2727.490 1104.110 2728.670 ;
        RECT 1102.930 2549.090 1104.110 2550.270 ;
        RECT 1102.930 2547.490 1104.110 2548.670 ;
        RECT 1102.930 2369.090 1104.110 2370.270 ;
        RECT 1102.930 2367.490 1104.110 2368.670 ;
        RECT 1102.930 2189.090 1104.110 2190.270 ;
        RECT 1102.930 2187.490 1104.110 2188.670 ;
        RECT 1102.930 2009.090 1104.110 2010.270 ;
        RECT 1102.930 2007.490 1104.110 2008.670 ;
        RECT 1102.930 1829.090 1104.110 1830.270 ;
        RECT 1102.930 1827.490 1104.110 1828.670 ;
        RECT 1102.930 1649.090 1104.110 1650.270 ;
        RECT 1102.930 1647.490 1104.110 1648.670 ;
        RECT 1102.930 1469.090 1104.110 1470.270 ;
        RECT 1102.930 1467.490 1104.110 1468.670 ;
        RECT 1102.930 1289.090 1104.110 1290.270 ;
        RECT 1102.930 1287.490 1104.110 1288.670 ;
        RECT 1102.930 1109.090 1104.110 1110.270 ;
        RECT 1102.930 1107.490 1104.110 1108.670 ;
        RECT 1102.930 929.090 1104.110 930.270 ;
        RECT 1102.930 927.490 1104.110 928.670 ;
        RECT 1102.930 749.090 1104.110 750.270 ;
        RECT 1102.930 747.490 1104.110 748.670 ;
        RECT 1102.930 569.090 1104.110 570.270 ;
        RECT 1102.930 567.490 1104.110 568.670 ;
        RECT 1102.930 389.090 1104.110 390.270 ;
        RECT 1102.930 387.490 1104.110 388.670 ;
        RECT 1102.930 209.090 1104.110 210.270 ;
        RECT 1102.930 207.490 1104.110 208.670 ;
        RECT 1102.930 29.090 1104.110 30.270 ;
        RECT 1102.930 27.490 1104.110 28.670 ;
        RECT 1102.930 -12.110 1104.110 -10.930 ;
        RECT 1102.930 -13.710 1104.110 -12.530 ;
        RECT 1282.930 3532.210 1284.110 3533.390 ;
        RECT 1282.930 3530.610 1284.110 3531.790 ;
        RECT 1282.930 3449.090 1284.110 3450.270 ;
        RECT 1282.930 3447.490 1284.110 3448.670 ;
        RECT 1282.930 3269.090 1284.110 3270.270 ;
        RECT 1282.930 3267.490 1284.110 3268.670 ;
        RECT 1282.930 3089.090 1284.110 3090.270 ;
        RECT 1282.930 3087.490 1284.110 3088.670 ;
        RECT 1282.930 2909.090 1284.110 2910.270 ;
        RECT 1282.930 2907.490 1284.110 2908.670 ;
        RECT 1282.930 2729.090 1284.110 2730.270 ;
        RECT 1282.930 2727.490 1284.110 2728.670 ;
        RECT 1282.930 2549.090 1284.110 2550.270 ;
        RECT 1282.930 2547.490 1284.110 2548.670 ;
        RECT 1282.930 2369.090 1284.110 2370.270 ;
        RECT 1282.930 2367.490 1284.110 2368.670 ;
        RECT 1282.930 2189.090 1284.110 2190.270 ;
        RECT 1282.930 2187.490 1284.110 2188.670 ;
        RECT 1282.930 2009.090 1284.110 2010.270 ;
        RECT 1282.930 2007.490 1284.110 2008.670 ;
        RECT 1282.930 1829.090 1284.110 1830.270 ;
        RECT 1282.930 1827.490 1284.110 1828.670 ;
        RECT 1282.930 1649.090 1284.110 1650.270 ;
        RECT 1282.930 1647.490 1284.110 1648.670 ;
        RECT 1282.930 1469.090 1284.110 1470.270 ;
        RECT 1282.930 1467.490 1284.110 1468.670 ;
        RECT 1282.930 1289.090 1284.110 1290.270 ;
        RECT 1282.930 1287.490 1284.110 1288.670 ;
        RECT 1282.930 1109.090 1284.110 1110.270 ;
        RECT 1282.930 1107.490 1284.110 1108.670 ;
        RECT 1282.930 929.090 1284.110 930.270 ;
        RECT 1282.930 927.490 1284.110 928.670 ;
        RECT 1282.930 749.090 1284.110 750.270 ;
        RECT 1282.930 747.490 1284.110 748.670 ;
        RECT 1282.930 569.090 1284.110 570.270 ;
        RECT 1282.930 567.490 1284.110 568.670 ;
        RECT 1282.930 389.090 1284.110 390.270 ;
        RECT 1282.930 387.490 1284.110 388.670 ;
        RECT 1282.930 209.090 1284.110 210.270 ;
        RECT 1282.930 207.490 1284.110 208.670 ;
        RECT 1282.930 29.090 1284.110 30.270 ;
        RECT 1282.930 27.490 1284.110 28.670 ;
        RECT 1282.930 -12.110 1284.110 -10.930 ;
        RECT 1282.930 -13.710 1284.110 -12.530 ;
        RECT 1462.930 3532.210 1464.110 3533.390 ;
        RECT 1462.930 3530.610 1464.110 3531.790 ;
        RECT 1462.930 3449.090 1464.110 3450.270 ;
        RECT 1462.930 3447.490 1464.110 3448.670 ;
        RECT 1462.930 3269.090 1464.110 3270.270 ;
        RECT 1462.930 3267.490 1464.110 3268.670 ;
        RECT 1462.930 3089.090 1464.110 3090.270 ;
        RECT 1462.930 3087.490 1464.110 3088.670 ;
        RECT 1462.930 2909.090 1464.110 2910.270 ;
        RECT 1462.930 2907.490 1464.110 2908.670 ;
        RECT 1462.930 2729.090 1464.110 2730.270 ;
        RECT 1462.930 2727.490 1464.110 2728.670 ;
        RECT 1462.930 2549.090 1464.110 2550.270 ;
        RECT 1462.930 2547.490 1464.110 2548.670 ;
        RECT 1462.930 2369.090 1464.110 2370.270 ;
        RECT 1462.930 2367.490 1464.110 2368.670 ;
        RECT 1462.930 2189.090 1464.110 2190.270 ;
        RECT 1462.930 2187.490 1464.110 2188.670 ;
        RECT 1462.930 2009.090 1464.110 2010.270 ;
        RECT 1462.930 2007.490 1464.110 2008.670 ;
        RECT 1462.930 1829.090 1464.110 1830.270 ;
        RECT 1462.930 1827.490 1464.110 1828.670 ;
        RECT 1462.930 1649.090 1464.110 1650.270 ;
        RECT 1462.930 1647.490 1464.110 1648.670 ;
        RECT 1462.930 1469.090 1464.110 1470.270 ;
        RECT 1462.930 1467.490 1464.110 1468.670 ;
        RECT 1462.930 1289.090 1464.110 1290.270 ;
        RECT 1462.930 1287.490 1464.110 1288.670 ;
        RECT 1462.930 1109.090 1464.110 1110.270 ;
        RECT 1462.930 1107.490 1464.110 1108.670 ;
        RECT 1462.930 929.090 1464.110 930.270 ;
        RECT 1462.930 927.490 1464.110 928.670 ;
        RECT 1462.930 749.090 1464.110 750.270 ;
        RECT 1462.930 747.490 1464.110 748.670 ;
        RECT 1462.930 569.090 1464.110 570.270 ;
        RECT 1462.930 567.490 1464.110 568.670 ;
        RECT 1462.930 389.090 1464.110 390.270 ;
        RECT 1462.930 387.490 1464.110 388.670 ;
        RECT 1462.930 209.090 1464.110 210.270 ;
        RECT 1462.930 207.490 1464.110 208.670 ;
        RECT 1462.930 29.090 1464.110 30.270 ;
        RECT 1462.930 27.490 1464.110 28.670 ;
        RECT 1462.930 -12.110 1464.110 -10.930 ;
        RECT 1462.930 -13.710 1464.110 -12.530 ;
        RECT 1642.930 3532.210 1644.110 3533.390 ;
        RECT 1642.930 3530.610 1644.110 3531.790 ;
        RECT 1642.930 3449.090 1644.110 3450.270 ;
        RECT 1642.930 3447.490 1644.110 3448.670 ;
        RECT 1642.930 3269.090 1644.110 3270.270 ;
        RECT 1642.930 3267.490 1644.110 3268.670 ;
        RECT 1642.930 3089.090 1644.110 3090.270 ;
        RECT 1642.930 3087.490 1644.110 3088.670 ;
        RECT 1642.930 2909.090 1644.110 2910.270 ;
        RECT 1642.930 2907.490 1644.110 2908.670 ;
        RECT 1642.930 2729.090 1644.110 2730.270 ;
        RECT 1642.930 2727.490 1644.110 2728.670 ;
        RECT 1642.930 2549.090 1644.110 2550.270 ;
        RECT 1642.930 2547.490 1644.110 2548.670 ;
        RECT 1642.930 2369.090 1644.110 2370.270 ;
        RECT 1642.930 2367.490 1644.110 2368.670 ;
        RECT 1642.930 2189.090 1644.110 2190.270 ;
        RECT 1642.930 2187.490 1644.110 2188.670 ;
        RECT 1642.930 2009.090 1644.110 2010.270 ;
        RECT 1642.930 2007.490 1644.110 2008.670 ;
        RECT 1642.930 1829.090 1644.110 1830.270 ;
        RECT 1642.930 1827.490 1644.110 1828.670 ;
        RECT 1642.930 1649.090 1644.110 1650.270 ;
        RECT 1642.930 1647.490 1644.110 1648.670 ;
        RECT 1642.930 1469.090 1644.110 1470.270 ;
        RECT 1642.930 1467.490 1644.110 1468.670 ;
        RECT 1642.930 1289.090 1644.110 1290.270 ;
        RECT 1642.930 1287.490 1644.110 1288.670 ;
        RECT 1642.930 1109.090 1644.110 1110.270 ;
        RECT 1642.930 1107.490 1644.110 1108.670 ;
        RECT 1642.930 929.090 1644.110 930.270 ;
        RECT 1642.930 927.490 1644.110 928.670 ;
        RECT 1642.930 749.090 1644.110 750.270 ;
        RECT 1642.930 747.490 1644.110 748.670 ;
        RECT 1642.930 569.090 1644.110 570.270 ;
        RECT 1642.930 567.490 1644.110 568.670 ;
        RECT 1642.930 389.090 1644.110 390.270 ;
        RECT 1642.930 387.490 1644.110 388.670 ;
        RECT 1642.930 209.090 1644.110 210.270 ;
        RECT 1642.930 207.490 1644.110 208.670 ;
        RECT 1642.930 29.090 1644.110 30.270 ;
        RECT 1642.930 27.490 1644.110 28.670 ;
        RECT 1642.930 -12.110 1644.110 -10.930 ;
        RECT 1642.930 -13.710 1644.110 -12.530 ;
        RECT 1822.930 3532.210 1824.110 3533.390 ;
        RECT 1822.930 3530.610 1824.110 3531.790 ;
        RECT 1822.930 3449.090 1824.110 3450.270 ;
        RECT 1822.930 3447.490 1824.110 3448.670 ;
        RECT 1822.930 3269.090 1824.110 3270.270 ;
        RECT 1822.930 3267.490 1824.110 3268.670 ;
        RECT 1822.930 3089.090 1824.110 3090.270 ;
        RECT 1822.930 3087.490 1824.110 3088.670 ;
        RECT 1822.930 2909.090 1824.110 2910.270 ;
        RECT 1822.930 2907.490 1824.110 2908.670 ;
        RECT 1822.930 2729.090 1824.110 2730.270 ;
        RECT 1822.930 2727.490 1824.110 2728.670 ;
        RECT 1822.930 2549.090 1824.110 2550.270 ;
        RECT 1822.930 2547.490 1824.110 2548.670 ;
        RECT 1822.930 2369.090 1824.110 2370.270 ;
        RECT 1822.930 2367.490 1824.110 2368.670 ;
        RECT 1822.930 2189.090 1824.110 2190.270 ;
        RECT 1822.930 2187.490 1824.110 2188.670 ;
        RECT 1822.930 2009.090 1824.110 2010.270 ;
        RECT 1822.930 2007.490 1824.110 2008.670 ;
        RECT 1822.930 1829.090 1824.110 1830.270 ;
        RECT 1822.930 1827.490 1824.110 1828.670 ;
        RECT 1822.930 1649.090 1824.110 1650.270 ;
        RECT 1822.930 1647.490 1824.110 1648.670 ;
        RECT 1822.930 1469.090 1824.110 1470.270 ;
        RECT 1822.930 1467.490 1824.110 1468.670 ;
        RECT 1822.930 1289.090 1824.110 1290.270 ;
        RECT 1822.930 1287.490 1824.110 1288.670 ;
        RECT 1822.930 1109.090 1824.110 1110.270 ;
        RECT 1822.930 1107.490 1824.110 1108.670 ;
        RECT 1822.930 929.090 1824.110 930.270 ;
        RECT 1822.930 927.490 1824.110 928.670 ;
        RECT 1822.930 749.090 1824.110 750.270 ;
        RECT 1822.930 747.490 1824.110 748.670 ;
        RECT 1822.930 569.090 1824.110 570.270 ;
        RECT 1822.930 567.490 1824.110 568.670 ;
        RECT 1822.930 389.090 1824.110 390.270 ;
        RECT 1822.930 387.490 1824.110 388.670 ;
        RECT 1822.930 209.090 1824.110 210.270 ;
        RECT 1822.930 207.490 1824.110 208.670 ;
        RECT 1822.930 29.090 1824.110 30.270 ;
        RECT 1822.930 27.490 1824.110 28.670 ;
        RECT 1822.930 -12.110 1824.110 -10.930 ;
        RECT 1822.930 -13.710 1824.110 -12.530 ;
        RECT 2002.930 3532.210 2004.110 3533.390 ;
        RECT 2002.930 3530.610 2004.110 3531.790 ;
        RECT 2002.930 3449.090 2004.110 3450.270 ;
        RECT 2002.930 3447.490 2004.110 3448.670 ;
        RECT 2002.930 3269.090 2004.110 3270.270 ;
        RECT 2002.930 3267.490 2004.110 3268.670 ;
        RECT 2002.930 3089.090 2004.110 3090.270 ;
        RECT 2002.930 3087.490 2004.110 3088.670 ;
        RECT 2002.930 2909.090 2004.110 2910.270 ;
        RECT 2002.930 2907.490 2004.110 2908.670 ;
        RECT 2002.930 2729.090 2004.110 2730.270 ;
        RECT 2002.930 2727.490 2004.110 2728.670 ;
        RECT 2002.930 2549.090 2004.110 2550.270 ;
        RECT 2002.930 2547.490 2004.110 2548.670 ;
        RECT 2002.930 2369.090 2004.110 2370.270 ;
        RECT 2002.930 2367.490 2004.110 2368.670 ;
        RECT 2002.930 2189.090 2004.110 2190.270 ;
        RECT 2002.930 2187.490 2004.110 2188.670 ;
        RECT 2002.930 2009.090 2004.110 2010.270 ;
        RECT 2002.930 2007.490 2004.110 2008.670 ;
        RECT 2002.930 1829.090 2004.110 1830.270 ;
        RECT 2002.930 1827.490 2004.110 1828.670 ;
        RECT 2002.930 1649.090 2004.110 1650.270 ;
        RECT 2002.930 1647.490 2004.110 1648.670 ;
        RECT 2002.930 1469.090 2004.110 1470.270 ;
        RECT 2002.930 1467.490 2004.110 1468.670 ;
        RECT 2002.930 1289.090 2004.110 1290.270 ;
        RECT 2002.930 1287.490 2004.110 1288.670 ;
        RECT 2002.930 1109.090 2004.110 1110.270 ;
        RECT 2002.930 1107.490 2004.110 1108.670 ;
        RECT 2002.930 929.090 2004.110 930.270 ;
        RECT 2002.930 927.490 2004.110 928.670 ;
        RECT 2002.930 749.090 2004.110 750.270 ;
        RECT 2002.930 747.490 2004.110 748.670 ;
        RECT 2002.930 569.090 2004.110 570.270 ;
        RECT 2002.930 567.490 2004.110 568.670 ;
        RECT 2002.930 389.090 2004.110 390.270 ;
        RECT 2002.930 387.490 2004.110 388.670 ;
        RECT 2002.930 209.090 2004.110 210.270 ;
        RECT 2002.930 207.490 2004.110 208.670 ;
        RECT 2002.930 29.090 2004.110 30.270 ;
        RECT 2002.930 27.490 2004.110 28.670 ;
        RECT 2002.930 -12.110 2004.110 -10.930 ;
        RECT 2002.930 -13.710 2004.110 -12.530 ;
        RECT 2182.930 3532.210 2184.110 3533.390 ;
        RECT 2182.930 3530.610 2184.110 3531.790 ;
        RECT 2182.930 3449.090 2184.110 3450.270 ;
        RECT 2182.930 3447.490 2184.110 3448.670 ;
        RECT 2182.930 3269.090 2184.110 3270.270 ;
        RECT 2182.930 3267.490 2184.110 3268.670 ;
        RECT 2182.930 3089.090 2184.110 3090.270 ;
        RECT 2182.930 3087.490 2184.110 3088.670 ;
        RECT 2182.930 2909.090 2184.110 2910.270 ;
        RECT 2182.930 2907.490 2184.110 2908.670 ;
        RECT 2182.930 2729.090 2184.110 2730.270 ;
        RECT 2182.930 2727.490 2184.110 2728.670 ;
        RECT 2182.930 2549.090 2184.110 2550.270 ;
        RECT 2182.930 2547.490 2184.110 2548.670 ;
        RECT 2182.930 2369.090 2184.110 2370.270 ;
        RECT 2182.930 2367.490 2184.110 2368.670 ;
        RECT 2182.930 2189.090 2184.110 2190.270 ;
        RECT 2182.930 2187.490 2184.110 2188.670 ;
        RECT 2182.930 2009.090 2184.110 2010.270 ;
        RECT 2182.930 2007.490 2184.110 2008.670 ;
        RECT 2182.930 1829.090 2184.110 1830.270 ;
        RECT 2182.930 1827.490 2184.110 1828.670 ;
        RECT 2182.930 1649.090 2184.110 1650.270 ;
        RECT 2182.930 1647.490 2184.110 1648.670 ;
        RECT 2182.930 1469.090 2184.110 1470.270 ;
        RECT 2182.930 1467.490 2184.110 1468.670 ;
        RECT 2182.930 1289.090 2184.110 1290.270 ;
        RECT 2182.930 1287.490 2184.110 1288.670 ;
        RECT 2182.930 1109.090 2184.110 1110.270 ;
        RECT 2182.930 1107.490 2184.110 1108.670 ;
        RECT 2182.930 929.090 2184.110 930.270 ;
        RECT 2182.930 927.490 2184.110 928.670 ;
        RECT 2182.930 749.090 2184.110 750.270 ;
        RECT 2182.930 747.490 2184.110 748.670 ;
        RECT 2182.930 569.090 2184.110 570.270 ;
        RECT 2182.930 567.490 2184.110 568.670 ;
        RECT 2182.930 389.090 2184.110 390.270 ;
        RECT 2182.930 387.490 2184.110 388.670 ;
        RECT 2182.930 209.090 2184.110 210.270 ;
        RECT 2182.930 207.490 2184.110 208.670 ;
        RECT 2182.930 29.090 2184.110 30.270 ;
        RECT 2182.930 27.490 2184.110 28.670 ;
        RECT 2182.930 -12.110 2184.110 -10.930 ;
        RECT 2182.930 -13.710 2184.110 -12.530 ;
        RECT 2362.930 3532.210 2364.110 3533.390 ;
        RECT 2362.930 3530.610 2364.110 3531.790 ;
        RECT 2362.930 3449.090 2364.110 3450.270 ;
        RECT 2362.930 3447.490 2364.110 3448.670 ;
        RECT 2362.930 3269.090 2364.110 3270.270 ;
        RECT 2362.930 3267.490 2364.110 3268.670 ;
        RECT 2362.930 3089.090 2364.110 3090.270 ;
        RECT 2362.930 3087.490 2364.110 3088.670 ;
        RECT 2362.930 2909.090 2364.110 2910.270 ;
        RECT 2362.930 2907.490 2364.110 2908.670 ;
        RECT 2362.930 2729.090 2364.110 2730.270 ;
        RECT 2362.930 2727.490 2364.110 2728.670 ;
        RECT 2362.930 2549.090 2364.110 2550.270 ;
        RECT 2362.930 2547.490 2364.110 2548.670 ;
        RECT 2362.930 2369.090 2364.110 2370.270 ;
        RECT 2362.930 2367.490 2364.110 2368.670 ;
        RECT 2362.930 2189.090 2364.110 2190.270 ;
        RECT 2362.930 2187.490 2364.110 2188.670 ;
        RECT 2362.930 2009.090 2364.110 2010.270 ;
        RECT 2362.930 2007.490 2364.110 2008.670 ;
        RECT 2362.930 1829.090 2364.110 1830.270 ;
        RECT 2362.930 1827.490 2364.110 1828.670 ;
        RECT 2362.930 1649.090 2364.110 1650.270 ;
        RECT 2362.930 1647.490 2364.110 1648.670 ;
        RECT 2362.930 1469.090 2364.110 1470.270 ;
        RECT 2362.930 1467.490 2364.110 1468.670 ;
        RECT 2362.930 1289.090 2364.110 1290.270 ;
        RECT 2362.930 1287.490 2364.110 1288.670 ;
        RECT 2362.930 1109.090 2364.110 1110.270 ;
        RECT 2362.930 1107.490 2364.110 1108.670 ;
        RECT 2362.930 929.090 2364.110 930.270 ;
        RECT 2362.930 927.490 2364.110 928.670 ;
        RECT 2362.930 749.090 2364.110 750.270 ;
        RECT 2362.930 747.490 2364.110 748.670 ;
        RECT 2362.930 569.090 2364.110 570.270 ;
        RECT 2362.930 567.490 2364.110 568.670 ;
        RECT 2362.930 389.090 2364.110 390.270 ;
        RECT 2362.930 387.490 2364.110 388.670 ;
        RECT 2362.930 209.090 2364.110 210.270 ;
        RECT 2362.930 207.490 2364.110 208.670 ;
        RECT 2362.930 29.090 2364.110 30.270 ;
        RECT 2362.930 27.490 2364.110 28.670 ;
        RECT 2362.930 -12.110 2364.110 -10.930 ;
        RECT 2362.930 -13.710 2364.110 -12.530 ;
        RECT 2542.930 3532.210 2544.110 3533.390 ;
        RECT 2542.930 3530.610 2544.110 3531.790 ;
        RECT 2542.930 3449.090 2544.110 3450.270 ;
        RECT 2542.930 3447.490 2544.110 3448.670 ;
        RECT 2542.930 3269.090 2544.110 3270.270 ;
        RECT 2542.930 3267.490 2544.110 3268.670 ;
        RECT 2542.930 3089.090 2544.110 3090.270 ;
        RECT 2542.930 3087.490 2544.110 3088.670 ;
        RECT 2542.930 2909.090 2544.110 2910.270 ;
        RECT 2542.930 2907.490 2544.110 2908.670 ;
        RECT 2542.930 2729.090 2544.110 2730.270 ;
        RECT 2542.930 2727.490 2544.110 2728.670 ;
        RECT 2542.930 2549.090 2544.110 2550.270 ;
        RECT 2542.930 2547.490 2544.110 2548.670 ;
        RECT 2542.930 2369.090 2544.110 2370.270 ;
        RECT 2542.930 2367.490 2544.110 2368.670 ;
        RECT 2542.930 2189.090 2544.110 2190.270 ;
        RECT 2542.930 2187.490 2544.110 2188.670 ;
        RECT 2542.930 2009.090 2544.110 2010.270 ;
        RECT 2542.930 2007.490 2544.110 2008.670 ;
        RECT 2542.930 1829.090 2544.110 1830.270 ;
        RECT 2542.930 1827.490 2544.110 1828.670 ;
        RECT 2542.930 1649.090 2544.110 1650.270 ;
        RECT 2542.930 1647.490 2544.110 1648.670 ;
        RECT 2542.930 1469.090 2544.110 1470.270 ;
        RECT 2542.930 1467.490 2544.110 1468.670 ;
        RECT 2542.930 1289.090 2544.110 1290.270 ;
        RECT 2542.930 1287.490 2544.110 1288.670 ;
        RECT 2542.930 1109.090 2544.110 1110.270 ;
        RECT 2542.930 1107.490 2544.110 1108.670 ;
        RECT 2542.930 929.090 2544.110 930.270 ;
        RECT 2542.930 927.490 2544.110 928.670 ;
        RECT 2542.930 749.090 2544.110 750.270 ;
        RECT 2542.930 747.490 2544.110 748.670 ;
        RECT 2542.930 569.090 2544.110 570.270 ;
        RECT 2542.930 567.490 2544.110 568.670 ;
        RECT 2542.930 389.090 2544.110 390.270 ;
        RECT 2542.930 387.490 2544.110 388.670 ;
        RECT 2542.930 209.090 2544.110 210.270 ;
        RECT 2542.930 207.490 2544.110 208.670 ;
        RECT 2542.930 29.090 2544.110 30.270 ;
        RECT 2542.930 27.490 2544.110 28.670 ;
        RECT 2542.930 -12.110 2544.110 -10.930 ;
        RECT 2542.930 -13.710 2544.110 -12.530 ;
        RECT 2722.930 3532.210 2724.110 3533.390 ;
        RECT 2722.930 3530.610 2724.110 3531.790 ;
        RECT 2722.930 3449.090 2724.110 3450.270 ;
        RECT 2722.930 3447.490 2724.110 3448.670 ;
        RECT 2722.930 3269.090 2724.110 3270.270 ;
        RECT 2722.930 3267.490 2724.110 3268.670 ;
        RECT 2722.930 3089.090 2724.110 3090.270 ;
        RECT 2722.930 3087.490 2724.110 3088.670 ;
        RECT 2722.930 2909.090 2724.110 2910.270 ;
        RECT 2722.930 2907.490 2724.110 2908.670 ;
        RECT 2722.930 2729.090 2724.110 2730.270 ;
        RECT 2722.930 2727.490 2724.110 2728.670 ;
        RECT 2722.930 2549.090 2724.110 2550.270 ;
        RECT 2722.930 2547.490 2724.110 2548.670 ;
        RECT 2722.930 2369.090 2724.110 2370.270 ;
        RECT 2722.930 2367.490 2724.110 2368.670 ;
        RECT 2722.930 2189.090 2724.110 2190.270 ;
        RECT 2722.930 2187.490 2724.110 2188.670 ;
        RECT 2722.930 2009.090 2724.110 2010.270 ;
        RECT 2722.930 2007.490 2724.110 2008.670 ;
        RECT 2722.930 1829.090 2724.110 1830.270 ;
        RECT 2722.930 1827.490 2724.110 1828.670 ;
        RECT 2722.930 1649.090 2724.110 1650.270 ;
        RECT 2722.930 1647.490 2724.110 1648.670 ;
        RECT 2722.930 1469.090 2724.110 1470.270 ;
        RECT 2722.930 1467.490 2724.110 1468.670 ;
        RECT 2722.930 1289.090 2724.110 1290.270 ;
        RECT 2722.930 1287.490 2724.110 1288.670 ;
        RECT 2722.930 1109.090 2724.110 1110.270 ;
        RECT 2722.930 1107.490 2724.110 1108.670 ;
        RECT 2722.930 929.090 2724.110 930.270 ;
        RECT 2722.930 927.490 2724.110 928.670 ;
        RECT 2722.930 749.090 2724.110 750.270 ;
        RECT 2722.930 747.490 2724.110 748.670 ;
        RECT 2722.930 569.090 2724.110 570.270 ;
        RECT 2722.930 567.490 2724.110 568.670 ;
        RECT 2722.930 389.090 2724.110 390.270 ;
        RECT 2722.930 387.490 2724.110 388.670 ;
        RECT 2722.930 209.090 2724.110 210.270 ;
        RECT 2722.930 207.490 2724.110 208.670 ;
        RECT 2722.930 29.090 2724.110 30.270 ;
        RECT 2722.930 27.490 2724.110 28.670 ;
        RECT 2722.930 -12.110 2724.110 -10.930 ;
        RECT 2722.930 -13.710 2724.110 -12.530 ;
        RECT 2902.930 3532.210 2904.110 3533.390 ;
        RECT 2902.930 3530.610 2904.110 3531.790 ;
        RECT 2902.930 3449.090 2904.110 3450.270 ;
        RECT 2902.930 3447.490 2904.110 3448.670 ;
        RECT 2902.930 3269.090 2904.110 3270.270 ;
        RECT 2902.930 3267.490 2904.110 3268.670 ;
        RECT 2902.930 3089.090 2904.110 3090.270 ;
        RECT 2902.930 3087.490 2904.110 3088.670 ;
        RECT 2902.930 2909.090 2904.110 2910.270 ;
        RECT 2902.930 2907.490 2904.110 2908.670 ;
        RECT 2902.930 2729.090 2904.110 2730.270 ;
        RECT 2902.930 2727.490 2904.110 2728.670 ;
        RECT 2902.930 2549.090 2904.110 2550.270 ;
        RECT 2902.930 2547.490 2904.110 2548.670 ;
        RECT 2902.930 2369.090 2904.110 2370.270 ;
        RECT 2902.930 2367.490 2904.110 2368.670 ;
        RECT 2902.930 2189.090 2904.110 2190.270 ;
        RECT 2902.930 2187.490 2904.110 2188.670 ;
        RECT 2902.930 2009.090 2904.110 2010.270 ;
        RECT 2902.930 2007.490 2904.110 2008.670 ;
        RECT 2902.930 1829.090 2904.110 1830.270 ;
        RECT 2902.930 1827.490 2904.110 1828.670 ;
        RECT 2902.930 1649.090 2904.110 1650.270 ;
        RECT 2902.930 1647.490 2904.110 1648.670 ;
        RECT 2902.930 1469.090 2904.110 1470.270 ;
        RECT 2902.930 1467.490 2904.110 1468.670 ;
        RECT 2902.930 1289.090 2904.110 1290.270 ;
        RECT 2902.930 1287.490 2904.110 1288.670 ;
        RECT 2902.930 1109.090 2904.110 1110.270 ;
        RECT 2902.930 1107.490 2904.110 1108.670 ;
        RECT 2902.930 929.090 2904.110 930.270 ;
        RECT 2902.930 927.490 2904.110 928.670 ;
        RECT 2902.930 749.090 2904.110 750.270 ;
        RECT 2902.930 747.490 2904.110 748.670 ;
        RECT 2902.930 569.090 2904.110 570.270 ;
        RECT 2902.930 567.490 2904.110 568.670 ;
        RECT 2902.930 389.090 2904.110 390.270 ;
        RECT 2902.930 387.490 2904.110 388.670 ;
        RECT 2902.930 209.090 2904.110 210.270 ;
        RECT 2902.930 207.490 2904.110 208.670 ;
        RECT 2902.930 29.090 2904.110 30.270 ;
        RECT 2902.930 27.490 2904.110 28.670 ;
        RECT 2902.930 -12.110 2904.110 -10.930 ;
        RECT 2902.930 -13.710 2904.110 -12.530 ;
        RECT 2936.710 3532.210 2937.890 3533.390 ;
        RECT 2936.710 3530.610 2937.890 3531.790 ;
        RECT 2936.710 3449.090 2937.890 3450.270 ;
        RECT 2936.710 3447.490 2937.890 3448.670 ;
        RECT 2936.710 3269.090 2937.890 3270.270 ;
        RECT 2936.710 3267.490 2937.890 3268.670 ;
        RECT 2936.710 3089.090 2937.890 3090.270 ;
        RECT 2936.710 3087.490 2937.890 3088.670 ;
        RECT 2936.710 2909.090 2937.890 2910.270 ;
        RECT 2936.710 2907.490 2937.890 2908.670 ;
        RECT 2936.710 2729.090 2937.890 2730.270 ;
        RECT 2936.710 2727.490 2937.890 2728.670 ;
        RECT 2936.710 2549.090 2937.890 2550.270 ;
        RECT 2936.710 2547.490 2937.890 2548.670 ;
        RECT 2936.710 2369.090 2937.890 2370.270 ;
        RECT 2936.710 2367.490 2937.890 2368.670 ;
        RECT 2936.710 2189.090 2937.890 2190.270 ;
        RECT 2936.710 2187.490 2937.890 2188.670 ;
        RECT 2936.710 2009.090 2937.890 2010.270 ;
        RECT 2936.710 2007.490 2937.890 2008.670 ;
        RECT 2936.710 1829.090 2937.890 1830.270 ;
        RECT 2936.710 1827.490 2937.890 1828.670 ;
        RECT 2936.710 1649.090 2937.890 1650.270 ;
        RECT 2936.710 1647.490 2937.890 1648.670 ;
        RECT 2936.710 1469.090 2937.890 1470.270 ;
        RECT 2936.710 1467.490 2937.890 1468.670 ;
        RECT 2936.710 1289.090 2937.890 1290.270 ;
        RECT 2936.710 1287.490 2937.890 1288.670 ;
        RECT 2936.710 1109.090 2937.890 1110.270 ;
        RECT 2936.710 1107.490 2937.890 1108.670 ;
        RECT 2936.710 929.090 2937.890 930.270 ;
        RECT 2936.710 927.490 2937.890 928.670 ;
        RECT 2936.710 749.090 2937.890 750.270 ;
        RECT 2936.710 747.490 2937.890 748.670 ;
        RECT 2936.710 569.090 2937.890 570.270 ;
        RECT 2936.710 567.490 2937.890 568.670 ;
        RECT 2936.710 389.090 2937.890 390.270 ;
        RECT 2936.710 387.490 2937.890 388.670 ;
        RECT 2936.710 209.090 2937.890 210.270 ;
        RECT 2936.710 207.490 2937.890 208.670 ;
        RECT 2936.710 29.090 2937.890 30.270 ;
        RECT 2936.710 27.490 2937.890 28.670 ;
        RECT 2936.710 -12.110 2937.890 -10.930 ;
        RECT 2936.710 -13.710 2937.890 -12.530 ;
      LAYER met5 ;
        RECT -19.180 3533.500 -16.180 3533.510 ;
        RECT 22.020 3533.500 25.020 3533.510 ;
        RECT 202.020 3533.500 205.020 3533.510 ;
        RECT 382.020 3533.500 385.020 3533.510 ;
        RECT 562.020 3533.500 565.020 3533.510 ;
        RECT 742.020 3533.500 745.020 3533.510 ;
        RECT 922.020 3533.500 925.020 3533.510 ;
        RECT 1102.020 3533.500 1105.020 3533.510 ;
        RECT 1282.020 3533.500 1285.020 3533.510 ;
        RECT 1462.020 3533.500 1465.020 3533.510 ;
        RECT 1642.020 3533.500 1645.020 3533.510 ;
        RECT 1822.020 3533.500 1825.020 3533.510 ;
        RECT 2002.020 3533.500 2005.020 3533.510 ;
        RECT 2182.020 3533.500 2185.020 3533.510 ;
        RECT 2362.020 3533.500 2365.020 3533.510 ;
        RECT 2542.020 3533.500 2545.020 3533.510 ;
        RECT 2722.020 3533.500 2725.020 3533.510 ;
        RECT 2902.020 3533.500 2905.020 3533.510 ;
        RECT 2935.800 3533.500 2938.800 3533.510 ;
        RECT -19.180 3530.500 2938.800 3533.500 ;
        RECT -19.180 3530.490 -16.180 3530.500 ;
        RECT 22.020 3530.490 25.020 3530.500 ;
        RECT 202.020 3530.490 205.020 3530.500 ;
        RECT 382.020 3530.490 385.020 3530.500 ;
        RECT 562.020 3530.490 565.020 3530.500 ;
        RECT 742.020 3530.490 745.020 3530.500 ;
        RECT 922.020 3530.490 925.020 3530.500 ;
        RECT 1102.020 3530.490 1105.020 3530.500 ;
        RECT 1282.020 3530.490 1285.020 3530.500 ;
        RECT 1462.020 3530.490 1465.020 3530.500 ;
        RECT 1642.020 3530.490 1645.020 3530.500 ;
        RECT 1822.020 3530.490 1825.020 3530.500 ;
        RECT 2002.020 3530.490 2005.020 3530.500 ;
        RECT 2182.020 3530.490 2185.020 3530.500 ;
        RECT 2362.020 3530.490 2365.020 3530.500 ;
        RECT 2542.020 3530.490 2545.020 3530.500 ;
        RECT 2722.020 3530.490 2725.020 3530.500 ;
        RECT 2902.020 3530.490 2905.020 3530.500 ;
        RECT 2935.800 3530.490 2938.800 3530.500 ;
        RECT -19.180 3450.380 -16.180 3450.390 ;
        RECT 22.020 3450.380 25.020 3450.390 ;
        RECT 202.020 3450.380 205.020 3450.390 ;
        RECT 382.020 3450.380 385.020 3450.390 ;
        RECT 562.020 3450.380 565.020 3450.390 ;
        RECT 742.020 3450.380 745.020 3450.390 ;
        RECT 922.020 3450.380 925.020 3450.390 ;
        RECT 1102.020 3450.380 1105.020 3450.390 ;
        RECT 1282.020 3450.380 1285.020 3450.390 ;
        RECT 1462.020 3450.380 1465.020 3450.390 ;
        RECT 1642.020 3450.380 1645.020 3450.390 ;
        RECT 1822.020 3450.380 1825.020 3450.390 ;
        RECT 2002.020 3450.380 2005.020 3450.390 ;
        RECT 2182.020 3450.380 2185.020 3450.390 ;
        RECT 2362.020 3450.380 2365.020 3450.390 ;
        RECT 2542.020 3450.380 2545.020 3450.390 ;
        RECT 2722.020 3450.380 2725.020 3450.390 ;
        RECT 2902.020 3450.380 2905.020 3450.390 ;
        RECT 2935.800 3450.380 2938.800 3450.390 ;
        RECT -23.780 3447.380 2943.400 3450.380 ;
        RECT -19.180 3447.370 -16.180 3447.380 ;
        RECT 22.020 3447.370 25.020 3447.380 ;
        RECT 202.020 3447.370 205.020 3447.380 ;
        RECT 382.020 3447.370 385.020 3447.380 ;
        RECT 562.020 3447.370 565.020 3447.380 ;
        RECT 742.020 3447.370 745.020 3447.380 ;
        RECT 922.020 3447.370 925.020 3447.380 ;
        RECT 1102.020 3447.370 1105.020 3447.380 ;
        RECT 1282.020 3447.370 1285.020 3447.380 ;
        RECT 1462.020 3447.370 1465.020 3447.380 ;
        RECT 1642.020 3447.370 1645.020 3447.380 ;
        RECT 1822.020 3447.370 1825.020 3447.380 ;
        RECT 2002.020 3447.370 2005.020 3447.380 ;
        RECT 2182.020 3447.370 2185.020 3447.380 ;
        RECT 2362.020 3447.370 2365.020 3447.380 ;
        RECT 2542.020 3447.370 2545.020 3447.380 ;
        RECT 2722.020 3447.370 2725.020 3447.380 ;
        RECT 2902.020 3447.370 2905.020 3447.380 ;
        RECT 2935.800 3447.370 2938.800 3447.380 ;
        RECT -19.180 3270.380 -16.180 3270.390 ;
        RECT 22.020 3270.380 25.020 3270.390 ;
        RECT 202.020 3270.380 205.020 3270.390 ;
        RECT 382.020 3270.380 385.020 3270.390 ;
        RECT 562.020 3270.380 565.020 3270.390 ;
        RECT 742.020 3270.380 745.020 3270.390 ;
        RECT 922.020 3270.380 925.020 3270.390 ;
        RECT 1102.020 3270.380 1105.020 3270.390 ;
        RECT 1282.020 3270.380 1285.020 3270.390 ;
        RECT 1462.020 3270.380 1465.020 3270.390 ;
        RECT 1642.020 3270.380 1645.020 3270.390 ;
        RECT 1822.020 3270.380 1825.020 3270.390 ;
        RECT 2002.020 3270.380 2005.020 3270.390 ;
        RECT 2182.020 3270.380 2185.020 3270.390 ;
        RECT 2362.020 3270.380 2365.020 3270.390 ;
        RECT 2542.020 3270.380 2545.020 3270.390 ;
        RECT 2722.020 3270.380 2725.020 3270.390 ;
        RECT 2902.020 3270.380 2905.020 3270.390 ;
        RECT 2935.800 3270.380 2938.800 3270.390 ;
        RECT -23.780 3267.380 2943.400 3270.380 ;
        RECT -19.180 3267.370 -16.180 3267.380 ;
        RECT 22.020 3267.370 25.020 3267.380 ;
        RECT 202.020 3267.370 205.020 3267.380 ;
        RECT 382.020 3267.370 385.020 3267.380 ;
        RECT 562.020 3267.370 565.020 3267.380 ;
        RECT 742.020 3267.370 745.020 3267.380 ;
        RECT 922.020 3267.370 925.020 3267.380 ;
        RECT 1102.020 3267.370 1105.020 3267.380 ;
        RECT 1282.020 3267.370 1285.020 3267.380 ;
        RECT 1462.020 3267.370 1465.020 3267.380 ;
        RECT 1642.020 3267.370 1645.020 3267.380 ;
        RECT 1822.020 3267.370 1825.020 3267.380 ;
        RECT 2002.020 3267.370 2005.020 3267.380 ;
        RECT 2182.020 3267.370 2185.020 3267.380 ;
        RECT 2362.020 3267.370 2365.020 3267.380 ;
        RECT 2542.020 3267.370 2545.020 3267.380 ;
        RECT 2722.020 3267.370 2725.020 3267.380 ;
        RECT 2902.020 3267.370 2905.020 3267.380 ;
        RECT 2935.800 3267.370 2938.800 3267.380 ;
        RECT -19.180 3090.380 -16.180 3090.390 ;
        RECT 22.020 3090.380 25.020 3090.390 ;
        RECT 202.020 3090.380 205.020 3090.390 ;
        RECT 382.020 3090.380 385.020 3090.390 ;
        RECT 562.020 3090.380 565.020 3090.390 ;
        RECT 742.020 3090.380 745.020 3090.390 ;
        RECT 922.020 3090.380 925.020 3090.390 ;
        RECT 1102.020 3090.380 1105.020 3090.390 ;
        RECT 1282.020 3090.380 1285.020 3090.390 ;
        RECT 1462.020 3090.380 1465.020 3090.390 ;
        RECT 1642.020 3090.380 1645.020 3090.390 ;
        RECT 1822.020 3090.380 1825.020 3090.390 ;
        RECT 2002.020 3090.380 2005.020 3090.390 ;
        RECT 2182.020 3090.380 2185.020 3090.390 ;
        RECT 2362.020 3090.380 2365.020 3090.390 ;
        RECT 2542.020 3090.380 2545.020 3090.390 ;
        RECT 2722.020 3090.380 2725.020 3090.390 ;
        RECT 2902.020 3090.380 2905.020 3090.390 ;
        RECT 2935.800 3090.380 2938.800 3090.390 ;
        RECT -23.780 3087.380 2943.400 3090.380 ;
        RECT -19.180 3087.370 -16.180 3087.380 ;
        RECT 22.020 3087.370 25.020 3087.380 ;
        RECT 202.020 3087.370 205.020 3087.380 ;
        RECT 382.020 3087.370 385.020 3087.380 ;
        RECT 562.020 3087.370 565.020 3087.380 ;
        RECT 742.020 3087.370 745.020 3087.380 ;
        RECT 922.020 3087.370 925.020 3087.380 ;
        RECT 1102.020 3087.370 1105.020 3087.380 ;
        RECT 1282.020 3087.370 1285.020 3087.380 ;
        RECT 1462.020 3087.370 1465.020 3087.380 ;
        RECT 1642.020 3087.370 1645.020 3087.380 ;
        RECT 1822.020 3087.370 1825.020 3087.380 ;
        RECT 2002.020 3087.370 2005.020 3087.380 ;
        RECT 2182.020 3087.370 2185.020 3087.380 ;
        RECT 2362.020 3087.370 2365.020 3087.380 ;
        RECT 2542.020 3087.370 2545.020 3087.380 ;
        RECT 2722.020 3087.370 2725.020 3087.380 ;
        RECT 2902.020 3087.370 2905.020 3087.380 ;
        RECT 2935.800 3087.370 2938.800 3087.380 ;
        RECT -19.180 2910.380 -16.180 2910.390 ;
        RECT 22.020 2910.380 25.020 2910.390 ;
        RECT 202.020 2910.380 205.020 2910.390 ;
        RECT 382.020 2910.380 385.020 2910.390 ;
        RECT 562.020 2910.380 565.020 2910.390 ;
        RECT 742.020 2910.380 745.020 2910.390 ;
        RECT 922.020 2910.380 925.020 2910.390 ;
        RECT 1102.020 2910.380 1105.020 2910.390 ;
        RECT 1282.020 2910.380 1285.020 2910.390 ;
        RECT 1462.020 2910.380 1465.020 2910.390 ;
        RECT 1642.020 2910.380 1645.020 2910.390 ;
        RECT 1822.020 2910.380 1825.020 2910.390 ;
        RECT 2002.020 2910.380 2005.020 2910.390 ;
        RECT 2182.020 2910.380 2185.020 2910.390 ;
        RECT 2362.020 2910.380 2365.020 2910.390 ;
        RECT 2542.020 2910.380 2545.020 2910.390 ;
        RECT 2722.020 2910.380 2725.020 2910.390 ;
        RECT 2902.020 2910.380 2905.020 2910.390 ;
        RECT 2935.800 2910.380 2938.800 2910.390 ;
        RECT -23.780 2907.380 2943.400 2910.380 ;
        RECT -19.180 2907.370 -16.180 2907.380 ;
        RECT 22.020 2907.370 25.020 2907.380 ;
        RECT 202.020 2907.370 205.020 2907.380 ;
        RECT 382.020 2907.370 385.020 2907.380 ;
        RECT 562.020 2907.370 565.020 2907.380 ;
        RECT 742.020 2907.370 745.020 2907.380 ;
        RECT 922.020 2907.370 925.020 2907.380 ;
        RECT 1102.020 2907.370 1105.020 2907.380 ;
        RECT 1282.020 2907.370 1285.020 2907.380 ;
        RECT 1462.020 2907.370 1465.020 2907.380 ;
        RECT 1642.020 2907.370 1645.020 2907.380 ;
        RECT 1822.020 2907.370 1825.020 2907.380 ;
        RECT 2002.020 2907.370 2005.020 2907.380 ;
        RECT 2182.020 2907.370 2185.020 2907.380 ;
        RECT 2362.020 2907.370 2365.020 2907.380 ;
        RECT 2542.020 2907.370 2545.020 2907.380 ;
        RECT 2722.020 2907.370 2725.020 2907.380 ;
        RECT 2902.020 2907.370 2905.020 2907.380 ;
        RECT 2935.800 2907.370 2938.800 2907.380 ;
        RECT -19.180 2730.380 -16.180 2730.390 ;
        RECT 22.020 2730.380 25.020 2730.390 ;
        RECT 202.020 2730.380 205.020 2730.390 ;
        RECT 382.020 2730.380 385.020 2730.390 ;
        RECT 562.020 2730.380 565.020 2730.390 ;
        RECT 742.020 2730.380 745.020 2730.390 ;
        RECT 922.020 2730.380 925.020 2730.390 ;
        RECT 1102.020 2730.380 1105.020 2730.390 ;
        RECT 1282.020 2730.380 1285.020 2730.390 ;
        RECT 1462.020 2730.380 1465.020 2730.390 ;
        RECT 1642.020 2730.380 1645.020 2730.390 ;
        RECT 1822.020 2730.380 1825.020 2730.390 ;
        RECT 2002.020 2730.380 2005.020 2730.390 ;
        RECT 2182.020 2730.380 2185.020 2730.390 ;
        RECT 2362.020 2730.380 2365.020 2730.390 ;
        RECT 2542.020 2730.380 2545.020 2730.390 ;
        RECT 2722.020 2730.380 2725.020 2730.390 ;
        RECT 2902.020 2730.380 2905.020 2730.390 ;
        RECT 2935.800 2730.380 2938.800 2730.390 ;
        RECT -23.780 2727.380 2943.400 2730.380 ;
        RECT -19.180 2727.370 -16.180 2727.380 ;
        RECT 22.020 2727.370 25.020 2727.380 ;
        RECT 202.020 2727.370 205.020 2727.380 ;
        RECT 382.020 2727.370 385.020 2727.380 ;
        RECT 562.020 2727.370 565.020 2727.380 ;
        RECT 742.020 2727.370 745.020 2727.380 ;
        RECT 922.020 2727.370 925.020 2727.380 ;
        RECT 1102.020 2727.370 1105.020 2727.380 ;
        RECT 1282.020 2727.370 1285.020 2727.380 ;
        RECT 1462.020 2727.370 1465.020 2727.380 ;
        RECT 1642.020 2727.370 1645.020 2727.380 ;
        RECT 1822.020 2727.370 1825.020 2727.380 ;
        RECT 2002.020 2727.370 2005.020 2727.380 ;
        RECT 2182.020 2727.370 2185.020 2727.380 ;
        RECT 2362.020 2727.370 2365.020 2727.380 ;
        RECT 2542.020 2727.370 2545.020 2727.380 ;
        RECT 2722.020 2727.370 2725.020 2727.380 ;
        RECT 2902.020 2727.370 2905.020 2727.380 ;
        RECT 2935.800 2727.370 2938.800 2727.380 ;
        RECT -19.180 2550.380 -16.180 2550.390 ;
        RECT 22.020 2550.380 25.020 2550.390 ;
        RECT 202.020 2550.380 205.020 2550.390 ;
        RECT 382.020 2550.380 385.020 2550.390 ;
        RECT 562.020 2550.380 565.020 2550.390 ;
        RECT 742.020 2550.380 745.020 2550.390 ;
        RECT 922.020 2550.380 925.020 2550.390 ;
        RECT 1102.020 2550.380 1105.020 2550.390 ;
        RECT 1282.020 2550.380 1285.020 2550.390 ;
        RECT 1462.020 2550.380 1465.020 2550.390 ;
        RECT 1642.020 2550.380 1645.020 2550.390 ;
        RECT 1822.020 2550.380 1825.020 2550.390 ;
        RECT 2002.020 2550.380 2005.020 2550.390 ;
        RECT 2182.020 2550.380 2185.020 2550.390 ;
        RECT 2362.020 2550.380 2365.020 2550.390 ;
        RECT 2542.020 2550.380 2545.020 2550.390 ;
        RECT 2722.020 2550.380 2725.020 2550.390 ;
        RECT 2902.020 2550.380 2905.020 2550.390 ;
        RECT 2935.800 2550.380 2938.800 2550.390 ;
        RECT -23.780 2547.380 2943.400 2550.380 ;
        RECT -19.180 2547.370 -16.180 2547.380 ;
        RECT 22.020 2547.370 25.020 2547.380 ;
        RECT 202.020 2547.370 205.020 2547.380 ;
        RECT 382.020 2547.370 385.020 2547.380 ;
        RECT 562.020 2547.370 565.020 2547.380 ;
        RECT 742.020 2547.370 745.020 2547.380 ;
        RECT 922.020 2547.370 925.020 2547.380 ;
        RECT 1102.020 2547.370 1105.020 2547.380 ;
        RECT 1282.020 2547.370 1285.020 2547.380 ;
        RECT 1462.020 2547.370 1465.020 2547.380 ;
        RECT 1642.020 2547.370 1645.020 2547.380 ;
        RECT 1822.020 2547.370 1825.020 2547.380 ;
        RECT 2002.020 2547.370 2005.020 2547.380 ;
        RECT 2182.020 2547.370 2185.020 2547.380 ;
        RECT 2362.020 2547.370 2365.020 2547.380 ;
        RECT 2542.020 2547.370 2545.020 2547.380 ;
        RECT 2722.020 2547.370 2725.020 2547.380 ;
        RECT 2902.020 2547.370 2905.020 2547.380 ;
        RECT 2935.800 2547.370 2938.800 2547.380 ;
        RECT -19.180 2370.380 -16.180 2370.390 ;
        RECT 22.020 2370.380 25.020 2370.390 ;
        RECT 202.020 2370.380 205.020 2370.390 ;
        RECT 382.020 2370.380 385.020 2370.390 ;
        RECT 562.020 2370.380 565.020 2370.390 ;
        RECT 742.020 2370.380 745.020 2370.390 ;
        RECT 922.020 2370.380 925.020 2370.390 ;
        RECT 1102.020 2370.380 1105.020 2370.390 ;
        RECT 1282.020 2370.380 1285.020 2370.390 ;
        RECT 1462.020 2370.380 1465.020 2370.390 ;
        RECT 1642.020 2370.380 1645.020 2370.390 ;
        RECT 1822.020 2370.380 1825.020 2370.390 ;
        RECT 2002.020 2370.380 2005.020 2370.390 ;
        RECT 2182.020 2370.380 2185.020 2370.390 ;
        RECT 2362.020 2370.380 2365.020 2370.390 ;
        RECT 2542.020 2370.380 2545.020 2370.390 ;
        RECT 2722.020 2370.380 2725.020 2370.390 ;
        RECT 2902.020 2370.380 2905.020 2370.390 ;
        RECT 2935.800 2370.380 2938.800 2370.390 ;
        RECT -23.780 2367.380 2943.400 2370.380 ;
        RECT -19.180 2367.370 -16.180 2367.380 ;
        RECT 22.020 2367.370 25.020 2367.380 ;
        RECT 202.020 2367.370 205.020 2367.380 ;
        RECT 382.020 2367.370 385.020 2367.380 ;
        RECT 562.020 2367.370 565.020 2367.380 ;
        RECT 742.020 2367.370 745.020 2367.380 ;
        RECT 922.020 2367.370 925.020 2367.380 ;
        RECT 1102.020 2367.370 1105.020 2367.380 ;
        RECT 1282.020 2367.370 1285.020 2367.380 ;
        RECT 1462.020 2367.370 1465.020 2367.380 ;
        RECT 1642.020 2367.370 1645.020 2367.380 ;
        RECT 1822.020 2367.370 1825.020 2367.380 ;
        RECT 2002.020 2367.370 2005.020 2367.380 ;
        RECT 2182.020 2367.370 2185.020 2367.380 ;
        RECT 2362.020 2367.370 2365.020 2367.380 ;
        RECT 2542.020 2367.370 2545.020 2367.380 ;
        RECT 2722.020 2367.370 2725.020 2367.380 ;
        RECT 2902.020 2367.370 2905.020 2367.380 ;
        RECT 2935.800 2367.370 2938.800 2367.380 ;
        RECT -19.180 2190.380 -16.180 2190.390 ;
        RECT 22.020 2190.380 25.020 2190.390 ;
        RECT 202.020 2190.380 205.020 2190.390 ;
        RECT 382.020 2190.380 385.020 2190.390 ;
        RECT 562.020 2190.380 565.020 2190.390 ;
        RECT 742.020 2190.380 745.020 2190.390 ;
        RECT 922.020 2190.380 925.020 2190.390 ;
        RECT 1102.020 2190.380 1105.020 2190.390 ;
        RECT 1282.020 2190.380 1285.020 2190.390 ;
        RECT 1462.020 2190.380 1465.020 2190.390 ;
        RECT 1642.020 2190.380 1645.020 2190.390 ;
        RECT 1822.020 2190.380 1825.020 2190.390 ;
        RECT 2002.020 2190.380 2005.020 2190.390 ;
        RECT 2182.020 2190.380 2185.020 2190.390 ;
        RECT 2362.020 2190.380 2365.020 2190.390 ;
        RECT 2542.020 2190.380 2545.020 2190.390 ;
        RECT 2722.020 2190.380 2725.020 2190.390 ;
        RECT 2902.020 2190.380 2905.020 2190.390 ;
        RECT 2935.800 2190.380 2938.800 2190.390 ;
        RECT -23.780 2187.380 2943.400 2190.380 ;
        RECT -19.180 2187.370 -16.180 2187.380 ;
        RECT 22.020 2187.370 25.020 2187.380 ;
        RECT 202.020 2187.370 205.020 2187.380 ;
        RECT 382.020 2187.370 385.020 2187.380 ;
        RECT 562.020 2187.370 565.020 2187.380 ;
        RECT 742.020 2187.370 745.020 2187.380 ;
        RECT 922.020 2187.370 925.020 2187.380 ;
        RECT 1102.020 2187.370 1105.020 2187.380 ;
        RECT 1282.020 2187.370 1285.020 2187.380 ;
        RECT 1462.020 2187.370 1465.020 2187.380 ;
        RECT 1642.020 2187.370 1645.020 2187.380 ;
        RECT 1822.020 2187.370 1825.020 2187.380 ;
        RECT 2002.020 2187.370 2005.020 2187.380 ;
        RECT 2182.020 2187.370 2185.020 2187.380 ;
        RECT 2362.020 2187.370 2365.020 2187.380 ;
        RECT 2542.020 2187.370 2545.020 2187.380 ;
        RECT 2722.020 2187.370 2725.020 2187.380 ;
        RECT 2902.020 2187.370 2905.020 2187.380 ;
        RECT 2935.800 2187.370 2938.800 2187.380 ;
        RECT -19.180 2010.380 -16.180 2010.390 ;
        RECT 22.020 2010.380 25.020 2010.390 ;
        RECT 202.020 2010.380 205.020 2010.390 ;
        RECT 382.020 2010.380 385.020 2010.390 ;
        RECT 562.020 2010.380 565.020 2010.390 ;
        RECT 742.020 2010.380 745.020 2010.390 ;
        RECT 922.020 2010.380 925.020 2010.390 ;
        RECT 1102.020 2010.380 1105.020 2010.390 ;
        RECT 1282.020 2010.380 1285.020 2010.390 ;
        RECT 1462.020 2010.380 1465.020 2010.390 ;
        RECT 1642.020 2010.380 1645.020 2010.390 ;
        RECT 1822.020 2010.380 1825.020 2010.390 ;
        RECT 2002.020 2010.380 2005.020 2010.390 ;
        RECT 2182.020 2010.380 2185.020 2010.390 ;
        RECT 2362.020 2010.380 2365.020 2010.390 ;
        RECT 2542.020 2010.380 2545.020 2010.390 ;
        RECT 2722.020 2010.380 2725.020 2010.390 ;
        RECT 2902.020 2010.380 2905.020 2010.390 ;
        RECT 2935.800 2010.380 2938.800 2010.390 ;
        RECT -23.780 2007.380 2943.400 2010.380 ;
        RECT -19.180 2007.370 -16.180 2007.380 ;
        RECT 22.020 2007.370 25.020 2007.380 ;
        RECT 202.020 2007.370 205.020 2007.380 ;
        RECT 382.020 2007.370 385.020 2007.380 ;
        RECT 562.020 2007.370 565.020 2007.380 ;
        RECT 742.020 2007.370 745.020 2007.380 ;
        RECT 922.020 2007.370 925.020 2007.380 ;
        RECT 1102.020 2007.370 1105.020 2007.380 ;
        RECT 1282.020 2007.370 1285.020 2007.380 ;
        RECT 1462.020 2007.370 1465.020 2007.380 ;
        RECT 1642.020 2007.370 1645.020 2007.380 ;
        RECT 1822.020 2007.370 1825.020 2007.380 ;
        RECT 2002.020 2007.370 2005.020 2007.380 ;
        RECT 2182.020 2007.370 2185.020 2007.380 ;
        RECT 2362.020 2007.370 2365.020 2007.380 ;
        RECT 2542.020 2007.370 2545.020 2007.380 ;
        RECT 2722.020 2007.370 2725.020 2007.380 ;
        RECT 2902.020 2007.370 2905.020 2007.380 ;
        RECT 2935.800 2007.370 2938.800 2007.380 ;
        RECT -19.180 1830.380 -16.180 1830.390 ;
        RECT 22.020 1830.380 25.020 1830.390 ;
        RECT 202.020 1830.380 205.020 1830.390 ;
        RECT 382.020 1830.380 385.020 1830.390 ;
        RECT 562.020 1830.380 565.020 1830.390 ;
        RECT 742.020 1830.380 745.020 1830.390 ;
        RECT 922.020 1830.380 925.020 1830.390 ;
        RECT 1102.020 1830.380 1105.020 1830.390 ;
        RECT 1282.020 1830.380 1285.020 1830.390 ;
        RECT 1462.020 1830.380 1465.020 1830.390 ;
        RECT 1642.020 1830.380 1645.020 1830.390 ;
        RECT 1822.020 1830.380 1825.020 1830.390 ;
        RECT 2002.020 1830.380 2005.020 1830.390 ;
        RECT 2182.020 1830.380 2185.020 1830.390 ;
        RECT 2362.020 1830.380 2365.020 1830.390 ;
        RECT 2542.020 1830.380 2545.020 1830.390 ;
        RECT 2722.020 1830.380 2725.020 1830.390 ;
        RECT 2902.020 1830.380 2905.020 1830.390 ;
        RECT 2935.800 1830.380 2938.800 1830.390 ;
        RECT -23.780 1827.380 2943.400 1830.380 ;
        RECT -19.180 1827.370 -16.180 1827.380 ;
        RECT 22.020 1827.370 25.020 1827.380 ;
        RECT 202.020 1827.370 205.020 1827.380 ;
        RECT 382.020 1827.370 385.020 1827.380 ;
        RECT 562.020 1827.370 565.020 1827.380 ;
        RECT 742.020 1827.370 745.020 1827.380 ;
        RECT 922.020 1827.370 925.020 1827.380 ;
        RECT 1102.020 1827.370 1105.020 1827.380 ;
        RECT 1282.020 1827.370 1285.020 1827.380 ;
        RECT 1462.020 1827.370 1465.020 1827.380 ;
        RECT 1642.020 1827.370 1645.020 1827.380 ;
        RECT 1822.020 1827.370 1825.020 1827.380 ;
        RECT 2002.020 1827.370 2005.020 1827.380 ;
        RECT 2182.020 1827.370 2185.020 1827.380 ;
        RECT 2362.020 1827.370 2365.020 1827.380 ;
        RECT 2542.020 1827.370 2545.020 1827.380 ;
        RECT 2722.020 1827.370 2725.020 1827.380 ;
        RECT 2902.020 1827.370 2905.020 1827.380 ;
        RECT 2935.800 1827.370 2938.800 1827.380 ;
        RECT -19.180 1650.380 -16.180 1650.390 ;
        RECT 22.020 1650.380 25.020 1650.390 ;
        RECT 202.020 1650.380 205.020 1650.390 ;
        RECT 382.020 1650.380 385.020 1650.390 ;
        RECT 562.020 1650.380 565.020 1650.390 ;
        RECT 742.020 1650.380 745.020 1650.390 ;
        RECT 922.020 1650.380 925.020 1650.390 ;
        RECT 1102.020 1650.380 1105.020 1650.390 ;
        RECT 1282.020 1650.380 1285.020 1650.390 ;
        RECT 1462.020 1650.380 1465.020 1650.390 ;
        RECT 1642.020 1650.380 1645.020 1650.390 ;
        RECT 1822.020 1650.380 1825.020 1650.390 ;
        RECT 2002.020 1650.380 2005.020 1650.390 ;
        RECT 2182.020 1650.380 2185.020 1650.390 ;
        RECT 2362.020 1650.380 2365.020 1650.390 ;
        RECT 2542.020 1650.380 2545.020 1650.390 ;
        RECT 2722.020 1650.380 2725.020 1650.390 ;
        RECT 2902.020 1650.380 2905.020 1650.390 ;
        RECT 2935.800 1650.380 2938.800 1650.390 ;
        RECT -23.780 1647.380 2943.400 1650.380 ;
        RECT -19.180 1647.370 -16.180 1647.380 ;
        RECT 22.020 1647.370 25.020 1647.380 ;
        RECT 202.020 1647.370 205.020 1647.380 ;
        RECT 382.020 1647.370 385.020 1647.380 ;
        RECT 562.020 1647.370 565.020 1647.380 ;
        RECT 742.020 1647.370 745.020 1647.380 ;
        RECT 922.020 1647.370 925.020 1647.380 ;
        RECT 1102.020 1647.370 1105.020 1647.380 ;
        RECT 1282.020 1647.370 1285.020 1647.380 ;
        RECT 1462.020 1647.370 1465.020 1647.380 ;
        RECT 1642.020 1647.370 1645.020 1647.380 ;
        RECT 1822.020 1647.370 1825.020 1647.380 ;
        RECT 2002.020 1647.370 2005.020 1647.380 ;
        RECT 2182.020 1647.370 2185.020 1647.380 ;
        RECT 2362.020 1647.370 2365.020 1647.380 ;
        RECT 2542.020 1647.370 2545.020 1647.380 ;
        RECT 2722.020 1647.370 2725.020 1647.380 ;
        RECT 2902.020 1647.370 2905.020 1647.380 ;
        RECT 2935.800 1647.370 2938.800 1647.380 ;
        RECT -19.180 1470.380 -16.180 1470.390 ;
        RECT 22.020 1470.380 25.020 1470.390 ;
        RECT 202.020 1470.380 205.020 1470.390 ;
        RECT 382.020 1470.380 385.020 1470.390 ;
        RECT 562.020 1470.380 565.020 1470.390 ;
        RECT 742.020 1470.380 745.020 1470.390 ;
        RECT 922.020 1470.380 925.020 1470.390 ;
        RECT 1102.020 1470.380 1105.020 1470.390 ;
        RECT 1282.020 1470.380 1285.020 1470.390 ;
        RECT 1462.020 1470.380 1465.020 1470.390 ;
        RECT 1642.020 1470.380 1645.020 1470.390 ;
        RECT 1822.020 1470.380 1825.020 1470.390 ;
        RECT 2002.020 1470.380 2005.020 1470.390 ;
        RECT 2182.020 1470.380 2185.020 1470.390 ;
        RECT 2362.020 1470.380 2365.020 1470.390 ;
        RECT 2542.020 1470.380 2545.020 1470.390 ;
        RECT 2722.020 1470.380 2725.020 1470.390 ;
        RECT 2902.020 1470.380 2905.020 1470.390 ;
        RECT 2935.800 1470.380 2938.800 1470.390 ;
        RECT -23.780 1467.380 2943.400 1470.380 ;
        RECT -19.180 1467.370 -16.180 1467.380 ;
        RECT 22.020 1467.370 25.020 1467.380 ;
        RECT 202.020 1467.370 205.020 1467.380 ;
        RECT 382.020 1467.370 385.020 1467.380 ;
        RECT 562.020 1467.370 565.020 1467.380 ;
        RECT 742.020 1467.370 745.020 1467.380 ;
        RECT 922.020 1467.370 925.020 1467.380 ;
        RECT 1102.020 1467.370 1105.020 1467.380 ;
        RECT 1282.020 1467.370 1285.020 1467.380 ;
        RECT 1462.020 1467.370 1465.020 1467.380 ;
        RECT 1642.020 1467.370 1645.020 1467.380 ;
        RECT 1822.020 1467.370 1825.020 1467.380 ;
        RECT 2002.020 1467.370 2005.020 1467.380 ;
        RECT 2182.020 1467.370 2185.020 1467.380 ;
        RECT 2362.020 1467.370 2365.020 1467.380 ;
        RECT 2542.020 1467.370 2545.020 1467.380 ;
        RECT 2722.020 1467.370 2725.020 1467.380 ;
        RECT 2902.020 1467.370 2905.020 1467.380 ;
        RECT 2935.800 1467.370 2938.800 1467.380 ;
        RECT -19.180 1290.380 -16.180 1290.390 ;
        RECT 22.020 1290.380 25.020 1290.390 ;
        RECT 202.020 1290.380 205.020 1290.390 ;
        RECT 382.020 1290.380 385.020 1290.390 ;
        RECT 562.020 1290.380 565.020 1290.390 ;
        RECT 742.020 1290.380 745.020 1290.390 ;
        RECT 922.020 1290.380 925.020 1290.390 ;
        RECT 1102.020 1290.380 1105.020 1290.390 ;
        RECT 1282.020 1290.380 1285.020 1290.390 ;
        RECT 1462.020 1290.380 1465.020 1290.390 ;
        RECT 1642.020 1290.380 1645.020 1290.390 ;
        RECT 1822.020 1290.380 1825.020 1290.390 ;
        RECT 2002.020 1290.380 2005.020 1290.390 ;
        RECT 2182.020 1290.380 2185.020 1290.390 ;
        RECT 2362.020 1290.380 2365.020 1290.390 ;
        RECT 2542.020 1290.380 2545.020 1290.390 ;
        RECT 2722.020 1290.380 2725.020 1290.390 ;
        RECT 2902.020 1290.380 2905.020 1290.390 ;
        RECT 2935.800 1290.380 2938.800 1290.390 ;
        RECT -23.780 1287.380 2943.400 1290.380 ;
        RECT -19.180 1287.370 -16.180 1287.380 ;
        RECT 22.020 1287.370 25.020 1287.380 ;
        RECT 202.020 1287.370 205.020 1287.380 ;
        RECT 382.020 1287.370 385.020 1287.380 ;
        RECT 562.020 1287.370 565.020 1287.380 ;
        RECT 742.020 1287.370 745.020 1287.380 ;
        RECT 922.020 1287.370 925.020 1287.380 ;
        RECT 1102.020 1287.370 1105.020 1287.380 ;
        RECT 1282.020 1287.370 1285.020 1287.380 ;
        RECT 1462.020 1287.370 1465.020 1287.380 ;
        RECT 1642.020 1287.370 1645.020 1287.380 ;
        RECT 1822.020 1287.370 1825.020 1287.380 ;
        RECT 2002.020 1287.370 2005.020 1287.380 ;
        RECT 2182.020 1287.370 2185.020 1287.380 ;
        RECT 2362.020 1287.370 2365.020 1287.380 ;
        RECT 2542.020 1287.370 2545.020 1287.380 ;
        RECT 2722.020 1287.370 2725.020 1287.380 ;
        RECT 2902.020 1287.370 2905.020 1287.380 ;
        RECT 2935.800 1287.370 2938.800 1287.380 ;
        RECT -19.180 1110.380 -16.180 1110.390 ;
        RECT 22.020 1110.380 25.020 1110.390 ;
        RECT 202.020 1110.380 205.020 1110.390 ;
        RECT 382.020 1110.380 385.020 1110.390 ;
        RECT 562.020 1110.380 565.020 1110.390 ;
        RECT 742.020 1110.380 745.020 1110.390 ;
        RECT 922.020 1110.380 925.020 1110.390 ;
        RECT 1102.020 1110.380 1105.020 1110.390 ;
        RECT 1282.020 1110.380 1285.020 1110.390 ;
        RECT 1462.020 1110.380 1465.020 1110.390 ;
        RECT 1642.020 1110.380 1645.020 1110.390 ;
        RECT 1822.020 1110.380 1825.020 1110.390 ;
        RECT 2002.020 1110.380 2005.020 1110.390 ;
        RECT 2182.020 1110.380 2185.020 1110.390 ;
        RECT 2362.020 1110.380 2365.020 1110.390 ;
        RECT 2542.020 1110.380 2545.020 1110.390 ;
        RECT 2722.020 1110.380 2725.020 1110.390 ;
        RECT 2902.020 1110.380 2905.020 1110.390 ;
        RECT 2935.800 1110.380 2938.800 1110.390 ;
        RECT -23.780 1107.380 2943.400 1110.380 ;
        RECT -19.180 1107.370 -16.180 1107.380 ;
        RECT 22.020 1107.370 25.020 1107.380 ;
        RECT 202.020 1107.370 205.020 1107.380 ;
        RECT 382.020 1107.370 385.020 1107.380 ;
        RECT 562.020 1107.370 565.020 1107.380 ;
        RECT 742.020 1107.370 745.020 1107.380 ;
        RECT 922.020 1107.370 925.020 1107.380 ;
        RECT 1102.020 1107.370 1105.020 1107.380 ;
        RECT 1282.020 1107.370 1285.020 1107.380 ;
        RECT 1462.020 1107.370 1465.020 1107.380 ;
        RECT 1642.020 1107.370 1645.020 1107.380 ;
        RECT 1822.020 1107.370 1825.020 1107.380 ;
        RECT 2002.020 1107.370 2005.020 1107.380 ;
        RECT 2182.020 1107.370 2185.020 1107.380 ;
        RECT 2362.020 1107.370 2365.020 1107.380 ;
        RECT 2542.020 1107.370 2545.020 1107.380 ;
        RECT 2722.020 1107.370 2725.020 1107.380 ;
        RECT 2902.020 1107.370 2905.020 1107.380 ;
        RECT 2935.800 1107.370 2938.800 1107.380 ;
        RECT -19.180 930.380 -16.180 930.390 ;
        RECT 22.020 930.380 25.020 930.390 ;
        RECT 202.020 930.380 205.020 930.390 ;
        RECT 382.020 930.380 385.020 930.390 ;
        RECT 562.020 930.380 565.020 930.390 ;
        RECT 742.020 930.380 745.020 930.390 ;
        RECT 922.020 930.380 925.020 930.390 ;
        RECT 1102.020 930.380 1105.020 930.390 ;
        RECT 1282.020 930.380 1285.020 930.390 ;
        RECT 1462.020 930.380 1465.020 930.390 ;
        RECT 1642.020 930.380 1645.020 930.390 ;
        RECT 1822.020 930.380 1825.020 930.390 ;
        RECT 2002.020 930.380 2005.020 930.390 ;
        RECT 2182.020 930.380 2185.020 930.390 ;
        RECT 2362.020 930.380 2365.020 930.390 ;
        RECT 2542.020 930.380 2545.020 930.390 ;
        RECT 2722.020 930.380 2725.020 930.390 ;
        RECT 2902.020 930.380 2905.020 930.390 ;
        RECT 2935.800 930.380 2938.800 930.390 ;
        RECT -23.780 927.380 2943.400 930.380 ;
        RECT -19.180 927.370 -16.180 927.380 ;
        RECT 22.020 927.370 25.020 927.380 ;
        RECT 202.020 927.370 205.020 927.380 ;
        RECT 382.020 927.370 385.020 927.380 ;
        RECT 562.020 927.370 565.020 927.380 ;
        RECT 742.020 927.370 745.020 927.380 ;
        RECT 922.020 927.370 925.020 927.380 ;
        RECT 1102.020 927.370 1105.020 927.380 ;
        RECT 1282.020 927.370 1285.020 927.380 ;
        RECT 1462.020 927.370 1465.020 927.380 ;
        RECT 1642.020 927.370 1645.020 927.380 ;
        RECT 1822.020 927.370 1825.020 927.380 ;
        RECT 2002.020 927.370 2005.020 927.380 ;
        RECT 2182.020 927.370 2185.020 927.380 ;
        RECT 2362.020 927.370 2365.020 927.380 ;
        RECT 2542.020 927.370 2545.020 927.380 ;
        RECT 2722.020 927.370 2725.020 927.380 ;
        RECT 2902.020 927.370 2905.020 927.380 ;
        RECT 2935.800 927.370 2938.800 927.380 ;
        RECT -19.180 750.380 -16.180 750.390 ;
        RECT 22.020 750.380 25.020 750.390 ;
        RECT 202.020 750.380 205.020 750.390 ;
        RECT 382.020 750.380 385.020 750.390 ;
        RECT 562.020 750.380 565.020 750.390 ;
        RECT 742.020 750.380 745.020 750.390 ;
        RECT 922.020 750.380 925.020 750.390 ;
        RECT 1102.020 750.380 1105.020 750.390 ;
        RECT 1282.020 750.380 1285.020 750.390 ;
        RECT 1462.020 750.380 1465.020 750.390 ;
        RECT 1642.020 750.380 1645.020 750.390 ;
        RECT 1822.020 750.380 1825.020 750.390 ;
        RECT 2002.020 750.380 2005.020 750.390 ;
        RECT 2182.020 750.380 2185.020 750.390 ;
        RECT 2362.020 750.380 2365.020 750.390 ;
        RECT 2542.020 750.380 2545.020 750.390 ;
        RECT 2722.020 750.380 2725.020 750.390 ;
        RECT 2902.020 750.380 2905.020 750.390 ;
        RECT 2935.800 750.380 2938.800 750.390 ;
        RECT -23.780 747.380 2943.400 750.380 ;
        RECT -19.180 747.370 -16.180 747.380 ;
        RECT 22.020 747.370 25.020 747.380 ;
        RECT 202.020 747.370 205.020 747.380 ;
        RECT 382.020 747.370 385.020 747.380 ;
        RECT 562.020 747.370 565.020 747.380 ;
        RECT 742.020 747.370 745.020 747.380 ;
        RECT 922.020 747.370 925.020 747.380 ;
        RECT 1102.020 747.370 1105.020 747.380 ;
        RECT 1282.020 747.370 1285.020 747.380 ;
        RECT 1462.020 747.370 1465.020 747.380 ;
        RECT 1642.020 747.370 1645.020 747.380 ;
        RECT 1822.020 747.370 1825.020 747.380 ;
        RECT 2002.020 747.370 2005.020 747.380 ;
        RECT 2182.020 747.370 2185.020 747.380 ;
        RECT 2362.020 747.370 2365.020 747.380 ;
        RECT 2542.020 747.370 2545.020 747.380 ;
        RECT 2722.020 747.370 2725.020 747.380 ;
        RECT 2902.020 747.370 2905.020 747.380 ;
        RECT 2935.800 747.370 2938.800 747.380 ;
        RECT -19.180 570.380 -16.180 570.390 ;
        RECT 22.020 570.380 25.020 570.390 ;
        RECT 202.020 570.380 205.020 570.390 ;
        RECT 382.020 570.380 385.020 570.390 ;
        RECT 562.020 570.380 565.020 570.390 ;
        RECT 742.020 570.380 745.020 570.390 ;
        RECT 922.020 570.380 925.020 570.390 ;
        RECT 1102.020 570.380 1105.020 570.390 ;
        RECT 1282.020 570.380 1285.020 570.390 ;
        RECT 1462.020 570.380 1465.020 570.390 ;
        RECT 1642.020 570.380 1645.020 570.390 ;
        RECT 1822.020 570.380 1825.020 570.390 ;
        RECT 2002.020 570.380 2005.020 570.390 ;
        RECT 2182.020 570.380 2185.020 570.390 ;
        RECT 2362.020 570.380 2365.020 570.390 ;
        RECT 2542.020 570.380 2545.020 570.390 ;
        RECT 2722.020 570.380 2725.020 570.390 ;
        RECT 2902.020 570.380 2905.020 570.390 ;
        RECT 2935.800 570.380 2938.800 570.390 ;
        RECT -23.780 567.380 2943.400 570.380 ;
        RECT -19.180 567.370 -16.180 567.380 ;
        RECT 22.020 567.370 25.020 567.380 ;
        RECT 202.020 567.370 205.020 567.380 ;
        RECT 382.020 567.370 385.020 567.380 ;
        RECT 562.020 567.370 565.020 567.380 ;
        RECT 742.020 567.370 745.020 567.380 ;
        RECT 922.020 567.370 925.020 567.380 ;
        RECT 1102.020 567.370 1105.020 567.380 ;
        RECT 1282.020 567.370 1285.020 567.380 ;
        RECT 1462.020 567.370 1465.020 567.380 ;
        RECT 1642.020 567.370 1645.020 567.380 ;
        RECT 1822.020 567.370 1825.020 567.380 ;
        RECT 2002.020 567.370 2005.020 567.380 ;
        RECT 2182.020 567.370 2185.020 567.380 ;
        RECT 2362.020 567.370 2365.020 567.380 ;
        RECT 2542.020 567.370 2545.020 567.380 ;
        RECT 2722.020 567.370 2725.020 567.380 ;
        RECT 2902.020 567.370 2905.020 567.380 ;
        RECT 2935.800 567.370 2938.800 567.380 ;
        RECT -19.180 390.380 -16.180 390.390 ;
        RECT 22.020 390.380 25.020 390.390 ;
        RECT 202.020 390.380 205.020 390.390 ;
        RECT 382.020 390.380 385.020 390.390 ;
        RECT 562.020 390.380 565.020 390.390 ;
        RECT 742.020 390.380 745.020 390.390 ;
        RECT 922.020 390.380 925.020 390.390 ;
        RECT 1102.020 390.380 1105.020 390.390 ;
        RECT 1282.020 390.380 1285.020 390.390 ;
        RECT 1462.020 390.380 1465.020 390.390 ;
        RECT 1642.020 390.380 1645.020 390.390 ;
        RECT 1822.020 390.380 1825.020 390.390 ;
        RECT 2002.020 390.380 2005.020 390.390 ;
        RECT 2182.020 390.380 2185.020 390.390 ;
        RECT 2362.020 390.380 2365.020 390.390 ;
        RECT 2542.020 390.380 2545.020 390.390 ;
        RECT 2722.020 390.380 2725.020 390.390 ;
        RECT 2902.020 390.380 2905.020 390.390 ;
        RECT 2935.800 390.380 2938.800 390.390 ;
        RECT -23.780 387.380 2943.400 390.380 ;
        RECT -19.180 387.370 -16.180 387.380 ;
        RECT 22.020 387.370 25.020 387.380 ;
        RECT 202.020 387.370 205.020 387.380 ;
        RECT 382.020 387.370 385.020 387.380 ;
        RECT 562.020 387.370 565.020 387.380 ;
        RECT 742.020 387.370 745.020 387.380 ;
        RECT 922.020 387.370 925.020 387.380 ;
        RECT 1102.020 387.370 1105.020 387.380 ;
        RECT 1282.020 387.370 1285.020 387.380 ;
        RECT 1462.020 387.370 1465.020 387.380 ;
        RECT 1642.020 387.370 1645.020 387.380 ;
        RECT 1822.020 387.370 1825.020 387.380 ;
        RECT 2002.020 387.370 2005.020 387.380 ;
        RECT 2182.020 387.370 2185.020 387.380 ;
        RECT 2362.020 387.370 2365.020 387.380 ;
        RECT 2542.020 387.370 2545.020 387.380 ;
        RECT 2722.020 387.370 2725.020 387.380 ;
        RECT 2902.020 387.370 2905.020 387.380 ;
        RECT 2935.800 387.370 2938.800 387.380 ;
        RECT -19.180 210.380 -16.180 210.390 ;
        RECT 22.020 210.380 25.020 210.390 ;
        RECT 202.020 210.380 205.020 210.390 ;
        RECT 382.020 210.380 385.020 210.390 ;
        RECT 562.020 210.380 565.020 210.390 ;
        RECT 742.020 210.380 745.020 210.390 ;
        RECT 922.020 210.380 925.020 210.390 ;
        RECT 1102.020 210.380 1105.020 210.390 ;
        RECT 1282.020 210.380 1285.020 210.390 ;
        RECT 1462.020 210.380 1465.020 210.390 ;
        RECT 1642.020 210.380 1645.020 210.390 ;
        RECT 1822.020 210.380 1825.020 210.390 ;
        RECT 2002.020 210.380 2005.020 210.390 ;
        RECT 2182.020 210.380 2185.020 210.390 ;
        RECT 2362.020 210.380 2365.020 210.390 ;
        RECT 2542.020 210.380 2545.020 210.390 ;
        RECT 2722.020 210.380 2725.020 210.390 ;
        RECT 2902.020 210.380 2905.020 210.390 ;
        RECT 2935.800 210.380 2938.800 210.390 ;
        RECT -23.780 207.380 2943.400 210.380 ;
        RECT -19.180 207.370 -16.180 207.380 ;
        RECT 22.020 207.370 25.020 207.380 ;
        RECT 202.020 207.370 205.020 207.380 ;
        RECT 382.020 207.370 385.020 207.380 ;
        RECT 562.020 207.370 565.020 207.380 ;
        RECT 742.020 207.370 745.020 207.380 ;
        RECT 922.020 207.370 925.020 207.380 ;
        RECT 1102.020 207.370 1105.020 207.380 ;
        RECT 1282.020 207.370 1285.020 207.380 ;
        RECT 1462.020 207.370 1465.020 207.380 ;
        RECT 1642.020 207.370 1645.020 207.380 ;
        RECT 1822.020 207.370 1825.020 207.380 ;
        RECT 2002.020 207.370 2005.020 207.380 ;
        RECT 2182.020 207.370 2185.020 207.380 ;
        RECT 2362.020 207.370 2365.020 207.380 ;
        RECT 2542.020 207.370 2545.020 207.380 ;
        RECT 2722.020 207.370 2725.020 207.380 ;
        RECT 2902.020 207.370 2905.020 207.380 ;
        RECT 2935.800 207.370 2938.800 207.380 ;
        RECT -19.180 30.380 -16.180 30.390 ;
        RECT 22.020 30.380 25.020 30.390 ;
        RECT 202.020 30.380 205.020 30.390 ;
        RECT 382.020 30.380 385.020 30.390 ;
        RECT 562.020 30.380 565.020 30.390 ;
        RECT 742.020 30.380 745.020 30.390 ;
        RECT 922.020 30.380 925.020 30.390 ;
        RECT 1102.020 30.380 1105.020 30.390 ;
        RECT 1282.020 30.380 1285.020 30.390 ;
        RECT 1462.020 30.380 1465.020 30.390 ;
        RECT 1642.020 30.380 1645.020 30.390 ;
        RECT 1822.020 30.380 1825.020 30.390 ;
        RECT 2002.020 30.380 2005.020 30.390 ;
        RECT 2182.020 30.380 2185.020 30.390 ;
        RECT 2362.020 30.380 2365.020 30.390 ;
        RECT 2542.020 30.380 2545.020 30.390 ;
        RECT 2722.020 30.380 2725.020 30.390 ;
        RECT 2902.020 30.380 2905.020 30.390 ;
        RECT 2935.800 30.380 2938.800 30.390 ;
        RECT -23.780 27.380 2943.400 30.380 ;
        RECT -19.180 27.370 -16.180 27.380 ;
        RECT 22.020 27.370 25.020 27.380 ;
        RECT 202.020 27.370 205.020 27.380 ;
        RECT 382.020 27.370 385.020 27.380 ;
        RECT 562.020 27.370 565.020 27.380 ;
        RECT 742.020 27.370 745.020 27.380 ;
        RECT 922.020 27.370 925.020 27.380 ;
        RECT 1102.020 27.370 1105.020 27.380 ;
        RECT 1282.020 27.370 1285.020 27.380 ;
        RECT 1462.020 27.370 1465.020 27.380 ;
        RECT 1642.020 27.370 1645.020 27.380 ;
        RECT 1822.020 27.370 1825.020 27.380 ;
        RECT 2002.020 27.370 2005.020 27.380 ;
        RECT 2182.020 27.370 2185.020 27.380 ;
        RECT 2362.020 27.370 2365.020 27.380 ;
        RECT 2542.020 27.370 2545.020 27.380 ;
        RECT 2722.020 27.370 2725.020 27.380 ;
        RECT 2902.020 27.370 2905.020 27.380 ;
        RECT 2935.800 27.370 2938.800 27.380 ;
        RECT -19.180 -10.820 -16.180 -10.810 ;
        RECT 22.020 -10.820 25.020 -10.810 ;
        RECT 202.020 -10.820 205.020 -10.810 ;
        RECT 382.020 -10.820 385.020 -10.810 ;
        RECT 562.020 -10.820 565.020 -10.810 ;
        RECT 742.020 -10.820 745.020 -10.810 ;
        RECT 922.020 -10.820 925.020 -10.810 ;
        RECT 1102.020 -10.820 1105.020 -10.810 ;
        RECT 1282.020 -10.820 1285.020 -10.810 ;
        RECT 1462.020 -10.820 1465.020 -10.810 ;
        RECT 1642.020 -10.820 1645.020 -10.810 ;
        RECT 1822.020 -10.820 1825.020 -10.810 ;
        RECT 2002.020 -10.820 2005.020 -10.810 ;
        RECT 2182.020 -10.820 2185.020 -10.810 ;
        RECT 2362.020 -10.820 2365.020 -10.810 ;
        RECT 2542.020 -10.820 2545.020 -10.810 ;
        RECT 2722.020 -10.820 2725.020 -10.810 ;
        RECT 2902.020 -10.820 2905.020 -10.810 ;
        RECT 2935.800 -10.820 2938.800 -10.810 ;
        RECT -19.180 -13.820 2938.800 -10.820 ;
        RECT -19.180 -13.830 -16.180 -13.820 ;
        RECT 22.020 -13.830 25.020 -13.820 ;
        RECT 202.020 -13.830 205.020 -13.820 ;
        RECT 382.020 -13.830 385.020 -13.820 ;
        RECT 562.020 -13.830 565.020 -13.820 ;
        RECT 742.020 -13.830 745.020 -13.820 ;
        RECT 922.020 -13.830 925.020 -13.820 ;
        RECT 1102.020 -13.830 1105.020 -13.820 ;
        RECT 1282.020 -13.830 1285.020 -13.820 ;
        RECT 1462.020 -13.830 1465.020 -13.820 ;
        RECT 1642.020 -13.830 1645.020 -13.820 ;
        RECT 1822.020 -13.830 1825.020 -13.820 ;
        RECT 2002.020 -13.830 2005.020 -13.820 ;
        RECT 2182.020 -13.830 2185.020 -13.820 ;
        RECT 2362.020 -13.830 2365.020 -13.820 ;
        RECT 2542.020 -13.830 2545.020 -13.820 ;
        RECT 2722.020 -13.830 2725.020 -13.820 ;
        RECT 2902.020 -13.830 2905.020 -13.820 ;
        RECT 2935.800 -13.830 2938.800 -13.820 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -23.780 -18.420 -20.780 3538.100 ;
        RECT 112.020 -18.420 115.020 3538.100 ;
        RECT 292.020 -18.420 295.020 3538.100 ;
        RECT 472.020 -18.420 475.020 3538.100 ;
        RECT 652.020 -18.420 655.020 3538.100 ;
        RECT 832.020 -18.420 835.020 3538.100 ;
        RECT 1012.020 -18.420 1015.020 3538.100 ;
        RECT 1192.020 -18.420 1195.020 3538.100 ;
        RECT 1372.020 -18.420 1375.020 3538.100 ;
        RECT 1552.020 -18.420 1555.020 3538.100 ;
        RECT 1732.020 -18.420 1735.020 3538.100 ;
        RECT 1912.020 -18.420 1915.020 3538.100 ;
        RECT 2092.020 -18.420 2095.020 3538.100 ;
        RECT 2272.020 -18.420 2275.020 3538.100 ;
        RECT 2452.020 -18.420 2455.020 3538.100 ;
        RECT 2632.020 -18.420 2635.020 3538.100 ;
        RECT 2812.020 -18.420 2815.020 3538.100 ;
        RECT 2940.400 -18.420 2943.400 3538.100 ;
      LAYER via4 ;
        RECT -22.870 3536.810 -21.690 3537.990 ;
        RECT -22.870 3535.210 -21.690 3536.390 ;
        RECT -22.870 3359.090 -21.690 3360.270 ;
        RECT -22.870 3357.490 -21.690 3358.670 ;
        RECT -22.870 3179.090 -21.690 3180.270 ;
        RECT -22.870 3177.490 -21.690 3178.670 ;
        RECT -22.870 2999.090 -21.690 3000.270 ;
        RECT -22.870 2997.490 -21.690 2998.670 ;
        RECT -22.870 2819.090 -21.690 2820.270 ;
        RECT -22.870 2817.490 -21.690 2818.670 ;
        RECT -22.870 2639.090 -21.690 2640.270 ;
        RECT -22.870 2637.490 -21.690 2638.670 ;
        RECT -22.870 2459.090 -21.690 2460.270 ;
        RECT -22.870 2457.490 -21.690 2458.670 ;
        RECT -22.870 2279.090 -21.690 2280.270 ;
        RECT -22.870 2277.490 -21.690 2278.670 ;
        RECT -22.870 2099.090 -21.690 2100.270 ;
        RECT -22.870 2097.490 -21.690 2098.670 ;
        RECT -22.870 1919.090 -21.690 1920.270 ;
        RECT -22.870 1917.490 -21.690 1918.670 ;
        RECT -22.870 1739.090 -21.690 1740.270 ;
        RECT -22.870 1737.490 -21.690 1738.670 ;
        RECT -22.870 1559.090 -21.690 1560.270 ;
        RECT -22.870 1557.490 -21.690 1558.670 ;
        RECT -22.870 1379.090 -21.690 1380.270 ;
        RECT -22.870 1377.490 -21.690 1378.670 ;
        RECT -22.870 1199.090 -21.690 1200.270 ;
        RECT -22.870 1197.490 -21.690 1198.670 ;
        RECT -22.870 1019.090 -21.690 1020.270 ;
        RECT -22.870 1017.490 -21.690 1018.670 ;
        RECT -22.870 839.090 -21.690 840.270 ;
        RECT -22.870 837.490 -21.690 838.670 ;
        RECT -22.870 659.090 -21.690 660.270 ;
        RECT -22.870 657.490 -21.690 658.670 ;
        RECT -22.870 479.090 -21.690 480.270 ;
        RECT -22.870 477.490 -21.690 478.670 ;
        RECT -22.870 299.090 -21.690 300.270 ;
        RECT -22.870 297.490 -21.690 298.670 ;
        RECT -22.870 119.090 -21.690 120.270 ;
        RECT -22.870 117.490 -21.690 118.670 ;
        RECT -22.870 -16.710 -21.690 -15.530 ;
        RECT -22.870 -18.310 -21.690 -17.130 ;
        RECT 112.930 3536.810 114.110 3537.990 ;
        RECT 112.930 3535.210 114.110 3536.390 ;
        RECT 112.930 3359.090 114.110 3360.270 ;
        RECT 112.930 3357.490 114.110 3358.670 ;
        RECT 112.930 3179.090 114.110 3180.270 ;
        RECT 112.930 3177.490 114.110 3178.670 ;
        RECT 112.930 2999.090 114.110 3000.270 ;
        RECT 112.930 2997.490 114.110 2998.670 ;
        RECT 112.930 2819.090 114.110 2820.270 ;
        RECT 112.930 2817.490 114.110 2818.670 ;
        RECT 112.930 2639.090 114.110 2640.270 ;
        RECT 112.930 2637.490 114.110 2638.670 ;
        RECT 112.930 2459.090 114.110 2460.270 ;
        RECT 112.930 2457.490 114.110 2458.670 ;
        RECT 112.930 2279.090 114.110 2280.270 ;
        RECT 112.930 2277.490 114.110 2278.670 ;
        RECT 112.930 2099.090 114.110 2100.270 ;
        RECT 112.930 2097.490 114.110 2098.670 ;
        RECT 112.930 1919.090 114.110 1920.270 ;
        RECT 112.930 1917.490 114.110 1918.670 ;
        RECT 112.930 1739.090 114.110 1740.270 ;
        RECT 112.930 1737.490 114.110 1738.670 ;
        RECT 112.930 1559.090 114.110 1560.270 ;
        RECT 112.930 1557.490 114.110 1558.670 ;
        RECT 112.930 1379.090 114.110 1380.270 ;
        RECT 112.930 1377.490 114.110 1378.670 ;
        RECT 112.930 1199.090 114.110 1200.270 ;
        RECT 112.930 1197.490 114.110 1198.670 ;
        RECT 112.930 1019.090 114.110 1020.270 ;
        RECT 112.930 1017.490 114.110 1018.670 ;
        RECT 112.930 839.090 114.110 840.270 ;
        RECT 112.930 837.490 114.110 838.670 ;
        RECT 112.930 659.090 114.110 660.270 ;
        RECT 112.930 657.490 114.110 658.670 ;
        RECT 112.930 479.090 114.110 480.270 ;
        RECT 112.930 477.490 114.110 478.670 ;
        RECT 112.930 299.090 114.110 300.270 ;
        RECT 112.930 297.490 114.110 298.670 ;
        RECT 112.930 119.090 114.110 120.270 ;
        RECT 112.930 117.490 114.110 118.670 ;
        RECT 112.930 -16.710 114.110 -15.530 ;
        RECT 112.930 -18.310 114.110 -17.130 ;
        RECT 292.930 3536.810 294.110 3537.990 ;
        RECT 292.930 3535.210 294.110 3536.390 ;
        RECT 292.930 3359.090 294.110 3360.270 ;
        RECT 292.930 3357.490 294.110 3358.670 ;
        RECT 292.930 3179.090 294.110 3180.270 ;
        RECT 292.930 3177.490 294.110 3178.670 ;
        RECT 292.930 2999.090 294.110 3000.270 ;
        RECT 292.930 2997.490 294.110 2998.670 ;
        RECT 292.930 2819.090 294.110 2820.270 ;
        RECT 292.930 2817.490 294.110 2818.670 ;
        RECT 292.930 2639.090 294.110 2640.270 ;
        RECT 292.930 2637.490 294.110 2638.670 ;
        RECT 292.930 2459.090 294.110 2460.270 ;
        RECT 292.930 2457.490 294.110 2458.670 ;
        RECT 292.930 2279.090 294.110 2280.270 ;
        RECT 292.930 2277.490 294.110 2278.670 ;
        RECT 292.930 2099.090 294.110 2100.270 ;
        RECT 292.930 2097.490 294.110 2098.670 ;
        RECT 292.930 1919.090 294.110 1920.270 ;
        RECT 292.930 1917.490 294.110 1918.670 ;
        RECT 292.930 1739.090 294.110 1740.270 ;
        RECT 292.930 1737.490 294.110 1738.670 ;
        RECT 292.930 1559.090 294.110 1560.270 ;
        RECT 292.930 1557.490 294.110 1558.670 ;
        RECT 292.930 1379.090 294.110 1380.270 ;
        RECT 292.930 1377.490 294.110 1378.670 ;
        RECT 292.930 1199.090 294.110 1200.270 ;
        RECT 292.930 1197.490 294.110 1198.670 ;
        RECT 292.930 1019.090 294.110 1020.270 ;
        RECT 292.930 1017.490 294.110 1018.670 ;
        RECT 292.930 839.090 294.110 840.270 ;
        RECT 292.930 837.490 294.110 838.670 ;
        RECT 292.930 659.090 294.110 660.270 ;
        RECT 292.930 657.490 294.110 658.670 ;
        RECT 292.930 479.090 294.110 480.270 ;
        RECT 292.930 477.490 294.110 478.670 ;
        RECT 292.930 299.090 294.110 300.270 ;
        RECT 292.930 297.490 294.110 298.670 ;
        RECT 292.930 119.090 294.110 120.270 ;
        RECT 292.930 117.490 294.110 118.670 ;
        RECT 292.930 -16.710 294.110 -15.530 ;
        RECT 292.930 -18.310 294.110 -17.130 ;
        RECT 472.930 3536.810 474.110 3537.990 ;
        RECT 472.930 3535.210 474.110 3536.390 ;
        RECT 472.930 3359.090 474.110 3360.270 ;
        RECT 472.930 3357.490 474.110 3358.670 ;
        RECT 472.930 3179.090 474.110 3180.270 ;
        RECT 472.930 3177.490 474.110 3178.670 ;
        RECT 472.930 2999.090 474.110 3000.270 ;
        RECT 472.930 2997.490 474.110 2998.670 ;
        RECT 472.930 2819.090 474.110 2820.270 ;
        RECT 472.930 2817.490 474.110 2818.670 ;
        RECT 472.930 2639.090 474.110 2640.270 ;
        RECT 472.930 2637.490 474.110 2638.670 ;
        RECT 472.930 2459.090 474.110 2460.270 ;
        RECT 472.930 2457.490 474.110 2458.670 ;
        RECT 472.930 2279.090 474.110 2280.270 ;
        RECT 472.930 2277.490 474.110 2278.670 ;
        RECT 472.930 2099.090 474.110 2100.270 ;
        RECT 472.930 2097.490 474.110 2098.670 ;
        RECT 472.930 1919.090 474.110 1920.270 ;
        RECT 472.930 1917.490 474.110 1918.670 ;
        RECT 472.930 1739.090 474.110 1740.270 ;
        RECT 472.930 1737.490 474.110 1738.670 ;
        RECT 472.930 1559.090 474.110 1560.270 ;
        RECT 472.930 1557.490 474.110 1558.670 ;
        RECT 472.930 1379.090 474.110 1380.270 ;
        RECT 472.930 1377.490 474.110 1378.670 ;
        RECT 472.930 1199.090 474.110 1200.270 ;
        RECT 472.930 1197.490 474.110 1198.670 ;
        RECT 472.930 1019.090 474.110 1020.270 ;
        RECT 472.930 1017.490 474.110 1018.670 ;
        RECT 472.930 839.090 474.110 840.270 ;
        RECT 472.930 837.490 474.110 838.670 ;
        RECT 472.930 659.090 474.110 660.270 ;
        RECT 472.930 657.490 474.110 658.670 ;
        RECT 472.930 479.090 474.110 480.270 ;
        RECT 472.930 477.490 474.110 478.670 ;
        RECT 472.930 299.090 474.110 300.270 ;
        RECT 472.930 297.490 474.110 298.670 ;
        RECT 472.930 119.090 474.110 120.270 ;
        RECT 472.930 117.490 474.110 118.670 ;
        RECT 472.930 -16.710 474.110 -15.530 ;
        RECT 472.930 -18.310 474.110 -17.130 ;
        RECT 652.930 3536.810 654.110 3537.990 ;
        RECT 652.930 3535.210 654.110 3536.390 ;
        RECT 652.930 3359.090 654.110 3360.270 ;
        RECT 652.930 3357.490 654.110 3358.670 ;
        RECT 652.930 3179.090 654.110 3180.270 ;
        RECT 652.930 3177.490 654.110 3178.670 ;
        RECT 652.930 2999.090 654.110 3000.270 ;
        RECT 652.930 2997.490 654.110 2998.670 ;
        RECT 652.930 2819.090 654.110 2820.270 ;
        RECT 652.930 2817.490 654.110 2818.670 ;
        RECT 652.930 2639.090 654.110 2640.270 ;
        RECT 652.930 2637.490 654.110 2638.670 ;
        RECT 652.930 2459.090 654.110 2460.270 ;
        RECT 652.930 2457.490 654.110 2458.670 ;
        RECT 652.930 2279.090 654.110 2280.270 ;
        RECT 652.930 2277.490 654.110 2278.670 ;
        RECT 652.930 2099.090 654.110 2100.270 ;
        RECT 652.930 2097.490 654.110 2098.670 ;
        RECT 652.930 1919.090 654.110 1920.270 ;
        RECT 652.930 1917.490 654.110 1918.670 ;
        RECT 652.930 1739.090 654.110 1740.270 ;
        RECT 652.930 1737.490 654.110 1738.670 ;
        RECT 652.930 1559.090 654.110 1560.270 ;
        RECT 652.930 1557.490 654.110 1558.670 ;
        RECT 652.930 1379.090 654.110 1380.270 ;
        RECT 652.930 1377.490 654.110 1378.670 ;
        RECT 652.930 1199.090 654.110 1200.270 ;
        RECT 652.930 1197.490 654.110 1198.670 ;
        RECT 652.930 1019.090 654.110 1020.270 ;
        RECT 652.930 1017.490 654.110 1018.670 ;
        RECT 652.930 839.090 654.110 840.270 ;
        RECT 652.930 837.490 654.110 838.670 ;
        RECT 652.930 659.090 654.110 660.270 ;
        RECT 652.930 657.490 654.110 658.670 ;
        RECT 652.930 479.090 654.110 480.270 ;
        RECT 652.930 477.490 654.110 478.670 ;
        RECT 652.930 299.090 654.110 300.270 ;
        RECT 652.930 297.490 654.110 298.670 ;
        RECT 652.930 119.090 654.110 120.270 ;
        RECT 652.930 117.490 654.110 118.670 ;
        RECT 652.930 -16.710 654.110 -15.530 ;
        RECT 652.930 -18.310 654.110 -17.130 ;
        RECT 832.930 3536.810 834.110 3537.990 ;
        RECT 832.930 3535.210 834.110 3536.390 ;
        RECT 832.930 3359.090 834.110 3360.270 ;
        RECT 832.930 3357.490 834.110 3358.670 ;
        RECT 832.930 3179.090 834.110 3180.270 ;
        RECT 832.930 3177.490 834.110 3178.670 ;
        RECT 832.930 2999.090 834.110 3000.270 ;
        RECT 832.930 2997.490 834.110 2998.670 ;
        RECT 832.930 2819.090 834.110 2820.270 ;
        RECT 832.930 2817.490 834.110 2818.670 ;
        RECT 832.930 2639.090 834.110 2640.270 ;
        RECT 832.930 2637.490 834.110 2638.670 ;
        RECT 832.930 2459.090 834.110 2460.270 ;
        RECT 832.930 2457.490 834.110 2458.670 ;
        RECT 832.930 2279.090 834.110 2280.270 ;
        RECT 832.930 2277.490 834.110 2278.670 ;
        RECT 832.930 2099.090 834.110 2100.270 ;
        RECT 832.930 2097.490 834.110 2098.670 ;
        RECT 832.930 1919.090 834.110 1920.270 ;
        RECT 832.930 1917.490 834.110 1918.670 ;
        RECT 832.930 1739.090 834.110 1740.270 ;
        RECT 832.930 1737.490 834.110 1738.670 ;
        RECT 832.930 1559.090 834.110 1560.270 ;
        RECT 832.930 1557.490 834.110 1558.670 ;
        RECT 832.930 1379.090 834.110 1380.270 ;
        RECT 832.930 1377.490 834.110 1378.670 ;
        RECT 832.930 1199.090 834.110 1200.270 ;
        RECT 832.930 1197.490 834.110 1198.670 ;
        RECT 832.930 1019.090 834.110 1020.270 ;
        RECT 832.930 1017.490 834.110 1018.670 ;
        RECT 832.930 839.090 834.110 840.270 ;
        RECT 832.930 837.490 834.110 838.670 ;
        RECT 832.930 659.090 834.110 660.270 ;
        RECT 832.930 657.490 834.110 658.670 ;
        RECT 832.930 479.090 834.110 480.270 ;
        RECT 832.930 477.490 834.110 478.670 ;
        RECT 832.930 299.090 834.110 300.270 ;
        RECT 832.930 297.490 834.110 298.670 ;
        RECT 832.930 119.090 834.110 120.270 ;
        RECT 832.930 117.490 834.110 118.670 ;
        RECT 832.930 -16.710 834.110 -15.530 ;
        RECT 832.930 -18.310 834.110 -17.130 ;
        RECT 1012.930 3536.810 1014.110 3537.990 ;
        RECT 1012.930 3535.210 1014.110 3536.390 ;
        RECT 1012.930 3359.090 1014.110 3360.270 ;
        RECT 1012.930 3357.490 1014.110 3358.670 ;
        RECT 1012.930 3179.090 1014.110 3180.270 ;
        RECT 1012.930 3177.490 1014.110 3178.670 ;
        RECT 1012.930 2999.090 1014.110 3000.270 ;
        RECT 1012.930 2997.490 1014.110 2998.670 ;
        RECT 1012.930 2819.090 1014.110 2820.270 ;
        RECT 1012.930 2817.490 1014.110 2818.670 ;
        RECT 1012.930 2639.090 1014.110 2640.270 ;
        RECT 1012.930 2637.490 1014.110 2638.670 ;
        RECT 1012.930 2459.090 1014.110 2460.270 ;
        RECT 1012.930 2457.490 1014.110 2458.670 ;
        RECT 1012.930 2279.090 1014.110 2280.270 ;
        RECT 1012.930 2277.490 1014.110 2278.670 ;
        RECT 1012.930 2099.090 1014.110 2100.270 ;
        RECT 1012.930 2097.490 1014.110 2098.670 ;
        RECT 1012.930 1919.090 1014.110 1920.270 ;
        RECT 1012.930 1917.490 1014.110 1918.670 ;
        RECT 1012.930 1739.090 1014.110 1740.270 ;
        RECT 1012.930 1737.490 1014.110 1738.670 ;
        RECT 1012.930 1559.090 1014.110 1560.270 ;
        RECT 1012.930 1557.490 1014.110 1558.670 ;
        RECT 1012.930 1379.090 1014.110 1380.270 ;
        RECT 1012.930 1377.490 1014.110 1378.670 ;
        RECT 1012.930 1199.090 1014.110 1200.270 ;
        RECT 1012.930 1197.490 1014.110 1198.670 ;
        RECT 1012.930 1019.090 1014.110 1020.270 ;
        RECT 1012.930 1017.490 1014.110 1018.670 ;
        RECT 1012.930 839.090 1014.110 840.270 ;
        RECT 1012.930 837.490 1014.110 838.670 ;
        RECT 1012.930 659.090 1014.110 660.270 ;
        RECT 1012.930 657.490 1014.110 658.670 ;
        RECT 1012.930 479.090 1014.110 480.270 ;
        RECT 1012.930 477.490 1014.110 478.670 ;
        RECT 1012.930 299.090 1014.110 300.270 ;
        RECT 1012.930 297.490 1014.110 298.670 ;
        RECT 1012.930 119.090 1014.110 120.270 ;
        RECT 1012.930 117.490 1014.110 118.670 ;
        RECT 1012.930 -16.710 1014.110 -15.530 ;
        RECT 1012.930 -18.310 1014.110 -17.130 ;
        RECT 1192.930 3536.810 1194.110 3537.990 ;
        RECT 1192.930 3535.210 1194.110 3536.390 ;
        RECT 1192.930 3359.090 1194.110 3360.270 ;
        RECT 1192.930 3357.490 1194.110 3358.670 ;
        RECT 1192.930 3179.090 1194.110 3180.270 ;
        RECT 1192.930 3177.490 1194.110 3178.670 ;
        RECT 1192.930 2999.090 1194.110 3000.270 ;
        RECT 1192.930 2997.490 1194.110 2998.670 ;
        RECT 1192.930 2819.090 1194.110 2820.270 ;
        RECT 1192.930 2817.490 1194.110 2818.670 ;
        RECT 1192.930 2639.090 1194.110 2640.270 ;
        RECT 1192.930 2637.490 1194.110 2638.670 ;
        RECT 1192.930 2459.090 1194.110 2460.270 ;
        RECT 1192.930 2457.490 1194.110 2458.670 ;
        RECT 1192.930 2279.090 1194.110 2280.270 ;
        RECT 1192.930 2277.490 1194.110 2278.670 ;
        RECT 1192.930 2099.090 1194.110 2100.270 ;
        RECT 1192.930 2097.490 1194.110 2098.670 ;
        RECT 1192.930 1919.090 1194.110 1920.270 ;
        RECT 1192.930 1917.490 1194.110 1918.670 ;
        RECT 1192.930 1739.090 1194.110 1740.270 ;
        RECT 1192.930 1737.490 1194.110 1738.670 ;
        RECT 1192.930 1559.090 1194.110 1560.270 ;
        RECT 1192.930 1557.490 1194.110 1558.670 ;
        RECT 1192.930 1379.090 1194.110 1380.270 ;
        RECT 1192.930 1377.490 1194.110 1378.670 ;
        RECT 1192.930 1199.090 1194.110 1200.270 ;
        RECT 1192.930 1197.490 1194.110 1198.670 ;
        RECT 1192.930 1019.090 1194.110 1020.270 ;
        RECT 1192.930 1017.490 1194.110 1018.670 ;
        RECT 1192.930 839.090 1194.110 840.270 ;
        RECT 1192.930 837.490 1194.110 838.670 ;
        RECT 1192.930 659.090 1194.110 660.270 ;
        RECT 1192.930 657.490 1194.110 658.670 ;
        RECT 1192.930 479.090 1194.110 480.270 ;
        RECT 1192.930 477.490 1194.110 478.670 ;
        RECT 1192.930 299.090 1194.110 300.270 ;
        RECT 1192.930 297.490 1194.110 298.670 ;
        RECT 1192.930 119.090 1194.110 120.270 ;
        RECT 1192.930 117.490 1194.110 118.670 ;
        RECT 1192.930 -16.710 1194.110 -15.530 ;
        RECT 1192.930 -18.310 1194.110 -17.130 ;
        RECT 1372.930 3536.810 1374.110 3537.990 ;
        RECT 1372.930 3535.210 1374.110 3536.390 ;
        RECT 1372.930 3359.090 1374.110 3360.270 ;
        RECT 1372.930 3357.490 1374.110 3358.670 ;
        RECT 1372.930 3179.090 1374.110 3180.270 ;
        RECT 1372.930 3177.490 1374.110 3178.670 ;
        RECT 1372.930 2999.090 1374.110 3000.270 ;
        RECT 1372.930 2997.490 1374.110 2998.670 ;
        RECT 1372.930 2819.090 1374.110 2820.270 ;
        RECT 1372.930 2817.490 1374.110 2818.670 ;
        RECT 1372.930 2639.090 1374.110 2640.270 ;
        RECT 1372.930 2637.490 1374.110 2638.670 ;
        RECT 1372.930 2459.090 1374.110 2460.270 ;
        RECT 1372.930 2457.490 1374.110 2458.670 ;
        RECT 1372.930 2279.090 1374.110 2280.270 ;
        RECT 1372.930 2277.490 1374.110 2278.670 ;
        RECT 1372.930 2099.090 1374.110 2100.270 ;
        RECT 1372.930 2097.490 1374.110 2098.670 ;
        RECT 1372.930 1919.090 1374.110 1920.270 ;
        RECT 1372.930 1917.490 1374.110 1918.670 ;
        RECT 1372.930 1739.090 1374.110 1740.270 ;
        RECT 1372.930 1737.490 1374.110 1738.670 ;
        RECT 1372.930 1559.090 1374.110 1560.270 ;
        RECT 1372.930 1557.490 1374.110 1558.670 ;
        RECT 1372.930 1379.090 1374.110 1380.270 ;
        RECT 1372.930 1377.490 1374.110 1378.670 ;
        RECT 1372.930 1199.090 1374.110 1200.270 ;
        RECT 1372.930 1197.490 1374.110 1198.670 ;
        RECT 1372.930 1019.090 1374.110 1020.270 ;
        RECT 1372.930 1017.490 1374.110 1018.670 ;
        RECT 1372.930 839.090 1374.110 840.270 ;
        RECT 1372.930 837.490 1374.110 838.670 ;
        RECT 1372.930 659.090 1374.110 660.270 ;
        RECT 1372.930 657.490 1374.110 658.670 ;
        RECT 1372.930 479.090 1374.110 480.270 ;
        RECT 1372.930 477.490 1374.110 478.670 ;
        RECT 1372.930 299.090 1374.110 300.270 ;
        RECT 1372.930 297.490 1374.110 298.670 ;
        RECT 1372.930 119.090 1374.110 120.270 ;
        RECT 1372.930 117.490 1374.110 118.670 ;
        RECT 1372.930 -16.710 1374.110 -15.530 ;
        RECT 1372.930 -18.310 1374.110 -17.130 ;
        RECT 1552.930 3536.810 1554.110 3537.990 ;
        RECT 1552.930 3535.210 1554.110 3536.390 ;
        RECT 1552.930 3359.090 1554.110 3360.270 ;
        RECT 1552.930 3357.490 1554.110 3358.670 ;
        RECT 1552.930 3179.090 1554.110 3180.270 ;
        RECT 1552.930 3177.490 1554.110 3178.670 ;
        RECT 1552.930 2999.090 1554.110 3000.270 ;
        RECT 1552.930 2997.490 1554.110 2998.670 ;
        RECT 1552.930 2819.090 1554.110 2820.270 ;
        RECT 1552.930 2817.490 1554.110 2818.670 ;
        RECT 1552.930 2639.090 1554.110 2640.270 ;
        RECT 1552.930 2637.490 1554.110 2638.670 ;
        RECT 1552.930 2459.090 1554.110 2460.270 ;
        RECT 1552.930 2457.490 1554.110 2458.670 ;
        RECT 1552.930 2279.090 1554.110 2280.270 ;
        RECT 1552.930 2277.490 1554.110 2278.670 ;
        RECT 1552.930 2099.090 1554.110 2100.270 ;
        RECT 1552.930 2097.490 1554.110 2098.670 ;
        RECT 1552.930 1919.090 1554.110 1920.270 ;
        RECT 1552.930 1917.490 1554.110 1918.670 ;
        RECT 1552.930 1739.090 1554.110 1740.270 ;
        RECT 1552.930 1737.490 1554.110 1738.670 ;
        RECT 1552.930 1559.090 1554.110 1560.270 ;
        RECT 1552.930 1557.490 1554.110 1558.670 ;
        RECT 1552.930 1379.090 1554.110 1380.270 ;
        RECT 1552.930 1377.490 1554.110 1378.670 ;
        RECT 1552.930 1199.090 1554.110 1200.270 ;
        RECT 1552.930 1197.490 1554.110 1198.670 ;
        RECT 1552.930 1019.090 1554.110 1020.270 ;
        RECT 1552.930 1017.490 1554.110 1018.670 ;
        RECT 1552.930 839.090 1554.110 840.270 ;
        RECT 1552.930 837.490 1554.110 838.670 ;
        RECT 1552.930 659.090 1554.110 660.270 ;
        RECT 1552.930 657.490 1554.110 658.670 ;
        RECT 1552.930 479.090 1554.110 480.270 ;
        RECT 1552.930 477.490 1554.110 478.670 ;
        RECT 1552.930 299.090 1554.110 300.270 ;
        RECT 1552.930 297.490 1554.110 298.670 ;
        RECT 1552.930 119.090 1554.110 120.270 ;
        RECT 1552.930 117.490 1554.110 118.670 ;
        RECT 1552.930 -16.710 1554.110 -15.530 ;
        RECT 1552.930 -18.310 1554.110 -17.130 ;
        RECT 1732.930 3536.810 1734.110 3537.990 ;
        RECT 1732.930 3535.210 1734.110 3536.390 ;
        RECT 1732.930 3359.090 1734.110 3360.270 ;
        RECT 1732.930 3357.490 1734.110 3358.670 ;
        RECT 1732.930 3179.090 1734.110 3180.270 ;
        RECT 1732.930 3177.490 1734.110 3178.670 ;
        RECT 1732.930 2999.090 1734.110 3000.270 ;
        RECT 1732.930 2997.490 1734.110 2998.670 ;
        RECT 1732.930 2819.090 1734.110 2820.270 ;
        RECT 1732.930 2817.490 1734.110 2818.670 ;
        RECT 1732.930 2639.090 1734.110 2640.270 ;
        RECT 1732.930 2637.490 1734.110 2638.670 ;
        RECT 1732.930 2459.090 1734.110 2460.270 ;
        RECT 1732.930 2457.490 1734.110 2458.670 ;
        RECT 1732.930 2279.090 1734.110 2280.270 ;
        RECT 1732.930 2277.490 1734.110 2278.670 ;
        RECT 1732.930 2099.090 1734.110 2100.270 ;
        RECT 1732.930 2097.490 1734.110 2098.670 ;
        RECT 1732.930 1919.090 1734.110 1920.270 ;
        RECT 1732.930 1917.490 1734.110 1918.670 ;
        RECT 1732.930 1739.090 1734.110 1740.270 ;
        RECT 1732.930 1737.490 1734.110 1738.670 ;
        RECT 1732.930 1559.090 1734.110 1560.270 ;
        RECT 1732.930 1557.490 1734.110 1558.670 ;
        RECT 1732.930 1379.090 1734.110 1380.270 ;
        RECT 1732.930 1377.490 1734.110 1378.670 ;
        RECT 1732.930 1199.090 1734.110 1200.270 ;
        RECT 1732.930 1197.490 1734.110 1198.670 ;
        RECT 1732.930 1019.090 1734.110 1020.270 ;
        RECT 1732.930 1017.490 1734.110 1018.670 ;
        RECT 1732.930 839.090 1734.110 840.270 ;
        RECT 1732.930 837.490 1734.110 838.670 ;
        RECT 1732.930 659.090 1734.110 660.270 ;
        RECT 1732.930 657.490 1734.110 658.670 ;
        RECT 1732.930 479.090 1734.110 480.270 ;
        RECT 1732.930 477.490 1734.110 478.670 ;
        RECT 1732.930 299.090 1734.110 300.270 ;
        RECT 1732.930 297.490 1734.110 298.670 ;
        RECT 1732.930 119.090 1734.110 120.270 ;
        RECT 1732.930 117.490 1734.110 118.670 ;
        RECT 1732.930 -16.710 1734.110 -15.530 ;
        RECT 1732.930 -18.310 1734.110 -17.130 ;
        RECT 1912.930 3536.810 1914.110 3537.990 ;
        RECT 1912.930 3535.210 1914.110 3536.390 ;
        RECT 1912.930 3359.090 1914.110 3360.270 ;
        RECT 1912.930 3357.490 1914.110 3358.670 ;
        RECT 1912.930 3179.090 1914.110 3180.270 ;
        RECT 1912.930 3177.490 1914.110 3178.670 ;
        RECT 1912.930 2999.090 1914.110 3000.270 ;
        RECT 1912.930 2997.490 1914.110 2998.670 ;
        RECT 1912.930 2819.090 1914.110 2820.270 ;
        RECT 1912.930 2817.490 1914.110 2818.670 ;
        RECT 1912.930 2639.090 1914.110 2640.270 ;
        RECT 1912.930 2637.490 1914.110 2638.670 ;
        RECT 1912.930 2459.090 1914.110 2460.270 ;
        RECT 1912.930 2457.490 1914.110 2458.670 ;
        RECT 1912.930 2279.090 1914.110 2280.270 ;
        RECT 1912.930 2277.490 1914.110 2278.670 ;
        RECT 1912.930 2099.090 1914.110 2100.270 ;
        RECT 1912.930 2097.490 1914.110 2098.670 ;
        RECT 1912.930 1919.090 1914.110 1920.270 ;
        RECT 1912.930 1917.490 1914.110 1918.670 ;
        RECT 1912.930 1739.090 1914.110 1740.270 ;
        RECT 1912.930 1737.490 1914.110 1738.670 ;
        RECT 1912.930 1559.090 1914.110 1560.270 ;
        RECT 1912.930 1557.490 1914.110 1558.670 ;
        RECT 1912.930 1379.090 1914.110 1380.270 ;
        RECT 1912.930 1377.490 1914.110 1378.670 ;
        RECT 1912.930 1199.090 1914.110 1200.270 ;
        RECT 1912.930 1197.490 1914.110 1198.670 ;
        RECT 1912.930 1019.090 1914.110 1020.270 ;
        RECT 1912.930 1017.490 1914.110 1018.670 ;
        RECT 1912.930 839.090 1914.110 840.270 ;
        RECT 1912.930 837.490 1914.110 838.670 ;
        RECT 1912.930 659.090 1914.110 660.270 ;
        RECT 1912.930 657.490 1914.110 658.670 ;
        RECT 1912.930 479.090 1914.110 480.270 ;
        RECT 1912.930 477.490 1914.110 478.670 ;
        RECT 1912.930 299.090 1914.110 300.270 ;
        RECT 1912.930 297.490 1914.110 298.670 ;
        RECT 1912.930 119.090 1914.110 120.270 ;
        RECT 1912.930 117.490 1914.110 118.670 ;
        RECT 1912.930 -16.710 1914.110 -15.530 ;
        RECT 1912.930 -18.310 1914.110 -17.130 ;
        RECT 2092.930 3536.810 2094.110 3537.990 ;
        RECT 2092.930 3535.210 2094.110 3536.390 ;
        RECT 2092.930 3359.090 2094.110 3360.270 ;
        RECT 2092.930 3357.490 2094.110 3358.670 ;
        RECT 2092.930 3179.090 2094.110 3180.270 ;
        RECT 2092.930 3177.490 2094.110 3178.670 ;
        RECT 2092.930 2999.090 2094.110 3000.270 ;
        RECT 2092.930 2997.490 2094.110 2998.670 ;
        RECT 2092.930 2819.090 2094.110 2820.270 ;
        RECT 2092.930 2817.490 2094.110 2818.670 ;
        RECT 2092.930 2639.090 2094.110 2640.270 ;
        RECT 2092.930 2637.490 2094.110 2638.670 ;
        RECT 2092.930 2459.090 2094.110 2460.270 ;
        RECT 2092.930 2457.490 2094.110 2458.670 ;
        RECT 2092.930 2279.090 2094.110 2280.270 ;
        RECT 2092.930 2277.490 2094.110 2278.670 ;
        RECT 2092.930 2099.090 2094.110 2100.270 ;
        RECT 2092.930 2097.490 2094.110 2098.670 ;
        RECT 2092.930 1919.090 2094.110 1920.270 ;
        RECT 2092.930 1917.490 2094.110 1918.670 ;
        RECT 2092.930 1739.090 2094.110 1740.270 ;
        RECT 2092.930 1737.490 2094.110 1738.670 ;
        RECT 2092.930 1559.090 2094.110 1560.270 ;
        RECT 2092.930 1557.490 2094.110 1558.670 ;
        RECT 2092.930 1379.090 2094.110 1380.270 ;
        RECT 2092.930 1377.490 2094.110 1378.670 ;
        RECT 2092.930 1199.090 2094.110 1200.270 ;
        RECT 2092.930 1197.490 2094.110 1198.670 ;
        RECT 2092.930 1019.090 2094.110 1020.270 ;
        RECT 2092.930 1017.490 2094.110 1018.670 ;
        RECT 2092.930 839.090 2094.110 840.270 ;
        RECT 2092.930 837.490 2094.110 838.670 ;
        RECT 2092.930 659.090 2094.110 660.270 ;
        RECT 2092.930 657.490 2094.110 658.670 ;
        RECT 2092.930 479.090 2094.110 480.270 ;
        RECT 2092.930 477.490 2094.110 478.670 ;
        RECT 2092.930 299.090 2094.110 300.270 ;
        RECT 2092.930 297.490 2094.110 298.670 ;
        RECT 2092.930 119.090 2094.110 120.270 ;
        RECT 2092.930 117.490 2094.110 118.670 ;
        RECT 2092.930 -16.710 2094.110 -15.530 ;
        RECT 2092.930 -18.310 2094.110 -17.130 ;
        RECT 2272.930 3536.810 2274.110 3537.990 ;
        RECT 2272.930 3535.210 2274.110 3536.390 ;
        RECT 2272.930 3359.090 2274.110 3360.270 ;
        RECT 2272.930 3357.490 2274.110 3358.670 ;
        RECT 2272.930 3179.090 2274.110 3180.270 ;
        RECT 2272.930 3177.490 2274.110 3178.670 ;
        RECT 2272.930 2999.090 2274.110 3000.270 ;
        RECT 2272.930 2997.490 2274.110 2998.670 ;
        RECT 2272.930 2819.090 2274.110 2820.270 ;
        RECT 2272.930 2817.490 2274.110 2818.670 ;
        RECT 2272.930 2639.090 2274.110 2640.270 ;
        RECT 2272.930 2637.490 2274.110 2638.670 ;
        RECT 2272.930 2459.090 2274.110 2460.270 ;
        RECT 2272.930 2457.490 2274.110 2458.670 ;
        RECT 2272.930 2279.090 2274.110 2280.270 ;
        RECT 2272.930 2277.490 2274.110 2278.670 ;
        RECT 2272.930 2099.090 2274.110 2100.270 ;
        RECT 2272.930 2097.490 2274.110 2098.670 ;
        RECT 2272.930 1919.090 2274.110 1920.270 ;
        RECT 2272.930 1917.490 2274.110 1918.670 ;
        RECT 2272.930 1739.090 2274.110 1740.270 ;
        RECT 2272.930 1737.490 2274.110 1738.670 ;
        RECT 2272.930 1559.090 2274.110 1560.270 ;
        RECT 2272.930 1557.490 2274.110 1558.670 ;
        RECT 2272.930 1379.090 2274.110 1380.270 ;
        RECT 2272.930 1377.490 2274.110 1378.670 ;
        RECT 2272.930 1199.090 2274.110 1200.270 ;
        RECT 2272.930 1197.490 2274.110 1198.670 ;
        RECT 2272.930 1019.090 2274.110 1020.270 ;
        RECT 2272.930 1017.490 2274.110 1018.670 ;
        RECT 2272.930 839.090 2274.110 840.270 ;
        RECT 2272.930 837.490 2274.110 838.670 ;
        RECT 2272.930 659.090 2274.110 660.270 ;
        RECT 2272.930 657.490 2274.110 658.670 ;
        RECT 2272.930 479.090 2274.110 480.270 ;
        RECT 2272.930 477.490 2274.110 478.670 ;
        RECT 2272.930 299.090 2274.110 300.270 ;
        RECT 2272.930 297.490 2274.110 298.670 ;
        RECT 2272.930 119.090 2274.110 120.270 ;
        RECT 2272.930 117.490 2274.110 118.670 ;
        RECT 2272.930 -16.710 2274.110 -15.530 ;
        RECT 2272.930 -18.310 2274.110 -17.130 ;
        RECT 2452.930 3536.810 2454.110 3537.990 ;
        RECT 2452.930 3535.210 2454.110 3536.390 ;
        RECT 2452.930 3359.090 2454.110 3360.270 ;
        RECT 2452.930 3357.490 2454.110 3358.670 ;
        RECT 2452.930 3179.090 2454.110 3180.270 ;
        RECT 2452.930 3177.490 2454.110 3178.670 ;
        RECT 2452.930 2999.090 2454.110 3000.270 ;
        RECT 2452.930 2997.490 2454.110 2998.670 ;
        RECT 2452.930 2819.090 2454.110 2820.270 ;
        RECT 2452.930 2817.490 2454.110 2818.670 ;
        RECT 2452.930 2639.090 2454.110 2640.270 ;
        RECT 2452.930 2637.490 2454.110 2638.670 ;
        RECT 2452.930 2459.090 2454.110 2460.270 ;
        RECT 2452.930 2457.490 2454.110 2458.670 ;
        RECT 2452.930 2279.090 2454.110 2280.270 ;
        RECT 2452.930 2277.490 2454.110 2278.670 ;
        RECT 2452.930 2099.090 2454.110 2100.270 ;
        RECT 2452.930 2097.490 2454.110 2098.670 ;
        RECT 2452.930 1919.090 2454.110 1920.270 ;
        RECT 2452.930 1917.490 2454.110 1918.670 ;
        RECT 2452.930 1739.090 2454.110 1740.270 ;
        RECT 2452.930 1737.490 2454.110 1738.670 ;
        RECT 2452.930 1559.090 2454.110 1560.270 ;
        RECT 2452.930 1557.490 2454.110 1558.670 ;
        RECT 2452.930 1379.090 2454.110 1380.270 ;
        RECT 2452.930 1377.490 2454.110 1378.670 ;
        RECT 2452.930 1199.090 2454.110 1200.270 ;
        RECT 2452.930 1197.490 2454.110 1198.670 ;
        RECT 2452.930 1019.090 2454.110 1020.270 ;
        RECT 2452.930 1017.490 2454.110 1018.670 ;
        RECT 2452.930 839.090 2454.110 840.270 ;
        RECT 2452.930 837.490 2454.110 838.670 ;
        RECT 2452.930 659.090 2454.110 660.270 ;
        RECT 2452.930 657.490 2454.110 658.670 ;
        RECT 2452.930 479.090 2454.110 480.270 ;
        RECT 2452.930 477.490 2454.110 478.670 ;
        RECT 2452.930 299.090 2454.110 300.270 ;
        RECT 2452.930 297.490 2454.110 298.670 ;
        RECT 2452.930 119.090 2454.110 120.270 ;
        RECT 2452.930 117.490 2454.110 118.670 ;
        RECT 2452.930 -16.710 2454.110 -15.530 ;
        RECT 2452.930 -18.310 2454.110 -17.130 ;
        RECT 2632.930 3536.810 2634.110 3537.990 ;
        RECT 2632.930 3535.210 2634.110 3536.390 ;
        RECT 2632.930 3359.090 2634.110 3360.270 ;
        RECT 2632.930 3357.490 2634.110 3358.670 ;
        RECT 2632.930 3179.090 2634.110 3180.270 ;
        RECT 2632.930 3177.490 2634.110 3178.670 ;
        RECT 2632.930 2999.090 2634.110 3000.270 ;
        RECT 2632.930 2997.490 2634.110 2998.670 ;
        RECT 2632.930 2819.090 2634.110 2820.270 ;
        RECT 2632.930 2817.490 2634.110 2818.670 ;
        RECT 2632.930 2639.090 2634.110 2640.270 ;
        RECT 2632.930 2637.490 2634.110 2638.670 ;
        RECT 2632.930 2459.090 2634.110 2460.270 ;
        RECT 2632.930 2457.490 2634.110 2458.670 ;
        RECT 2632.930 2279.090 2634.110 2280.270 ;
        RECT 2632.930 2277.490 2634.110 2278.670 ;
        RECT 2632.930 2099.090 2634.110 2100.270 ;
        RECT 2632.930 2097.490 2634.110 2098.670 ;
        RECT 2632.930 1919.090 2634.110 1920.270 ;
        RECT 2632.930 1917.490 2634.110 1918.670 ;
        RECT 2632.930 1739.090 2634.110 1740.270 ;
        RECT 2632.930 1737.490 2634.110 1738.670 ;
        RECT 2632.930 1559.090 2634.110 1560.270 ;
        RECT 2632.930 1557.490 2634.110 1558.670 ;
        RECT 2632.930 1379.090 2634.110 1380.270 ;
        RECT 2632.930 1377.490 2634.110 1378.670 ;
        RECT 2632.930 1199.090 2634.110 1200.270 ;
        RECT 2632.930 1197.490 2634.110 1198.670 ;
        RECT 2632.930 1019.090 2634.110 1020.270 ;
        RECT 2632.930 1017.490 2634.110 1018.670 ;
        RECT 2632.930 839.090 2634.110 840.270 ;
        RECT 2632.930 837.490 2634.110 838.670 ;
        RECT 2632.930 659.090 2634.110 660.270 ;
        RECT 2632.930 657.490 2634.110 658.670 ;
        RECT 2632.930 479.090 2634.110 480.270 ;
        RECT 2632.930 477.490 2634.110 478.670 ;
        RECT 2632.930 299.090 2634.110 300.270 ;
        RECT 2632.930 297.490 2634.110 298.670 ;
        RECT 2632.930 119.090 2634.110 120.270 ;
        RECT 2632.930 117.490 2634.110 118.670 ;
        RECT 2632.930 -16.710 2634.110 -15.530 ;
        RECT 2632.930 -18.310 2634.110 -17.130 ;
        RECT 2812.930 3536.810 2814.110 3537.990 ;
        RECT 2812.930 3535.210 2814.110 3536.390 ;
        RECT 2812.930 3359.090 2814.110 3360.270 ;
        RECT 2812.930 3357.490 2814.110 3358.670 ;
        RECT 2812.930 3179.090 2814.110 3180.270 ;
        RECT 2812.930 3177.490 2814.110 3178.670 ;
        RECT 2812.930 2999.090 2814.110 3000.270 ;
        RECT 2812.930 2997.490 2814.110 2998.670 ;
        RECT 2812.930 2819.090 2814.110 2820.270 ;
        RECT 2812.930 2817.490 2814.110 2818.670 ;
        RECT 2812.930 2639.090 2814.110 2640.270 ;
        RECT 2812.930 2637.490 2814.110 2638.670 ;
        RECT 2812.930 2459.090 2814.110 2460.270 ;
        RECT 2812.930 2457.490 2814.110 2458.670 ;
        RECT 2812.930 2279.090 2814.110 2280.270 ;
        RECT 2812.930 2277.490 2814.110 2278.670 ;
        RECT 2812.930 2099.090 2814.110 2100.270 ;
        RECT 2812.930 2097.490 2814.110 2098.670 ;
        RECT 2812.930 1919.090 2814.110 1920.270 ;
        RECT 2812.930 1917.490 2814.110 1918.670 ;
        RECT 2812.930 1739.090 2814.110 1740.270 ;
        RECT 2812.930 1737.490 2814.110 1738.670 ;
        RECT 2812.930 1559.090 2814.110 1560.270 ;
        RECT 2812.930 1557.490 2814.110 1558.670 ;
        RECT 2812.930 1379.090 2814.110 1380.270 ;
        RECT 2812.930 1377.490 2814.110 1378.670 ;
        RECT 2812.930 1199.090 2814.110 1200.270 ;
        RECT 2812.930 1197.490 2814.110 1198.670 ;
        RECT 2812.930 1019.090 2814.110 1020.270 ;
        RECT 2812.930 1017.490 2814.110 1018.670 ;
        RECT 2812.930 839.090 2814.110 840.270 ;
        RECT 2812.930 837.490 2814.110 838.670 ;
        RECT 2812.930 659.090 2814.110 660.270 ;
        RECT 2812.930 657.490 2814.110 658.670 ;
        RECT 2812.930 479.090 2814.110 480.270 ;
        RECT 2812.930 477.490 2814.110 478.670 ;
        RECT 2812.930 299.090 2814.110 300.270 ;
        RECT 2812.930 297.490 2814.110 298.670 ;
        RECT 2812.930 119.090 2814.110 120.270 ;
        RECT 2812.930 117.490 2814.110 118.670 ;
        RECT 2812.930 -16.710 2814.110 -15.530 ;
        RECT 2812.930 -18.310 2814.110 -17.130 ;
        RECT 2941.310 3536.810 2942.490 3537.990 ;
        RECT 2941.310 3535.210 2942.490 3536.390 ;
        RECT 2941.310 3359.090 2942.490 3360.270 ;
        RECT 2941.310 3357.490 2942.490 3358.670 ;
        RECT 2941.310 3179.090 2942.490 3180.270 ;
        RECT 2941.310 3177.490 2942.490 3178.670 ;
        RECT 2941.310 2999.090 2942.490 3000.270 ;
        RECT 2941.310 2997.490 2942.490 2998.670 ;
        RECT 2941.310 2819.090 2942.490 2820.270 ;
        RECT 2941.310 2817.490 2942.490 2818.670 ;
        RECT 2941.310 2639.090 2942.490 2640.270 ;
        RECT 2941.310 2637.490 2942.490 2638.670 ;
        RECT 2941.310 2459.090 2942.490 2460.270 ;
        RECT 2941.310 2457.490 2942.490 2458.670 ;
        RECT 2941.310 2279.090 2942.490 2280.270 ;
        RECT 2941.310 2277.490 2942.490 2278.670 ;
        RECT 2941.310 2099.090 2942.490 2100.270 ;
        RECT 2941.310 2097.490 2942.490 2098.670 ;
        RECT 2941.310 1919.090 2942.490 1920.270 ;
        RECT 2941.310 1917.490 2942.490 1918.670 ;
        RECT 2941.310 1739.090 2942.490 1740.270 ;
        RECT 2941.310 1737.490 2942.490 1738.670 ;
        RECT 2941.310 1559.090 2942.490 1560.270 ;
        RECT 2941.310 1557.490 2942.490 1558.670 ;
        RECT 2941.310 1379.090 2942.490 1380.270 ;
        RECT 2941.310 1377.490 2942.490 1378.670 ;
        RECT 2941.310 1199.090 2942.490 1200.270 ;
        RECT 2941.310 1197.490 2942.490 1198.670 ;
        RECT 2941.310 1019.090 2942.490 1020.270 ;
        RECT 2941.310 1017.490 2942.490 1018.670 ;
        RECT 2941.310 839.090 2942.490 840.270 ;
        RECT 2941.310 837.490 2942.490 838.670 ;
        RECT 2941.310 659.090 2942.490 660.270 ;
        RECT 2941.310 657.490 2942.490 658.670 ;
        RECT 2941.310 479.090 2942.490 480.270 ;
        RECT 2941.310 477.490 2942.490 478.670 ;
        RECT 2941.310 299.090 2942.490 300.270 ;
        RECT 2941.310 297.490 2942.490 298.670 ;
        RECT 2941.310 119.090 2942.490 120.270 ;
        RECT 2941.310 117.490 2942.490 118.670 ;
        RECT 2941.310 -16.710 2942.490 -15.530 ;
        RECT 2941.310 -18.310 2942.490 -17.130 ;
      LAYER met5 ;
        RECT -23.780 3538.100 -20.780 3538.110 ;
        RECT 112.020 3538.100 115.020 3538.110 ;
        RECT 292.020 3538.100 295.020 3538.110 ;
        RECT 472.020 3538.100 475.020 3538.110 ;
        RECT 652.020 3538.100 655.020 3538.110 ;
        RECT 832.020 3538.100 835.020 3538.110 ;
        RECT 1012.020 3538.100 1015.020 3538.110 ;
        RECT 1192.020 3538.100 1195.020 3538.110 ;
        RECT 1372.020 3538.100 1375.020 3538.110 ;
        RECT 1552.020 3538.100 1555.020 3538.110 ;
        RECT 1732.020 3538.100 1735.020 3538.110 ;
        RECT 1912.020 3538.100 1915.020 3538.110 ;
        RECT 2092.020 3538.100 2095.020 3538.110 ;
        RECT 2272.020 3538.100 2275.020 3538.110 ;
        RECT 2452.020 3538.100 2455.020 3538.110 ;
        RECT 2632.020 3538.100 2635.020 3538.110 ;
        RECT 2812.020 3538.100 2815.020 3538.110 ;
        RECT 2940.400 3538.100 2943.400 3538.110 ;
        RECT -23.780 3535.100 2943.400 3538.100 ;
        RECT -23.780 3535.090 -20.780 3535.100 ;
        RECT 112.020 3535.090 115.020 3535.100 ;
        RECT 292.020 3535.090 295.020 3535.100 ;
        RECT 472.020 3535.090 475.020 3535.100 ;
        RECT 652.020 3535.090 655.020 3535.100 ;
        RECT 832.020 3535.090 835.020 3535.100 ;
        RECT 1012.020 3535.090 1015.020 3535.100 ;
        RECT 1192.020 3535.090 1195.020 3535.100 ;
        RECT 1372.020 3535.090 1375.020 3535.100 ;
        RECT 1552.020 3535.090 1555.020 3535.100 ;
        RECT 1732.020 3535.090 1735.020 3535.100 ;
        RECT 1912.020 3535.090 1915.020 3535.100 ;
        RECT 2092.020 3535.090 2095.020 3535.100 ;
        RECT 2272.020 3535.090 2275.020 3535.100 ;
        RECT 2452.020 3535.090 2455.020 3535.100 ;
        RECT 2632.020 3535.090 2635.020 3535.100 ;
        RECT 2812.020 3535.090 2815.020 3535.100 ;
        RECT 2940.400 3535.090 2943.400 3535.100 ;
        RECT -23.780 3360.380 -20.780 3360.390 ;
        RECT 112.020 3360.380 115.020 3360.390 ;
        RECT 292.020 3360.380 295.020 3360.390 ;
        RECT 472.020 3360.380 475.020 3360.390 ;
        RECT 652.020 3360.380 655.020 3360.390 ;
        RECT 832.020 3360.380 835.020 3360.390 ;
        RECT 1012.020 3360.380 1015.020 3360.390 ;
        RECT 1192.020 3360.380 1195.020 3360.390 ;
        RECT 1372.020 3360.380 1375.020 3360.390 ;
        RECT 1552.020 3360.380 1555.020 3360.390 ;
        RECT 1732.020 3360.380 1735.020 3360.390 ;
        RECT 1912.020 3360.380 1915.020 3360.390 ;
        RECT 2092.020 3360.380 2095.020 3360.390 ;
        RECT 2272.020 3360.380 2275.020 3360.390 ;
        RECT 2452.020 3360.380 2455.020 3360.390 ;
        RECT 2632.020 3360.380 2635.020 3360.390 ;
        RECT 2812.020 3360.380 2815.020 3360.390 ;
        RECT 2940.400 3360.380 2943.400 3360.390 ;
        RECT -23.780 3357.380 2943.400 3360.380 ;
        RECT -23.780 3357.370 -20.780 3357.380 ;
        RECT 112.020 3357.370 115.020 3357.380 ;
        RECT 292.020 3357.370 295.020 3357.380 ;
        RECT 472.020 3357.370 475.020 3357.380 ;
        RECT 652.020 3357.370 655.020 3357.380 ;
        RECT 832.020 3357.370 835.020 3357.380 ;
        RECT 1012.020 3357.370 1015.020 3357.380 ;
        RECT 1192.020 3357.370 1195.020 3357.380 ;
        RECT 1372.020 3357.370 1375.020 3357.380 ;
        RECT 1552.020 3357.370 1555.020 3357.380 ;
        RECT 1732.020 3357.370 1735.020 3357.380 ;
        RECT 1912.020 3357.370 1915.020 3357.380 ;
        RECT 2092.020 3357.370 2095.020 3357.380 ;
        RECT 2272.020 3357.370 2275.020 3357.380 ;
        RECT 2452.020 3357.370 2455.020 3357.380 ;
        RECT 2632.020 3357.370 2635.020 3357.380 ;
        RECT 2812.020 3357.370 2815.020 3357.380 ;
        RECT 2940.400 3357.370 2943.400 3357.380 ;
        RECT -23.780 3180.380 -20.780 3180.390 ;
        RECT 112.020 3180.380 115.020 3180.390 ;
        RECT 292.020 3180.380 295.020 3180.390 ;
        RECT 472.020 3180.380 475.020 3180.390 ;
        RECT 652.020 3180.380 655.020 3180.390 ;
        RECT 832.020 3180.380 835.020 3180.390 ;
        RECT 1012.020 3180.380 1015.020 3180.390 ;
        RECT 1192.020 3180.380 1195.020 3180.390 ;
        RECT 1372.020 3180.380 1375.020 3180.390 ;
        RECT 1552.020 3180.380 1555.020 3180.390 ;
        RECT 1732.020 3180.380 1735.020 3180.390 ;
        RECT 1912.020 3180.380 1915.020 3180.390 ;
        RECT 2092.020 3180.380 2095.020 3180.390 ;
        RECT 2272.020 3180.380 2275.020 3180.390 ;
        RECT 2452.020 3180.380 2455.020 3180.390 ;
        RECT 2632.020 3180.380 2635.020 3180.390 ;
        RECT 2812.020 3180.380 2815.020 3180.390 ;
        RECT 2940.400 3180.380 2943.400 3180.390 ;
        RECT -23.780 3177.380 2943.400 3180.380 ;
        RECT -23.780 3177.370 -20.780 3177.380 ;
        RECT 112.020 3177.370 115.020 3177.380 ;
        RECT 292.020 3177.370 295.020 3177.380 ;
        RECT 472.020 3177.370 475.020 3177.380 ;
        RECT 652.020 3177.370 655.020 3177.380 ;
        RECT 832.020 3177.370 835.020 3177.380 ;
        RECT 1012.020 3177.370 1015.020 3177.380 ;
        RECT 1192.020 3177.370 1195.020 3177.380 ;
        RECT 1372.020 3177.370 1375.020 3177.380 ;
        RECT 1552.020 3177.370 1555.020 3177.380 ;
        RECT 1732.020 3177.370 1735.020 3177.380 ;
        RECT 1912.020 3177.370 1915.020 3177.380 ;
        RECT 2092.020 3177.370 2095.020 3177.380 ;
        RECT 2272.020 3177.370 2275.020 3177.380 ;
        RECT 2452.020 3177.370 2455.020 3177.380 ;
        RECT 2632.020 3177.370 2635.020 3177.380 ;
        RECT 2812.020 3177.370 2815.020 3177.380 ;
        RECT 2940.400 3177.370 2943.400 3177.380 ;
        RECT -23.780 3000.380 -20.780 3000.390 ;
        RECT 112.020 3000.380 115.020 3000.390 ;
        RECT 292.020 3000.380 295.020 3000.390 ;
        RECT 472.020 3000.380 475.020 3000.390 ;
        RECT 652.020 3000.380 655.020 3000.390 ;
        RECT 832.020 3000.380 835.020 3000.390 ;
        RECT 1012.020 3000.380 1015.020 3000.390 ;
        RECT 1192.020 3000.380 1195.020 3000.390 ;
        RECT 1372.020 3000.380 1375.020 3000.390 ;
        RECT 1552.020 3000.380 1555.020 3000.390 ;
        RECT 1732.020 3000.380 1735.020 3000.390 ;
        RECT 1912.020 3000.380 1915.020 3000.390 ;
        RECT 2092.020 3000.380 2095.020 3000.390 ;
        RECT 2272.020 3000.380 2275.020 3000.390 ;
        RECT 2452.020 3000.380 2455.020 3000.390 ;
        RECT 2632.020 3000.380 2635.020 3000.390 ;
        RECT 2812.020 3000.380 2815.020 3000.390 ;
        RECT 2940.400 3000.380 2943.400 3000.390 ;
        RECT -23.780 2997.380 2943.400 3000.380 ;
        RECT -23.780 2997.370 -20.780 2997.380 ;
        RECT 112.020 2997.370 115.020 2997.380 ;
        RECT 292.020 2997.370 295.020 2997.380 ;
        RECT 472.020 2997.370 475.020 2997.380 ;
        RECT 652.020 2997.370 655.020 2997.380 ;
        RECT 832.020 2997.370 835.020 2997.380 ;
        RECT 1012.020 2997.370 1015.020 2997.380 ;
        RECT 1192.020 2997.370 1195.020 2997.380 ;
        RECT 1372.020 2997.370 1375.020 2997.380 ;
        RECT 1552.020 2997.370 1555.020 2997.380 ;
        RECT 1732.020 2997.370 1735.020 2997.380 ;
        RECT 1912.020 2997.370 1915.020 2997.380 ;
        RECT 2092.020 2997.370 2095.020 2997.380 ;
        RECT 2272.020 2997.370 2275.020 2997.380 ;
        RECT 2452.020 2997.370 2455.020 2997.380 ;
        RECT 2632.020 2997.370 2635.020 2997.380 ;
        RECT 2812.020 2997.370 2815.020 2997.380 ;
        RECT 2940.400 2997.370 2943.400 2997.380 ;
        RECT -23.780 2820.380 -20.780 2820.390 ;
        RECT 112.020 2820.380 115.020 2820.390 ;
        RECT 292.020 2820.380 295.020 2820.390 ;
        RECT 472.020 2820.380 475.020 2820.390 ;
        RECT 652.020 2820.380 655.020 2820.390 ;
        RECT 832.020 2820.380 835.020 2820.390 ;
        RECT 1012.020 2820.380 1015.020 2820.390 ;
        RECT 1192.020 2820.380 1195.020 2820.390 ;
        RECT 1372.020 2820.380 1375.020 2820.390 ;
        RECT 1552.020 2820.380 1555.020 2820.390 ;
        RECT 1732.020 2820.380 1735.020 2820.390 ;
        RECT 1912.020 2820.380 1915.020 2820.390 ;
        RECT 2092.020 2820.380 2095.020 2820.390 ;
        RECT 2272.020 2820.380 2275.020 2820.390 ;
        RECT 2452.020 2820.380 2455.020 2820.390 ;
        RECT 2632.020 2820.380 2635.020 2820.390 ;
        RECT 2812.020 2820.380 2815.020 2820.390 ;
        RECT 2940.400 2820.380 2943.400 2820.390 ;
        RECT -23.780 2817.380 2943.400 2820.380 ;
        RECT -23.780 2817.370 -20.780 2817.380 ;
        RECT 112.020 2817.370 115.020 2817.380 ;
        RECT 292.020 2817.370 295.020 2817.380 ;
        RECT 472.020 2817.370 475.020 2817.380 ;
        RECT 652.020 2817.370 655.020 2817.380 ;
        RECT 832.020 2817.370 835.020 2817.380 ;
        RECT 1012.020 2817.370 1015.020 2817.380 ;
        RECT 1192.020 2817.370 1195.020 2817.380 ;
        RECT 1372.020 2817.370 1375.020 2817.380 ;
        RECT 1552.020 2817.370 1555.020 2817.380 ;
        RECT 1732.020 2817.370 1735.020 2817.380 ;
        RECT 1912.020 2817.370 1915.020 2817.380 ;
        RECT 2092.020 2817.370 2095.020 2817.380 ;
        RECT 2272.020 2817.370 2275.020 2817.380 ;
        RECT 2452.020 2817.370 2455.020 2817.380 ;
        RECT 2632.020 2817.370 2635.020 2817.380 ;
        RECT 2812.020 2817.370 2815.020 2817.380 ;
        RECT 2940.400 2817.370 2943.400 2817.380 ;
        RECT -23.780 2640.380 -20.780 2640.390 ;
        RECT 112.020 2640.380 115.020 2640.390 ;
        RECT 292.020 2640.380 295.020 2640.390 ;
        RECT 472.020 2640.380 475.020 2640.390 ;
        RECT 652.020 2640.380 655.020 2640.390 ;
        RECT 832.020 2640.380 835.020 2640.390 ;
        RECT 1012.020 2640.380 1015.020 2640.390 ;
        RECT 1192.020 2640.380 1195.020 2640.390 ;
        RECT 1372.020 2640.380 1375.020 2640.390 ;
        RECT 1552.020 2640.380 1555.020 2640.390 ;
        RECT 1732.020 2640.380 1735.020 2640.390 ;
        RECT 1912.020 2640.380 1915.020 2640.390 ;
        RECT 2092.020 2640.380 2095.020 2640.390 ;
        RECT 2272.020 2640.380 2275.020 2640.390 ;
        RECT 2452.020 2640.380 2455.020 2640.390 ;
        RECT 2632.020 2640.380 2635.020 2640.390 ;
        RECT 2812.020 2640.380 2815.020 2640.390 ;
        RECT 2940.400 2640.380 2943.400 2640.390 ;
        RECT -23.780 2637.380 2943.400 2640.380 ;
        RECT -23.780 2637.370 -20.780 2637.380 ;
        RECT 112.020 2637.370 115.020 2637.380 ;
        RECT 292.020 2637.370 295.020 2637.380 ;
        RECT 472.020 2637.370 475.020 2637.380 ;
        RECT 652.020 2637.370 655.020 2637.380 ;
        RECT 832.020 2637.370 835.020 2637.380 ;
        RECT 1012.020 2637.370 1015.020 2637.380 ;
        RECT 1192.020 2637.370 1195.020 2637.380 ;
        RECT 1372.020 2637.370 1375.020 2637.380 ;
        RECT 1552.020 2637.370 1555.020 2637.380 ;
        RECT 1732.020 2637.370 1735.020 2637.380 ;
        RECT 1912.020 2637.370 1915.020 2637.380 ;
        RECT 2092.020 2637.370 2095.020 2637.380 ;
        RECT 2272.020 2637.370 2275.020 2637.380 ;
        RECT 2452.020 2637.370 2455.020 2637.380 ;
        RECT 2632.020 2637.370 2635.020 2637.380 ;
        RECT 2812.020 2637.370 2815.020 2637.380 ;
        RECT 2940.400 2637.370 2943.400 2637.380 ;
        RECT -23.780 2460.380 -20.780 2460.390 ;
        RECT 112.020 2460.380 115.020 2460.390 ;
        RECT 292.020 2460.380 295.020 2460.390 ;
        RECT 472.020 2460.380 475.020 2460.390 ;
        RECT 652.020 2460.380 655.020 2460.390 ;
        RECT 832.020 2460.380 835.020 2460.390 ;
        RECT 1012.020 2460.380 1015.020 2460.390 ;
        RECT 1192.020 2460.380 1195.020 2460.390 ;
        RECT 1372.020 2460.380 1375.020 2460.390 ;
        RECT 1552.020 2460.380 1555.020 2460.390 ;
        RECT 1732.020 2460.380 1735.020 2460.390 ;
        RECT 1912.020 2460.380 1915.020 2460.390 ;
        RECT 2092.020 2460.380 2095.020 2460.390 ;
        RECT 2272.020 2460.380 2275.020 2460.390 ;
        RECT 2452.020 2460.380 2455.020 2460.390 ;
        RECT 2632.020 2460.380 2635.020 2460.390 ;
        RECT 2812.020 2460.380 2815.020 2460.390 ;
        RECT 2940.400 2460.380 2943.400 2460.390 ;
        RECT -23.780 2457.380 2943.400 2460.380 ;
        RECT -23.780 2457.370 -20.780 2457.380 ;
        RECT 112.020 2457.370 115.020 2457.380 ;
        RECT 292.020 2457.370 295.020 2457.380 ;
        RECT 472.020 2457.370 475.020 2457.380 ;
        RECT 652.020 2457.370 655.020 2457.380 ;
        RECT 832.020 2457.370 835.020 2457.380 ;
        RECT 1012.020 2457.370 1015.020 2457.380 ;
        RECT 1192.020 2457.370 1195.020 2457.380 ;
        RECT 1372.020 2457.370 1375.020 2457.380 ;
        RECT 1552.020 2457.370 1555.020 2457.380 ;
        RECT 1732.020 2457.370 1735.020 2457.380 ;
        RECT 1912.020 2457.370 1915.020 2457.380 ;
        RECT 2092.020 2457.370 2095.020 2457.380 ;
        RECT 2272.020 2457.370 2275.020 2457.380 ;
        RECT 2452.020 2457.370 2455.020 2457.380 ;
        RECT 2632.020 2457.370 2635.020 2457.380 ;
        RECT 2812.020 2457.370 2815.020 2457.380 ;
        RECT 2940.400 2457.370 2943.400 2457.380 ;
        RECT -23.780 2280.380 -20.780 2280.390 ;
        RECT 112.020 2280.380 115.020 2280.390 ;
        RECT 292.020 2280.380 295.020 2280.390 ;
        RECT 472.020 2280.380 475.020 2280.390 ;
        RECT 652.020 2280.380 655.020 2280.390 ;
        RECT 832.020 2280.380 835.020 2280.390 ;
        RECT 1012.020 2280.380 1015.020 2280.390 ;
        RECT 1192.020 2280.380 1195.020 2280.390 ;
        RECT 1372.020 2280.380 1375.020 2280.390 ;
        RECT 1552.020 2280.380 1555.020 2280.390 ;
        RECT 1732.020 2280.380 1735.020 2280.390 ;
        RECT 1912.020 2280.380 1915.020 2280.390 ;
        RECT 2092.020 2280.380 2095.020 2280.390 ;
        RECT 2272.020 2280.380 2275.020 2280.390 ;
        RECT 2452.020 2280.380 2455.020 2280.390 ;
        RECT 2632.020 2280.380 2635.020 2280.390 ;
        RECT 2812.020 2280.380 2815.020 2280.390 ;
        RECT 2940.400 2280.380 2943.400 2280.390 ;
        RECT -23.780 2277.380 2943.400 2280.380 ;
        RECT -23.780 2277.370 -20.780 2277.380 ;
        RECT 112.020 2277.370 115.020 2277.380 ;
        RECT 292.020 2277.370 295.020 2277.380 ;
        RECT 472.020 2277.370 475.020 2277.380 ;
        RECT 652.020 2277.370 655.020 2277.380 ;
        RECT 832.020 2277.370 835.020 2277.380 ;
        RECT 1012.020 2277.370 1015.020 2277.380 ;
        RECT 1192.020 2277.370 1195.020 2277.380 ;
        RECT 1372.020 2277.370 1375.020 2277.380 ;
        RECT 1552.020 2277.370 1555.020 2277.380 ;
        RECT 1732.020 2277.370 1735.020 2277.380 ;
        RECT 1912.020 2277.370 1915.020 2277.380 ;
        RECT 2092.020 2277.370 2095.020 2277.380 ;
        RECT 2272.020 2277.370 2275.020 2277.380 ;
        RECT 2452.020 2277.370 2455.020 2277.380 ;
        RECT 2632.020 2277.370 2635.020 2277.380 ;
        RECT 2812.020 2277.370 2815.020 2277.380 ;
        RECT 2940.400 2277.370 2943.400 2277.380 ;
        RECT -23.780 2100.380 -20.780 2100.390 ;
        RECT 112.020 2100.380 115.020 2100.390 ;
        RECT 292.020 2100.380 295.020 2100.390 ;
        RECT 472.020 2100.380 475.020 2100.390 ;
        RECT 652.020 2100.380 655.020 2100.390 ;
        RECT 832.020 2100.380 835.020 2100.390 ;
        RECT 1012.020 2100.380 1015.020 2100.390 ;
        RECT 1192.020 2100.380 1195.020 2100.390 ;
        RECT 1372.020 2100.380 1375.020 2100.390 ;
        RECT 1552.020 2100.380 1555.020 2100.390 ;
        RECT 1732.020 2100.380 1735.020 2100.390 ;
        RECT 1912.020 2100.380 1915.020 2100.390 ;
        RECT 2092.020 2100.380 2095.020 2100.390 ;
        RECT 2272.020 2100.380 2275.020 2100.390 ;
        RECT 2452.020 2100.380 2455.020 2100.390 ;
        RECT 2632.020 2100.380 2635.020 2100.390 ;
        RECT 2812.020 2100.380 2815.020 2100.390 ;
        RECT 2940.400 2100.380 2943.400 2100.390 ;
        RECT -23.780 2097.380 2943.400 2100.380 ;
        RECT -23.780 2097.370 -20.780 2097.380 ;
        RECT 112.020 2097.370 115.020 2097.380 ;
        RECT 292.020 2097.370 295.020 2097.380 ;
        RECT 472.020 2097.370 475.020 2097.380 ;
        RECT 652.020 2097.370 655.020 2097.380 ;
        RECT 832.020 2097.370 835.020 2097.380 ;
        RECT 1012.020 2097.370 1015.020 2097.380 ;
        RECT 1192.020 2097.370 1195.020 2097.380 ;
        RECT 1372.020 2097.370 1375.020 2097.380 ;
        RECT 1552.020 2097.370 1555.020 2097.380 ;
        RECT 1732.020 2097.370 1735.020 2097.380 ;
        RECT 1912.020 2097.370 1915.020 2097.380 ;
        RECT 2092.020 2097.370 2095.020 2097.380 ;
        RECT 2272.020 2097.370 2275.020 2097.380 ;
        RECT 2452.020 2097.370 2455.020 2097.380 ;
        RECT 2632.020 2097.370 2635.020 2097.380 ;
        RECT 2812.020 2097.370 2815.020 2097.380 ;
        RECT 2940.400 2097.370 2943.400 2097.380 ;
        RECT -23.780 1920.380 -20.780 1920.390 ;
        RECT 112.020 1920.380 115.020 1920.390 ;
        RECT 292.020 1920.380 295.020 1920.390 ;
        RECT 472.020 1920.380 475.020 1920.390 ;
        RECT 652.020 1920.380 655.020 1920.390 ;
        RECT 832.020 1920.380 835.020 1920.390 ;
        RECT 1012.020 1920.380 1015.020 1920.390 ;
        RECT 1192.020 1920.380 1195.020 1920.390 ;
        RECT 1372.020 1920.380 1375.020 1920.390 ;
        RECT 1552.020 1920.380 1555.020 1920.390 ;
        RECT 1732.020 1920.380 1735.020 1920.390 ;
        RECT 1912.020 1920.380 1915.020 1920.390 ;
        RECT 2092.020 1920.380 2095.020 1920.390 ;
        RECT 2272.020 1920.380 2275.020 1920.390 ;
        RECT 2452.020 1920.380 2455.020 1920.390 ;
        RECT 2632.020 1920.380 2635.020 1920.390 ;
        RECT 2812.020 1920.380 2815.020 1920.390 ;
        RECT 2940.400 1920.380 2943.400 1920.390 ;
        RECT -23.780 1917.380 2943.400 1920.380 ;
        RECT -23.780 1917.370 -20.780 1917.380 ;
        RECT 112.020 1917.370 115.020 1917.380 ;
        RECT 292.020 1917.370 295.020 1917.380 ;
        RECT 472.020 1917.370 475.020 1917.380 ;
        RECT 652.020 1917.370 655.020 1917.380 ;
        RECT 832.020 1917.370 835.020 1917.380 ;
        RECT 1012.020 1917.370 1015.020 1917.380 ;
        RECT 1192.020 1917.370 1195.020 1917.380 ;
        RECT 1372.020 1917.370 1375.020 1917.380 ;
        RECT 1552.020 1917.370 1555.020 1917.380 ;
        RECT 1732.020 1917.370 1735.020 1917.380 ;
        RECT 1912.020 1917.370 1915.020 1917.380 ;
        RECT 2092.020 1917.370 2095.020 1917.380 ;
        RECT 2272.020 1917.370 2275.020 1917.380 ;
        RECT 2452.020 1917.370 2455.020 1917.380 ;
        RECT 2632.020 1917.370 2635.020 1917.380 ;
        RECT 2812.020 1917.370 2815.020 1917.380 ;
        RECT 2940.400 1917.370 2943.400 1917.380 ;
        RECT -23.780 1740.380 -20.780 1740.390 ;
        RECT 112.020 1740.380 115.020 1740.390 ;
        RECT 292.020 1740.380 295.020 1740.390 ;
        RECT 472.020 1740.380 475.020 1740.390 ;
        RECT 652.020 1740.380 655.020 1740.390 ;
        RECT 832.020 1740.380 835.020 1740.390 ;
        RECT 1012.020 1740.380 1015.020 1740.390 ;
        RECT 1192.020 1740.380 1195.020 1740.390 ;
        RECT 1372.020 1740.380 1375.020 1740.390 ;
        RECT 1552.020 1740.380 1555.020 1740.390 ;
        RECT 1732.020 1740.380 1735.020 1740.390 ;
        RECT 1912.020 1740.380 1915.020 1740.390 ;
        RECT 2092.020 1740.380 2095.020 1740.390 ;
        RECT 2272.020 1740.380 2275.020 1740.390 ;
        RECT 2452.020 1740.380 2455.020 1740.390 ;
        RECT 2632.020 1740.380 2635.020 1740.390 ;
        RECT 2812.020 1740.380 2815.020 1740.390 ;
        RECT 2940.400 1740.380 2943.400 1740.390 ;
        RECT -23.780 1737.380 2943.400 1740.380 ;
        RECT -23.780 1737.370 -20.780 1737.380 ;
        RECT 112.020 1737.370 115.020 1737.380 ;
        RECT 292.020 1737.370 295.020 1737.380 ;
        RECT 472.020 1737.370 475.020 1737.380 ;
        RECT 652.020 1737.370 655.020 1737.380 ;
        RECT 832.020 1737.370 835.020 1737.380 ;
        RECT 1012.020 1737.370 1015.020 1737.380 ;
        RECT 1192.020 1737.370 1195.020 1737.380 ;
        RECT 1372.020 1737.370 1375.020 1737.380 ;
        RECT 1552.020 1737.370 1555.020 1737.380 ;
        RECT 1732.020 1737.370 1735.020 1737.380 ;
        RECT 1912.020 1737.370 1915.020 1737.380 ;
        RECT 2092.020 1737.370 2095.020 1737.380 ;
        RECT 2272.020 1737.370 2275.020 1737.380 ;
        RECT 2452.020 1737.370 2455.020 1737.380 ;
        RECT 2632.020 1737.370 2635.020 1737.380 ;
        RECT 2812.020 1737.370 2815.020 1737.380 ;
        RECT 2940.400 1737.370 2943.400 1737.380 ;
        RECT -23.780 1560.380 -20.780 1560.390 ;
        RECT 112.020 1560.380 115.020 1560.390 ;
        RECT 292.020 1560.380 295.020 1560.390 ;
        RECT 472.020 1560.380 475.020 1560.390 ;
        RECT 652.020 1560.380 655.020 1560.390 ;
        RECT 832.020 1560.380 835.020 1560.390 ;
        RECT 1012.020 1560.380 1015.020 1560.390 ;
        RECT 1192.020 1560.380 1195.020 1560.390 ;
        RECT 1372.020 1560.380 1375.020 1560.390 ;
        RECT 1552.020 1560.380 1555.020 1560.390 ;
        RECT 1732.020 1560.380 1735.020 1560.390 ;
        RECT 1912.020 1560.380 1915.020 1560.390 ;
        RECT 2092.020 1560.380 2095.020 1560.390 ;
        RECT 2272.020 1560.380 2275.020 1560.390 ;
        RECT 2452.020 1560.380 2455.020 1560.390 ;
        RECT 2632.020 1560.380 2635.020 1560.390 ;
        RECT 2812.020 1560.380 2815.020 1560.390 ;
        RECT 2940.400 1560.380 2943.400 1560.390 ;
        RECT -23.780 1557.380 2943.400 1560.380 ;
        RECT -23.780 1557.370 -20.780 1557.380 ;
        RECT 112.020 1557.370 115.020 1557.380 ;
        RECT 292.020 1557.370 295.020 1557.380 ;
        RECT 472.020 1557.370 475.020 1557.380 ;
        RECT 652.020 1557.370 655.020 1557.380 ;
        RECT 832.020 1557.370 835.020 1557.380 ;
        RECT 1012.020 1557.370 1015.020 1557.380 ;
        RECT 1192.020 1557.370 1195.020 1557.380 ;
        RECT 1372.020 1557.370 1375.020 1557.380 ;
        RECT 1552.020 1557.370 1555.020 1557.380 ;
        RECT 1732.020 1557.370 1735.020 1557.380 ;
        RECT 1912.020 1557.370 1915.020 1557.380 ;
        RECT 2092.020 1557.370 2095.020 1557.380 ;
        RECT 2272.020 1557.370 2275.020 1557.380 ;
        RECT 2452.020 1557.370 2455.020 1557.380 ;
        RECT 2632.020 1557.370 2635.020 1557.380 ;
        RECT 2812.020 1557.370 2815.020 1557.380 ;
        RECT 2940.400 1557.370 2943.400 1557.380 ;
        RECT -23.780 1380.380 -20.780 1380.390 ;
        RECT 112.020 1380.380 115.020 1380.390 ;
        RECT 292.020 1380.380 295.020 1380.390 ;
        RECT 472.020 1380.380 475.020 1380.390 ;
        RECT 652.020 1380.380 655.020 1380.390 ;
        RECT 832.020 1380.380 835.020 1380.390 ;
        RECT 1012.020 1380.380 1015.020 1380.390 ;
        RECT 1192.020 1380.380 1195.020 1380.390 ;
        RECT 1372.020 1380.380 1375.020 1380.390 ;
        RECT 1552.020 1380.380 1555.020 1380.390 ;
        RECT 1732.020 1380.380 1735.020 1380.390 ;
        RECT 1912.020 1380.380 1915.020 1380.390 ;
        RECT 2092.020 1380.380 2095.020 1380.390 ;
        RECT 2272.020 1380.380 2275.020 1380.390 ;
        RECT 2452.020 1380.380 2455.020 1380.390 ;
        RECT 2632.020 1380.380 2635.020 1380.390 ;
        RECT 2812.020 1380.380 2815.020 1380.390 ;
        RECT 2940.400 1380.380 2943.400 1380.390 ;
        RECT -23.780 1377.380 2943.400 1380.380 ;
        RECT -23.780 1377.370 -20.780 1377.380 ;
        RECT 112.020 1377.370 115.020 1377.380 ;
        RECT 292.020 1377.370 295.020 1377.380 ;
        RECT 472.020 1377.370 475.020 1377.380 ;
        RECT 652.020 1377.370 655.020 1377.380 ;
        RECT 832.020 1377.370 835.020 1377.380 ;
        RECT 1012.020 1377.370 1015.020 1377.380 ;
        RECT 1192.020 1377.370 1195.020 1377.380 ;
        RECT 1372.020 1377.370 1375.020 1377.380 ;
        RECT 1552.020 1377.370 1555.020 1377.380 ;
        RECT 1732.020 1377.370 1735.020 1377.380 ;
        RECT 1912.020 1377.370 1915.020 1377.380 ;
        RECT 2092.020 1377.370 2095.020 1377.380 ;
        RECT 2272.020 1377.370 2275.020 1377.380 ;
        RECT 2452.020 1377.370 2455.020 1377.380 ;
        RECT 2632.020 1377.370 2635.020 1377.380 ;
        RECT 2812.020 1377.370 2815.020 1377.380 ;
        RECT 2940.400 1377.370 2943.400 1377.380 ;
        RECT -23.780 1200.380 -20.780 1200.390 ;
        RECT 112.020 1200.380 115.020 1200.390 ;
        RECT 292.020 1200.380 295.020 1200.390 ;
        RECT 472.020 1200.380 475.020 1200.390 ;
        RECT 652.020 1200.380 655.020 1200.390 ;
        RECT 832.020 1200.380 835.020 1200.390 ;
        RECT 1012.020 1200.380 1015.020 1200.390 ;
        RECT 1192.020 1200.380 1195.020 1200.390 ;
        RECT 1372.020 1200.380 1375.020 1200.390 ;
        RECT 1552.020 1200.380 1555.020 1200.390 ;
        RECT 1732.020 1200.380 1735.020 1200.390 ;
        RECT 1912.020 1200.380 1915.020 1200.390 ;
        RECT 2092.020 1200.380 2095.020 1200.390 ;
        RECT 2272.020 1200.380 2275.020 1200.390 ;
        RECT 2452.020 1200.380 2455.020 1200.390 ;
        RECT 2632.020 1200.380 2635.020 1200.390 ;
        RECT 2812.020 1200.380 2815.020 1200.390 ;
        RECT 2940.400 1200.380 2943.400 1200.390 ;
        RECT -23.780 1197.380 2943.400 1200.380 ;
        RECT -23.780 1197.370 -20.780 1197.380 ;
        RECT 112.020 1197.370 115.020 1197.380 ;
        RECT 292.020 1197.370 295.020 1197.380 ;
        RECT 472.020 1197.370 475.020 1197.380 ;
        RECT 652.020 1197.370 655.020 1197.380 ;
        RECT 832.020 1197.370 835.020 1197.380 ;
        RECT 1012.020 1197.370 1015.020 1197.380 ;
        RECT 1192.020 1197.370 1195.020 1197.380 ;
        RECT 1372.020 1197.370 1375.020 1197.380 ;
        RECT 1552.020 1197.370 1555.020 1197.380 ;
        RECT 1732.020 1197.370 1735.020 1197.380 ;
        RECT 1912.020 1197.370 1915.020 1197.380 ;
        RECT 2092.020 1197.370 2095.020 1197.380 ;
        RECT 2272.020 1197.370 2275.020 1197.380 ;
        RECT 2452.020 1197.370 2455.020 1197.380 ;
        RECT 2632.020 1197.370 2635.020 1197.380 ;
        RECT 2812.020 1197.370 2815.020 1197.380 ;
        RECT 2940.400 1197.370 2943.400 1197.380 ;
        RECT -23.780 1020.380 -20.780 1020.390 ;
        RECT 112.020 1020.380 115.020 1020.390 ;
        RECT 292.020 1020.380 295.020 1020.390 ;
        RECT 472.020 1020.380 475.020 1020.390 ;
        RECT 652.020 1020.380 655.020 1020.390 ;
        RECT 832.020 1020.380 835.020 1020.390 ;
        RECT 1012.020 1020.380 1015.020 1020.390 ;
        RECT 1192.020 1020.380 1195.020 1020.390 ;
        RECT 1372.020 1020.380 1375.020 1020.390 ;
        RECT 1552.020 1020.380 1555.020 1020.390 ;
        RECT 1732.020 1020.380 1735.020 1020.390 ;
        RECT 1912.020 1020.380 1915.020 1020.390 ;
        RECT 2092.020 1020.380 2095.020 1020.390 ;
        RECT 2272.020 1020.380 2275.020 1020.390 ;
        RECT 2452.020 1020.380 2455.020 1020.390 ;
        RECT 2632.020 1020.380 2635.020 1020.390 ;
        RECT 2812.020 1020.380 2815.020 1020.390 ;
        RECT 2940.400 1020.380 2943.400 1020.390 ;
        RECT -23.780 1017.380 2943.400 1020.380 ;
        RECT -23.780 1017.370 -20.780 1017.380 ;
        RECT 112.020 1017.370 115.020 1017.380 ;
        RECT 292.020 1017.370 295.020 1017.380 ;
        RECT 472.020 1017.370 475.020 1017.380 ;
        RECT 652.020 1017.370 655.020 1017.380 ;
        RECT 832.020 1017.370 835.020 1017.380 ;
        RECT 1012.020 1017.370 1015.020 1017.380 ;
        RECT 1192.020 1017.370 1195.020 1017.380 ;
        RECT 1372.020 1017.370 1375.020 1017.380 ;
        RECT 1552.020 1017.370 1555.020 1017.380 ;
        RECT 1732.020 1017.370 1735.020 1017.380 ;
        RECT 1912.020 1017.370 1915.020 1017.380 ;
        RECT 2092.020 1017.370 2095.020 1017.380 ;
        RECT 2272.020 1017.370 2275.020 1017.380 ;
        RECT 2452.020 1017.370 2455.020 1017.380 ;
        RECT 2632.020 1017.370 2635.020 1017.380 ;
        RECT 2812.020 1017.370 2815.020 1017.380 ;
        RECT 2940.400 1017.370 2943.400 1017.380 ;
        RECT -23.780 840.380 -20.780 840.390 ;
        RECT 112.020 840.380 115.020 840.390 ;
        RECT 292.020 840.380 295.020 840.390 ;
        RECT 472.020 840.380 475.020 840.390 ;
        RECT 652.020 840.380 655.020 840.390 ;
        RECT 832.020 840.380 835.020 840.390 ;
        RECT 1012.020 840.380 1015.020 840.390 ;
        RECT 1192.020 840.380 1195.020 840.390 ;
        RECT 1372.020 840.380 1375.020 840.390 ;
        RECT 1552.020 840.380 1555.020 840.390 ;
        RECT 1732.020 840.380 1735.020 840.390 ;
        RECT 1912.020 840.380 1915.020 840.390 ;
        RECT 2092.020 840.380 2095.020 840.390 ;
        RECT 2272.020 840.380 2275.020 840.390 ;
        RECT 2452.020 840.380 2455.020 840.390 ;
        RECT 2632.020 840.380 2635.020 840.390 ;
        RECT 2812.020 840.380 2815.020 840.390 ;
        RECT 2940.400 840.380 2943.400 840.390 ;
        RECT -23.780 837.380 2943.400 840.380 ;
        RECT -23.780 837.370 -20.780 837.380 ;
        RECT 112.020 837.370 115.020 837.380 ;
        RECT 292.020 837.370 295.020 837.380 ;
        RECT 472.020 837.370 475.020 837.380 ;
        RECT 652.020 837.370 655.020 837.380 ;
        RECT 832.020 837.370 835.020 837.380 ;
        RECT 1012.020 837.370 1015.020 837.380 ;
        RECT 1192.020 837.370 1195.020 837.380 ;
        RECT 1372.020 837.370 1375.020 837.380 ;
        RECT 1552.020 837.370 1555.020 837.380 ;
        RECT 1732.020 837.370 1735.020 837.380 ;
        RECT 1912.020 837.370 1915.020 837.380 ;
        RECT 2092.020 837.370 2095.020 837.380 ;
        RECT 2272.020 837.370 2275.020 837.380 ;
        RECT 2452.020 837.370 2455.020 837.380 ;
        RECT 2632.020 837.370 2635.020 837.380 ;
        RECT 2812.020 837.370 2815.020 837.380 ;
        RECT 2940.400 837.370 2943.400 837.380 ;
        RECT -23.780 660.380 -20.780 660.390 ;
        RECT 112.020 660.380 115.020 660.390 ;
        RECT 292.020 660.380 295.020 660.390 ;
        RECT 472.020 660.380 475.020 660.390 ;
        RECT 652.020 660.380 655.020 660.390 ;
        RECT 832.020 660.380 835.020 660.390 ;
        RECT 1012.020 660.380 1015.020 660.390 ;
        RECT 1192.020 660.380 1195.020 660.390 ;
        RECT 1372.020 660.380 1375.020 660.390 ;
        RECT 1552.020 660.380 1555.020 660.390 ;
        RECT 1732.020 660.380 1735.020 660.390 ;
        RECT 1912.020 660.380 1915.020 660.390 ;
        RECT 2092.020 660.380 2095.020 660.390 ;
        RECT 2272.020 660.380 2275.020 660.390 ;
        RECT 2452.020 660.380 2455.020 660.390 ;
        RECT 2632.020 660.380 2635.020 660.390 ;
        RECT 2812.020 660.380 2815.020 660.390 ;
        RECT 2940.400 660.380 2943.400 660.390 ;
        RECT -23.780 657.380 2943.400 660.380 ;
        RECT -23.780 657.370 -20.780 657.380 ;
        RECT 112.020 657.370 115.020 657.380 ;
        RECT 292.020 657.370 295.020 657.380 ;
        RECT 472.020 657.370 475.020 657.380 ;
        RECT 652.020 657.370 655.020 657.380 ;
        RECT 832.020 657.370 835.020 657.380 ;
        RECT 1012.020 657.370 1015.020 657.380 ;
        RECT 1192.020 657.370 1195.020 657.380 ;
        RECT 1372.020 657.370 1375.020 657.380 ;
        RECT 1552.020 657.370 1555.020 657.380 ;
        RECT 1732.020 657.370 1735.020 657.380 ;
        RECT 1912.020 657.370 1915.020 657.380 ;
        RECT 2092.020 657.370 2095.020 657.380 ;
        RECT 2272.020 657.370 2275.020 657.380 ;
        RECT 2452.020 657.370 2455.020 657.380 ;
        RECT 2632.020 657.370 2635.020 657.380 ;
        RECT 2812.020 657.370 2815.020 657.380 ;
        RECT 2940.400 657.370 2943.400 657.380 ;
        RECT -23.780 480.380 -20.780 480.390 ;
        RECT 112.020 480.380 115.020 480.390 ;
        RECT 292.020 480.380 295.020 480.390 ;
        RECT 472.020 480.380 475.020 480.390 ;
        RECT 652.020 480.380 655.020 480.390 ;
        RECT 832.020 480.380 835.020 480.390 ;
        RECT 1012.020 480.380 1015.020 480.390 ;
        RECT 1192.020 480.380 1195.020 480.390 ;
        RECT 1372.020 480.380 1375.020 480.390 ;
        RECT 1552.020 480.380 1555.020 480.390 ;
        RECT 1732.020 480.380 1735.020 480.390 ;
        RECT 1912.020 480.380 1915.020 480.390 ;
        RECT 2092.020 480.380 2095.020 480.390 ;
        RECT 2272.020 480.380 2275.020 480.390 ;
        RECT 2452.020 480.380 2455.020 480.390 ;
        RECT 2632.020 480.380 2635.020 480.390 ;
        RECT 2812.020 480.380 2815.020 480.390 ;
        RECT 2940.400 480.380 2943.400 480.390 ;
        RECT -23.780 477.380 2943.400 480.380 ;
        RECT -23.780 477.370 -20.780 477.380 ;
        RECT 112.020 477.370 115.020 477.380 ;
        RECT 292.020 477.370 295.020 477.380 ;
        RECT 472.020 477.370 475.020 477.380 ;
        RECT 652.020 477.370 655.020 477.380 ;
        RECT 832.020 477.370 835.020 477.380 ;
        RECT 1012.020 477.370 1015.020 477.380 ;
        RECT 1192.020 477.370 1195.020 477.380 ;
        RECT 1372.020 477.370 1375.020 477.380 ;
        RECT 1552.020 477.370 1555.020 477.380 ;
        RECT 1732.020 477.370 1735.020 477.380 ;
        RECT 1912.020 477.370 1915.020 477.380 ;
        RECT 2092.020 477.370 2095.020 477.380 ;
        RECT 2272.020 477.370 2275.020 477.380 ;
        RECT 2452.020 477.370 2455.020 477.380 ;
        RECT 2632.020 477.370 2635.020 477.380 ;
        RECT 2812.020 477.370 2815.020 477.380 ;
        RECT 2940.400 477.370 2943.400 477.380 ;
        RECT -23.780 300.380 -20.780 300.390 ;
        RECT 112.020 300.380 115.020 300.390 ;
        RECT 292.020 300.380 295.020 300.390 ;
        RECT 472.020 300.380 475.020 300.390 ;
        RECT 652.020 300.380 655.020 300.390 ;
        RECT 832.020 300.380 835.020 300.390 ;
        RECT 1012.020 300.380 1015.020 300.390 ;
        RECT 1192.020 300.380 1195.020 300.390 ;
        RECT 1372.020 300.380 1375.020 300.390 ;
        RECT 1552.020 300.380 1555.020 300.390 ;
        RECT 1732.020 300.380 1735.020 300.390 ;
        RECT 1912.020 300.380 1915.020 300.390 ;
        RECT 2092.020 300.380 2095.020 300.390 ;
        RECT 2272.020 300.380 2275.020 300.390 ;
        RECT 2452.020 300.380 2455.020 300.390 ;
        RECT 2632.020 300.380 2635.020 300.390 ;
        RECT 2812.020 300.380 2815.020 300.390 ;
        RECT 2940.400 300.380 2943.400 300.390 ;
        RECT -23.780 297.380 2943.400 300.380 ;
        RECT -23.780 297.370 -20.780 297.380 ;
        RECT 112.020 297.370 115.020 297.380 ;
        RECT 292.020 297.370 295.020 297.380 ;
        RECT 472.020 297.370 475.020 297.380 ;
        RECT 652.020 297.370 655.020 297.380 ;
        RECT 832.020 297.370 835.020 297.380 ;
        RECT 1012.020 297.370 1015.020 297.380 ;
        RECT 1192.020 297.370 1195.020 297.380 ;
        RECT 1372.020 297.370 1375.020 297.380 ;
        RECT 1552.020 297.370 1555.020 297.380 ;
        RECT 1732.020 297.370 1735.020 297.380 ;
        RECT 1912.020 297.370 1915.020 297.380 ;
        RECT 2092.020 297.370 2095.020 297.380 ;
        RECT 2272.020 297.370 2275.020 297.380 ;
        RECT 2452.020 297.370 2455.020 297.380 ;
        RECT 2632.020 297.370 2635.020 297.380 ;
        RECT 2812.020 297.370 2815.020 297.380 ;
        RECT 2940.400 297.370 2943.400 297.380 ;
        RECT -23.780 120.380 -20.780 120.390 ;
        RECT 112.020 120.380 115.020 120.390 ;
        RECT 292.020 120.380 295.020 120.390 ;
        RECT 472.020 120.380 475.020 120.390 ;
        RECT 652.020 120.380 655.020 120.390 ;
        RECT 832.020 120.380 835.020 120.390 ;
        RECT 1012.020 120.380 1015.020 120.390 ;
        RECT 1192.020 120.380 1195.020 120.390 ;
        RECT 1372.020 120.380 1375.020 120.390 ;
        RECT 1552.020 120.380 1555.020 120.390 ;
        RECT 1732.020 120.380 1735.020 120.390 ;
        RECT 1912.020 120.380 1915.020 120.390 ;
        RECT 2092.020 120.380 2095.020 120.390 ;
        RECT 2272.020 120.380 2275.020 120.390 ;
        RECT 2452.020 120.380 2455.020 120.390 ;
        RECT 2632.020 120.380 2635.020 120.390 ;
        RECT 2812.020 120.380 2815.020 120.390 ;
        RECT 2940.400 120.380 2943.400 120.390 ;
        RECT -23.780 117.380 2943.400 120.380 ;
        RECT -23.780 117.370 -20.780 117.380 ;
        RECT 112.020 117.370 115.020 117.380 ;
        RECT 292.020 117.370 295.020 117.380 ;
        RECT 472.020 117.370 475.020 117.380 ;
        RECT 652.020 117.370 655.020 117.380 ;
        RECT 832.020 117.370 835.020 117.380 ;
        RECT 1012.020 117.370 1015.020 117.380 ;
        RECT 1192.020 117.370 1195.020 117.380 ;
        RECT 1372.020 117.370 1375.020 117.380 ;
        RECT 1552.020 117.370 1555.020 117.380 ;
        RECT 1732.020 117.370 1735.020 117.380 ;
        RECT 1912.020 117.370 1915.020 117.380 ;
        RECT 2092.020 117.370 2095.020 117.380 ;
        RECT 2272.020 117.370 2275.020 117.380 ;
        RECT 2452.020 117.370 2455.020 117.380 ;
        RECT 2632.020 117.370 2635.020 117.380 ;
        RECT 2812.020 117.370 2815.020 117.380 ;
        RECT 2940.400 117.370 2943.400 117.380 ;
        RECT -23.780 -15.420 -20.780 -15.410 ;
        RECT 112.020 -15.420 115.020 -15.410 ;
        RECT 292.020 -15.420 295.020 -15.410 ;
        RECT 472.020 -15.420 475.020 -15.410 ;
        RECT 652.020 -15.420 655.020 -15.410 ;
        RECT 832.020 -15.420 835.020 -15.410 ;
        RECT 1012.020 -15.420 1015.020 -15.410 ;
        RECT 1192.020 -15.420 1195.020 -15.410 ;
        RECT 1372.020 -15.420 1375.020 -15.410 ;
        RECT 1552.020 -15.420 1555.020 -15.410 ;
        RECT 1732.020 -15.420 1735.020 -15.410 ;
        RECT 1912.020 -15.420 1915.020 -15.410 ;
        RECT 2092.020 -15.420 2095.020 -15.410 ;
        RECT 2272.020 -15.420 2275.020 -15.410 ;
        RECT 2452.020 -15.420 2455.020 -15.410 ;
        RECT 2632.020 -15.420 2635.020 -15.410 ;
        RECT 2812.020 -15.420 2815.020 -15.410 ;
        RECT 2940.400 -15.420 2943.400 -15.410 ;
        RECT -23.780 -18.420 2943.400 -15.420 ;
        RECT -23.780 -18.430 -20.780 -18.420 ;
        RECT 112.020 -18.430 115.020 -18.420 ;
        RECT 292.020 -18.430 295.020 -18.420 ;
        RECT 472.020 -18.430 475.020 -18.420 ;
        RECT 652.020 -18.430 655.020 -18.420 ;
        RECT 832.020 -18.430 835.020 -18.420 ;
        RECT 1012.020 -18.430 1015.020 -18.420 ;
        RECT 1192.020 -18.430 1195.020 -18.420 ;
        RECT 1372.020 -18.430 1375.020 -18.420 ;
        RECT 1552.020 -18.430 1555.020 -18.420 ;
        RECT 1732.020 -18.430 1735.020 -18.420 ;
        RECT 1912.020 -18.430 1915.020 -18.420 ;
        RECT 2092.020 -18.430 2095.020 -18.420 ;
        RECT 2272.020 -18.430 2275.020 -18.420 ;
        RECT 2452.020 -18.430 2455.020 -18.420 ;
        RECT 2632.020 -18.430 2635.020 -18.420 ;
        RECT 2812.020 -18.430 2815.020 -18.420 ;
        RECT 2940.400 -18.430 2943.400 -18.420 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -28.380 -23.020 -25.380 3542.700 ;
        RECT 40.020 -27.620 43.020 3547.300 ;
        RECT 220.020 -27.620 223.020 3547.300 ;
        RECT 400.020 -27.620 403.020 3547.300 ;
        RECT 580.020 -27.620 583.020 3547.300 ;
        RECT 760.020 -27.620 763.020 3547.300 ;
        RECT 940.020 -27.620 943.020 3547.300 ;
        RECT 1120.020 -27.620 1123.020 3547.300 ;
        RECT 1300.020 -27.620 1303.020 3547.300 ;
        RECT 1480.020 -27.620 1483.020 3547.300 ;
        RECT 1660.020 -27.620 1663.020 3547.300 ;
        RECT 1840.020 -27.620 1843.020 3547.300 ;
        RECT 2020.020 -27.620 2023.020 3547.300 ;
        RECT 2200.020 -27.620 2203.020 3547.300 ;
        RECT 2380.020 -27.620 2383.020 3547.300 ;
        RECT 2560.020 -27.620 2563.020 3547.300 ;
        RECT 2740.020 -27.620 2743.020 3547.300 ;
        RECT 2945.000 -23.020 2948.000 3542.700 ;
      LAYER via4 ;
        RECT -27.470 3541.410 -26.290 3542.590 ;
        RECT -27.470 3539.810 -26.290 3540.990 ;
        RECT -27.470 3467.090 -26.290 3468.270 ;
        RECT -27.470 3465.490 -26.290 3466.670 ;
        RECT -27.470 3287.090 -26.290 3288.270 ;
        RECT -27.470 3285.490 -26.290 3286.670 ;
        RECT -27.470 3107.090 -26.290 3108.270 ;
        RECT -27.470 3105.490 -26.290 3106.670 ;
        RECT -27.470 2927.090 -26.290 2928.270 ;
        RECT -27.470 2925.490 -26.290 2926.670 ;
        RECT -27.470 2747.090 -26.290 2748.270 ;
        RECT -27.470 2745.490 -26.290 2746.670 ;
        RECT -27.470 2567.090 -26.290 2568.270 ;
        RECT -27.470 2565.490 -26.290 2566.670 ;
        RECT -27.470 2387.090 -26.290 2388.270 ;
        RECT -27.470 2385.490 -26.290 2386.670 ;
        RECT -27.470 2207.090 -26.290 2208.270 ;
        RECT -27.470 2205.490 -26.290 2206.670 ;
        RECT -27.470 2027.090 -26.290 2028.270 ;
        RECT -27.470 2025.490 -26.290 2026.670 ;
        RECT -27.470 1847.090 -26.290 1848.270 ;
        RECT -27.470 1845.490 -26.290 1846.670 ;
        RECT -27.470 1667.090 -26.290 1668.270 ;
        RECT -27.470 1665.490 -26.290 1666.670 ;
        RECT -27.470 1487.090 -26.290 1488.270 ;
        RECT -27.470 1485.490 -26.290 1486.670 ;
        RECT -27.470 1307.090 -26.290 1308.270 ;
        RECT -27.470 1305.490 -26.290 1306.670 ;
        RECT -27.470 1127.090 -26.290 1128.270 ;
        RECT -27.470 1125.490 -26.290 1126.670 ;
        RECT -27.470 947.090 -26.290 948.270 ;
        RECT -27.470 945.490 -26.290 946.670 ;
        RECT -27.470 767.090 -26.290 768.270 ;
        RECT -27.470 765.490 -26.290 766.670 ;
        RECT -27.470 587.090 -26.290 588.270 ;
        RECT -27.470 585.490 -26.290 586.670 ;
        RECT -27.470 407.090 -26.290 408.270 ;
        RECT -27.470 405.490 -26.290 406.670 ;
        RECT -27.470 227.090 -26.290 228.270 ;
        RECT -27.470 225.490 -26.290 226.670 ;
        RECT -27.470 47.090 -26.290 48.270 ;
        RECT -27.470 45.490 -26.290 46.670 ;
        RECT -27.470 -21.310 -26.290 -20.130 ;
        RECT -27.470 -22.910 -26.290 -21.730 ;
        RECT 40.930 3541.410 42.110 3542.590 ;
        RECT 40.930 3539.810 42.110 3540.990 ;
        RECT 40.930 3467.090 42.110 3468.270 ;
        RECT 40.930 3465.490 42.110 3466.670 ;
        RECT 40.930 3287.090 42.110 3288.270 ;
        RECT 40.930 3285.490 42.110 3286.670 ;
        RECT 40.930 3107.090 42.110 3108.270 ;
        RECT 40.930 3105.490 42.110 3106.670 ;
        RECT 40.930 2927.090 42.110 2928.270 ;
        RECT 40.930 2925.490 42.110 2926.670 ;
        RECT 40.930 2747.090 42.110 2748.270 ;
        RECT 40.930 2745.490 42.110 2746.670 ;
        RECT 40.930 2567.090 42.110 2568.270 ;
        RECT 40.930 2565.490 42.110 2566.670 ;
        RECT 40.930 2387.090 42.110 2388.270 ;
        RECT 40.930 2385.490 42.110 2386.670 ;
        RECT 40.930 2207.090 42.110 2208.270 ;
        RECT 40.930 2205.490 42.110 2206.670 ;
        RECT 40.930 2027.090 42.110 2028.270 ;
        RECT 40.930 2025.490 42.110 2026.670 ;
        RECT 40.930 1847.090 42.110 1848.270 ;
        RECT 40.930 1845.490 42.110 1846.670 ;
        RECT 40.930 1667.090 42.110 1668.270 ;
        RECT 40.930 1665.490 42.110 1666.670 ;
        RECT 40.930 1487.090 42.110 1488.270 ;
        RECT 40.930 1485.490 42.110 1486.670 ;
        RECT 40.930 1307.090 42.110 1308.270 ;
        RECT 40.930 1305.490 42.110 1306.670 ;
        RECT 40.930 1127.090 42.110 1128.270 ;
        RECT 40.930 1125.490 42.110 1126.670 ;
        RECT 40.930 947.090 42.110 948.270 ;
        RECT 40.930 945.490 42.110 946.670 ;
        RECT 40.930 767.090 42.110 768.270 ;
        RECT 40.930 765.490 42.110 766.670 ;
        RECT 40.930 587.090 42.110 588.270 ;
        RECT 40.930 585.490 42.110 586.670 ;
        RECT 40.930 407.090 42.110 408.270 ;
        RECT 40.930 405.490 42.110 406.670 ;
        RECT 40.930 227.090 42.110 228.270 ;
        RECT 40.930 225.490 42.110 226.670 ;
        RECT 40.930 47.090 42.110 48.270 ;
        RECT 40.930 45.490 42.110 46.670 ;
        RECT 40.930 -21.310 42.110 -20.130 ;
        RECT 40.930 -22.910 42.110 -21.730 ;
        RECT 220.930 3541.410 222.110 3542.590 ;
        RECT 220.930 3539.810 222.110 3540.990 ;
        RECT 220.930 3467.090 222.110 3468.270 ;
        RECT 220.930 3465.490 222.110 3466.670 ;
        RECT 220.930 3287.090 222.110 3288.270 ;
        RECT 220.930 3285.490 222.110 3286.670 ;
        RECT 220.930 3107.090 222.110 3108.270 ;
        RECT 220.930 3105.490 222.110 3106.670 ;
        RECT 220.930 2927.090 222.110 2928.270 ;
        RECT 220.930 2925.490 222.110 2926.670 ;
        RECT 220.930 2747.090 222.110 2748.270 ;
        RECT 220.930 2745.490 222.110 2746.670 ;
        RECT 220.930 2567.090 222.110 2568.270 ;
        RECT 220.930 2565.490 222.110 2566.670 ;
        RECT 220.930 2387.090 222.110 2388.270 ;
        RECT 220.930 2385.490 222.110 2386.670 ;
        RECT 220.930 2207.090 222.110 2208.270 ;
        RECT 220.930 2205.490 222.110 2206.670 ;
        RECT 220.930 2027.090 222.110 2028.270 ;
        RECT 220.930 2025.490 222.110 2026.670 ;
        RECT 220.930 1847.090 222.110 1848.270 ;
        RECT 220.930 1845.490 222.110 1846.670 ;
        RECT 220.930 1667.090 222.110 1668.270 ;
        RECT 220.930 1665.490 222.110 1666.670 ;
        RECT 220.930 1487.090 222.110 1488.270 ;
        RECT 220.930 1485.490 222.110 1486.670 ;
        RECT 220.930 1307.090 222.110 1308.270 ;
        RECT 220.930 1305.490 222.110 1306.670 ;
        RECT 220.930 1127.090 222.110 1128.270 ;
        RECT 220.930 1125.490 222.110 1126.670 ;
        RECT 220.930 947.090 222.110 948.270 ;
        RECT 220.930 945.490 222.110 946.670 ;
        RECT 220.930 767.090 222.110 768.270 ;
        RECT 220.930 765.490 222.110 766.670 ;
        RECT 220.930 587.090 222.110 588.270 ;
        RECT 220.930 585.490 222.110 586.670 ;
        RECT 220.930 407.090 222.110 408.270 ;
        RECT 220.930 405.490 222.110 406.670 ;
        RECT 220.930 227.090 222.110 228.270 ;
        RECT 220.930 225.490 222.110 226.670 ;
        RECT 220.930 47.090 222.110 48.270 ;
        RECT 220.930 45.490 222.110 46.670 ;
        RECT 220.930 -21.310 222.110 -20.130 ;
        RECT 220.930 -22.910 222.110 -21.730 ;
        RECT 400.930 3541.410 402.110 3542.590 ;
        RECT 400.930 3539.810 402.110 3540.990 ;
        RECT 400.930 3467.090 402.110 3468.270 ;
        RECT 400.930 3465.490 402.110 3466.670 ;
        RECT 400.930 3287.090 402.110 3288.270 ;
        RECT 400.930 3285.490 402.110 3286.670 ;
        RECT 400.930 3107.090 402.110 3108.270 ;
        RECT 400.930 3105.490 402.110 3106.670 ;
        RECT 400.930 2927.090 402.110 2928.270 ;
        RECT 400.930 2925.490 402.110 2926.670 ;
        RECT 400.930 2747.090 402.110 2748.270 ;
        RECT 400.930 2745.490 402.110 2746.670 ;
        RECT 400.930 2567.090 402.110 2568.270 ;
        RECT 400.930 2565.490 402.110 2566.670 ;
        RECT 400.930 2387.090 402.110 2388.270 ;
        RECT 400.930 2385.490 402.110 2386.670 ;
        RECT 400.930 2207.090 402.110 2208.270 ;
        RECT 400.930 2205.490 402.110 2206.670 ;
        RECT 400.930 2027.090 402.110 2028.270 ;
        RECT 400.930 2025.490 402.110 2026.670 ;
        RECT 400.930 1847.090 402.110 1848.270 ;
        RECT 400.930 1845.490 402.110 1846.670 ;
        RECT 400.930 1667.090 402.110 1668.270 ;
        RECT 400.930 1665.490 402.110 1666.670 ;
        RECT 400.930 1487.090 402.110 1488.270 ;
        RECT 400.930 1485.490 402.110 1486.670 ;
        RECT 400.930 1307.090 402.110 1308.270 ;
        RECT 400.930 1305.490 402.110 1306.670 ;
        RECT 400.930 1127.090 402.110 1128.270 ;
        RECT 400.930 1125.490 402.110 1126.670 ;
        RECT 400.930 947.090 402.110 948.270 ;
        RECT 400.930 945.490 402.110 946.670 ;
        RECT 400.930 767.090 402.110 768.270 ;
        RECT 400.930 765.490 402.110 766.670 ;
        RECT 400.930 587.090 402.110 588.270 ;
        RECT 400.930 585.490 402.110 586.670 ;
        RECT 400.930 407.090 402.110 408.270 ;
        RECT 400.930 405.490 402.110 406.670 ;
        RECT 400.930 227.090 402.110 228.270 ;
        RECT 400.930 225.490 402.110 226.670 ;
        RECT 400.930 47.090 402.110 48.270 ;
        RECT 400.930 45.490 402.110 46.670 ;
        RECT 400.930 -21.310 402.110 -20.130 ;
        RECT 400.930 -22.910 402.110 -21.730 ;
        RECT 580.930 3541.410 582.110 3542.590 ;
        RECT 580.930 3539.810 582.110 3540.990 ;
        RECT 580.930 3467.090 582.110 3468.270 ;
        RECT 580.930 3465.490 582.110 3466.670 ;
        RECT 580.930 3287.090 582.110 3288.270 ;
        RECT 580.930 3285.490 582.110 3286.670 ;
        RECT 580.930 3107.090 582.110 3108.270 ;
        RECT 580.930 3105.490 582.110 3106.670 ;
        RECT 580.930 2927.090 582.110 2928.270 ;
        RECT 580.930 2925.490 582.110 2926.670 ;
        RECT 580.930 2747.090 582.110 2748.270 ;
        RECT 580.930 2745.490 582.110 2746.670 ;
        RECT 580.930 2567.090 582.110 2568.270 ;
        RECT 580.930 2565.490 582.110 2566.670 ;
        RECT 580.930 2387.090 582.110 2388.270 ;
        RECT 580.930 2385.490 582.110 2386.670 ;
        RECT 580.930 2207.090 582.110 2208.270 ;
        RECT 580.930 2205.490 582.110 2206.670 ;
        RECT 580.930 2027.090 582.110 2028.270 ;
        RECT 580.930 2025.490 582.110 2026.670 ;
        RECT 580.930 1847.090 582.110 1848.270 ;
        RECT 580.930 1845.490 582.110 1846.670 ;
        RECT 580.930 1667.090 582.110 1668.270 ;
        RECT 580.930 1665.490 582.110 1666.670 ;
        RECT 580.930 1487.090 582.110 1488.270 ;
        RECT 580.930 1485.490 582.110 1486.670 ;
        RECT 580.930 1307.090 582.110 1308.270 ;
        RECT 580.930 1305.490 582.110 1306.670 ;
        RECT 580.930 1127.090 582.110 1128.270 ;
        RECT 580.930 1125.490 582.110 1126.670 ;
        RECT 580.930 947.090 582.110 948.270 ;
        RECT 580.930 945.490 582.110 946.670 ;
        RECT 580.930 767.090 582.110 768.270 ;
        RECT 580.930 765.490 582.110 766.670 ;
        RECT 580.930 587.090 582.110 588.270 ;
        RECT 580.930 585.490 582.110 586.670 ;
        RECT 580.930 407.090 582.110 408.270 ;
        RECT 580.930 405.490 582.110 406.670 ;
        RECT 580.930 227.090 582.110 228.270 ;
        RECT 580.930 225.490 582.110 226.670 ;
        RECT 580.930 47.090 582.110 48.270 ;
        RECT 580.930 45.490 582.110 46.670 ;
        RECT 580.930 -21.310 582.110 -20.130 ;
        RECT 580.930 -22.910 582.110 -21.730 ;
        RECT 760.930 3541.410 762.110 3542.590 ;
        RECT 760.930 3539.810 762.110 3540.990 ;
        RECT 760.930 3467.090 762.110 3468.270 ;
        RECT 760.930 3465.490 762.110 3466.670 ;
        RECT 760.930 3287.090 762.110 3288.270 ;
        RECT 760.930 3285.490 762.110 3286.670 ;
        RECT 760.930 3107.090 762.110 3108.270 ;
        RECT 760.930 3105.490 762.110 3106.670 ;
        RECT 760.930 2927.090 762.110 2928.270 ;
        RECT 760.930 2925.490 762.110 2926.670 ;
        RECT 760.930 2747.090 762.110 2748.270 ;
        RECT 760.930 2745.490 762.110 2746.670 ;
        RECT 760.930 2567.090 762.110 2568.270 ;
        RECT 760.930 2565.490 762.110 2566.670 ;
        RECT 760.930 2387.090 762.110 2388.270 ;
        RECT 760.930 2385.490 762.110 2386.670 ;
        RECT 760.930 2207.090 762.110 2208.270 ;
        RECT 760.930 2205.490 762.110 2206.670 ;
        RECT 760.930 2027.090 762.110 2028.270 ;
        RECT 760.930 2025.490 762.110 2026.670 ;
        RECT 760.930 1847.090 762.110 1848.270 ;
        RECT 760.930 1845.490 762.110 1846.670 ;
        RECT 760.930 1667.090 762.110 1668.270 ;
        RECT 760.930 1665.490 762.110 1666.670 ;
        RECT 760.930 1487.090 762.110 1488.270 ;
        RECT 760.930 1485.490 762.110 1486.670 ;
        RECT 760.930 1307.090 762.110 1308.270 ;
        RECT 760.930 1305.490 762.110 1306.670 ;
        RECT 760.930 1127.090 762.110 1128.270 ;
        RECT 760.930 1125.490 762.110 1126.670 ;
        RECT 760.930 947.090 762.110 948.270 ;
        RECT 760.930 945.490 762.110 946.670 ;
        RECT 760.930 767.090 762.110 768.270 ;
        RECT 760.930 765.490 762.110 766.670 ;
        RECT 760.930 587.090 762.110 588.270 ;
        RECT 760.930 585.490 762.110 586.670 ;
        RECT 760.930 407.090 762.110 408.270 ;
        RECT 760.930 405.490 762.110 406.670 ;
        RECT 760.930 227.090 762.110 228.270 ;
        RECT 760.930 225.490 762.110 226.670 ;
        RECT 760.930 47.090 762.110 48.270 ;
        RECT 760.930 45.490 762.110 46.670 ;
        RECT 760.930 -21.310 762.110 -20.130 ;
        RECT 760.930 -22.910 762.110 -21.730 ;
        RECT 940.930 3541.410 942.110 3542.590 ;
        RECT 940.930 3539.810 942.110 3540.990 ;
        RECT 940.930 3467.090 942.110 3468.270 ;
        RECT 940.930 3465.490 942.110 3466.670 ;
        RECT 940.930 3287.090 942.110 3288.270 ;
        RECT 940.930 3285.490 942.110 3286.670 ;
        RECT 940.930 3107.090 942.110 3108.270 ;
        RECT 940.930 3105.490 942.110 3106.670 ;
        RECT 940.930 2927.090 942.110 2928.270 ;
        RECT 940.930 2925.490 942.110 2926.670 ;
        RECT 940.930 2747.090 942.110 2748.270 ;
        RECT 940.930 2745.490 942.110 2746.670 ;
        RECT 940.930 2567.090 942.110 2568.270 ;
        RECT 940.930 2565.490 942.110 2566.670 ;
        RECT 940.930 2387.090 942.110 2388.270 ;
        RECT 940.930 2385.490 942.110 2386.670 ;
        RECT 940.930 2207.090 942.110 2208.270 ;
        RECT 940.930 2205.490 942.110 2206.670 ;
        RECT 940.930 2027.090 942.110 2028.270 ;
        RECT 940.930 2025.490 942.110 2026.670 ;
        RECT 940.930 1847.090 942.110 1848.270 ;
        RECT 940.930 1845.490 942.110 1846.670 ;
        RECT 940.930 1667.090 942.110 1668.270 ;
        RECT 940.930 1665.490 942.110 1666.670 ;
        RECT 940.930 1487.090 942.110 1488.270 ;
        RECT 940.930 1485.490 942.110 1486.670 ;
        RECT 940.930 1307.090 942.110 1308.270 ;
        RECT 940.930 1305.490 942.110 1306.670 ;
        RECT 940.930 1127.090 942.110 1128.270 ;
        RECT 940.930 1125.490 942.110 1126.670 ;
        RECT 940.930 947.090 942.110 948.270 ;
        RECT 940.930 945.490 942.110 946.670 ;
        RECT 940.930 767.090 942.110 768.270 ;
        RECT 940.930 765.490 942.110 766.670 ;
        RECT 940.930 587.090 942.110 588.270 ;
        RECT 940.930 585.490 942.110 586.670 ;
        RECT 940.930 407.090 942.110 408.270 ;
        RECT 940.930 405.490 942.110 406.670 ;
        RECT 940.930 227.090 942.110 228.270 ;
        RECT 940.930 225.490 942.110 226.670 ;
        RECT 940.930 47.090 942.110 48.270 ;
        RECT 940.930 45.490 942.110 46.670 ;
        RECT 940.930 -21.310 942.110 -20.130 ;
        RECT 940.930 -22.910 942.110 -21.730 ;
        RECT 1120.930 3541.410 1122.110 3542.590 ;
        RECT 1120.930 3539.810 1122.110 3540.990 ;
        RECT 1120.930 3467.090 1122.110 3468.270 ;
        RECT 1120.930 3465.490 1122.110 3466.670 ;
        RECT 1120.930 3287.090 1122.110 3288.270 ;
        RECT 1120.930 3285.490 1122.110 3286.670 ;
        RECT 1120.930 3107.090 1122.110 3108.270 ;
        RECT 1120.930 3105.490 1122.110 3106.670 ;
        RECT 1120.930 2927.090 1122.110 2928.270 ;
        RECT 1120.930 2925.490 1122.110 2926.670 ;
        RECT 1120.930 2747.090 1122.110 2748.270 ;
        RECT 1120.930 2745.490 1122.110 2746.670 ;
        RECT 1120.930 2567.090 1122.110 2568.270 ;
        RECT 1120.930 2565.490 1122.110 2566.670 ;
        RECT 1120.930 2387.090 1122.110 2388.270 ;
        RECT 1120.930 2385.490 1122.110 2386.670 ;
        RECT 1120.930 2207.090 1122.110 2208.270 ;
        RECT 1120.930 2205.490 1122.110 2206.670 ;
        RECT 1120.930 2027.090 1122.110 2028.270 ;
        RECT 1120.930 2025.490 1122.110 2026.670 ;
        RECT 1120.930 1847.090 1122.110 1848.270 ;
        RECT 1120.930 1845.490 1122.110 1846.670 ;
        RECT 1120.930 1667.090 1122.110 1668.270 ;
        RECT 1120.930 1665.490 1122.110 1666.670 ;
        RECT 1120.930 1487.090 1122.110 1488.270 ;
        RECT 1120.930 1485.490 1122.110 1486.670 ;
        RECT 1120.930 1307.090 1122.110 1308.270 ;
        RECT 1120.930 1305.490 1122.110 1306.670 ;
        RECT 1120.930 1127.090 1122.110 1128.270 ;
        RECT 1120.930 1125.490 1122.110 1126.670 ;
        RECT 1120.930 947.090 1122.110 948.270 ;
        RECT 1120.930 945.490 1122.110 946.670 ;
        RECT 1120.930 767.090 1122.110 768.270 ;
        RECT 1120.930 765.490 1122.110 766.670 ;
        RECT 1120.930 587.090 1122.110 588.270 ;
        RECT 1120.930 585.490 1122.110 586.670 ;
        RECT 1120.930 407.090 1122.110 408.270 ;
        RECT 1120.930 405.490 1122.110 406.670 ;
        RECT 1120.930 227.090 1122.110 228.270 ;
        RECT 1120.930 225.490 1122.110 226.670 ;
        RECT 1120.930 47.090 1122.110 48.270 ;
        RECT 1120.930 45.490 1122.110 46.670 ;
        RECT 1120.930 -21.310 1122.110 -20.130 ;
        RECT 1120.930 -22.910 1122.110 -21.730 ;
        RECT 1300.930 3541.410 1302.110 3542.590 ;
        RECT 1300.930 3539.810 1302.110 3540.990 ;
        RECT 1300.930 3467.090 1302.110 3468.270 ;
        RECT 1300.930 3465.490 1302.110 3466.670 ;
        RECT 1300.930 3287.090 1302.110 3288.270 ;
        RECT 1300.930 3285.490 1302.110 3286.670 ;
        RECT 1300.930 3107.090 1302.110 3108.270 ;
        RECT 1300.930 3105.490 1302.110 3106.670 ;
        RECT 1300.930 2927.090 1302.110 2928.270 ;
        RECT 1300.930 2925.490 1302.110 2926.670 ;
        RECT 1300.930 2747.090 1302.110 2748.270 ;
        RECT 1300.930 2745.490 1302.110 2746.670 ;
        RECT 1300.930 2567.090 1302.110 2568.270 ;
        RECT 1300.930 2565.490 1302.110 2566.670 ;
        RECT 1300.930 2387.090 1302.110 2388.270 ;
        RECT 1300.930 2385.490 1302.110 2386.670 ;
        RECT 1300.930 2207.090 1302.110 2208.270 ;
        RECT 1300.930 2205.490 1302.110 2206.670 ;
        RECT 1300.930 2027.090 1302.110 2028.270 ;
        RECT 1300.930 2025.490 1302.110 2026.670 ;
        RECT 1300.930 1847.090 1302.110 1848.270 ;
        RECT 1300.930 1845.490 1302.110 1846.670 ;
        RECT 1300.930 1667.090 1302.110 1668.270 ;
        RECT 1300.930 1665.490 1302.110 1666.670 ;
        RECT 1300.930 1487.090 1302.110 1488.270 ;
        RECT 1300.930 1485.490 1302.110 1486.670 ;
        RECT 1300.930 1307.090 1302.110 1308.270 ;
        RECT 1300.930 1305.490 1302.110 1306.670 ;
        RECT 1300.930 1127.090 1302.110 1128.270 ;
        RECT 1300.930 1125.490 1302.110 1126.670 ;
        RECT 1300.930 947.090 1302.110 948.270 ;
        RECT 1300.930 945.490 1302.110 946.670 ;
        RECT 1300.930 767.090 1302.110 768.270 ;
        RECT 1300.930 765.490 1302.110 766.670 ;
        RECT 1300.930 587.090 1302.110 588.270 ;
        RECT 1300.930 585.490 1302.110 586.670 ;
        RECT 1300.930 407.090 1302.110 408.270 ;
        RECT 1300.930 405.490 1302.110 406.670 ;
        RECT 1300.930 227.090 1302.110 228.270 ;
        RECT 1300.930 225.490 1302.110 226.670 ;
        RECT 1300.930 47.090 1302.110 48.270 ;
        RECT 1300.930 45.490 1302.110 46.670 ;
        RECT 1300.930 -21.310 1302.110 -20.130 ;
        RECT 1300.930 -22.910 1302.110 -21.730 ;
        RECT 1480.930 3541.410 1482.110 3542.590 ;
        RECT 1480.930 3539.810 1482.110 3540.990 ;
        RECT 1480.930 3467.090 1482.110 3468.270 ;
        RECT 1480.930 3465.490 1482.110 3466.670 ;
        RECT 1480.930 3287.090 1482.110 3288.270 ;
        RECT 1480.930 3285.490 1482.110 3286.670 ;
        RECT 1480.930 3107.090 1482.110 3108.270 ;
        RECT 1480.930 3105.490 1482.110 3106.670 ;
        RECT 1480.930 2927.090 1482.110 2928.270 ;
        RECT 1480.930 2925.490 1482.110 2926.670 ;
        RECT 1480.930 2747.090 1482.110 2748.270 ;
        RECT 1480.930 2745.490 1482.110 2746.670 ;
        RECT 1480.930 2567.090 1482.110 2568.270 ;
        RECT 1480.930 2565.490 1482.110 2566.670 ;
        RECT 1480.930 2387.090 1482.110 2388.270 ;
        RECT 1480.930 2385.490 1482.110 2386.670 ;
        RECT 1480.930 2207.090 1482.110 2208.270 ;
        RECT 1480.930 2205.490 1482.110 2206.670 ;
        RECT 1480.930 2027.090 1482.110 2028.270 ;
        RECT 1480.930 2025.490 1482.110 2026.670 ;
        RECT 1480.930 1847.090 1482.110 1848.270 ;
        RECT 1480.930 1845.490 1482.110 1846.670 ;
        RECT 1480.930 1667.090 1482.110 1668.270 ;
        RECT 1480.930 1665.490 1482.110 1666.670 ;
        RECT 1480.930 1487.090 1482.110 1488.270 ;
        RECT 1480.930 1485.490 1482.110 1486.670 ;
        RECT 1480.930 1307.090 1482.110 1308.270 ;
        RECT 1480.930 1305.490 1482.110 1306.670 ;
        RECT 1480.930 1127.090 1482.110 1128.270 ;
        RECT 1480.930 1125.490 1482.110 1126.670 ;
        RECT 1480.930 947.090 1482.110 948.270 ;
        RECT 1480.930 945.490 1482.110 946.670 ;
        RECT 1480.930 767.090 1482.110 768.270 ;
        RECT 1480.930 765.490 1482.110 766.670 ;
        RECT 1480.930 587.090 1482.110 588.270 ;
        RECT 1480.930 585.490 1482.110 586.670 ;
        RECT 1480.930 407.090 1482.110 408.270 ;
        RECT 1480.930 405.490 1482.110 406.670 ;
        RECT 1480.930 227.090 1482.110 228.270 ;
        RECT 1480.930 225.490 1482.110 226.670 ;
        RECT 1480.930 47.090 1482.110 48.270 ;
        RECT 1480.930 45.490 1482.110 46.670 ;
        RECT 1480.930 -21.310 1482.110 -20.130 ;
        RECT 1480.930 -22.910 1482.110 -21.730 ;
        RECT 1660.930 3541.410 1662.110 3542.590 ;
        RECT 1660.930 3539.810 1662.110 3540.990 ;
        RECT 1660.930 3467.090 1662.110 3468.270 ;
        RECT 1660.930 3465.490 1662.110 3466.670 ;
        RECT 1660.930 3287.090 1662.110 3288.270 ;
        RECT 1660.930 3285.490 1662.110 3286.670 ;
        RECT 1660.930 3107.090 1662.110 3108.270 ;
        RECT 1660.930 3105.490 1662.110 3106.670 ;
        RECT 1660.930 2927.090 1662.110 2928.270 ;
        RECT 1660.930 2925.490 1662.110 2926.670 ;
        RECT 1660.930 2747.090 1662.110 2748.270 ;
        RECT 1660.930 2745.490 1662.110 2746.670 ;
        RECT 1660.930 2567.090 1662.110 2568.270 ;
        RECT 1660.930 2565.490 1662.110 2566.670 ;
        RECT 1660.930 2387.090 1662.110 2388.270 ;
        RECT 1660.930 2385.490 1662.110 2386.670 ;
        RECT 1660.930 2207.090 1662.110 2208.270 ;
        RECT 1660.930 2205.490 1662.110 2206.670 ;
        RECT 1660.930 2027.090 1662.110 2028.270 ;
        RECT 1660.930 2025.490 1662.110 2026.670 ;
        RECT 1660.930 1847.090 1662.110 1848.270 ;
        RECT 1660.930 1845.490 1662.110 1846.670 ;
        RECT 1660.930 1667.090 1662.110 1668.270 ;
        RECT 1660.930 1665.490 1662.110 1666.670 ;
        RECT 1660.930 1487.090 1662.110 1488.270 ;
        RECT 1660.930 1485.490 1662.110 1486.670 ;
        RECT 1660.930 1307.090 1662.110 1308.270 ;
        RECT 1660.930 1305.490 1662.110 1306.670 ;
        RECT 1660.930 1127.090 1662.110 1128.270 ;
        RECT 1660.930 1125.490 1662.110 1126.670 ;
        RECT 1660.930 947.090 1662.110 948.270 ;
        RECT 1660.930 945.490 1662.110 946.670 ;
        RECT 1660.930 767.090 1662.110 768.270 ;
        RECT 1660.930 765.490 1662.110 766.670 ;
        RECT 1660.930 587.090 1662.110 588.270 ;
        RECT 1660.930 585.490 1662.110 586.670 ;
        RECT 1660.930 407.090 1662.110 408.270 ;
        RECT 1660.930 405.490 1662.110 406.670 ;
        RECT 1660.930 227.090 1662.110 228.270 ;
        RECT 1660.930 225.490 1662.110 226.670 ;
        RECT 1660.930 47.090 1662.110 48.270 ;
        RECT 1660.930 45.490 1662.110 46.670 ;
        RECT 1660.930 -21.310 1662.110 -20.130 ;
        RECT 1660.930 -22.910 1662.110 -21.730 ;
        RECT 1840.930 3541.410 1842.110 3542.590 ;
        RECT 1840.930 3539.810 1842.110 3540.990 ;
        RECT 1840.930 3467.090 1842.110 3468.270 ;
        RECT 1840.930 3465.490 1842.110 3466.670 ;
        RECT 1840.930 3287.090 1842.110 3288.270 ;
        RECT 1840.930 3285.490 1842.110 3286.670 ;
        RECT 1840.930 3107.090 1842.110 3108.270 ;
        RECT 1840.930 3105.490 1842.110 3106.670 ;
        RECT 1840.930 2927.090 1842.110 2928.270 ;
        RECT 1840.930 2925.490 1842.110 2926.670 ;
        RECT 1840.930 2747.090 1842.110 2748.270 ;
        RECT 1840.930 2745.490 1842.110 2746.670 ;
        RECT 1840.930 2567.090 1842.110 2568.270 ;
        RECT 1840.930 2565.490 1842.110 2566.670 ;
        RECT 1840.930 2387.090 1842.110 2388.270 ;
        RECT 1840.930 2385.490 1842.110 2386.670 ;
        RECT 1840.930 2207.090 1842.110 2208.270 ;
        RECT 1840.930 2205.490 1842.110 2206.670 ;
        RECT 1840.930 2027.090 1842.110 2028.270 ;
        RECT 1840.930 2025.490 1842.110 2026.670 ;
        RECT 1840.930 1847.090 1842.110 1848.270 ;
        RECT 1840.930 1845.490 1842.110 1846.670 ;
        RECT 1840.930 1667.090 1842.110 1668.270 ;
        RECT 1840.930 1665.490 1842.110 1666.670 ;
        RECT 1840.930 1487.090 1842.110 1488.270 ;
        RECT 1840.930 1485.490 1842.110 1486.670 ;
        RECT 1840.930 1307.090 1842.110 1308.270 ;
        RECT 1840.930 1305.490 1842.110 1306.670 ;
        RECT 1840.930 1127.090 1842.110 1128.270 ;
        RECT 1840.930 1125.490 1842.110 1126.670 ;
        RECT 1840.930 947.090 1842.110 948.270 ;
        RECT 1840.930 945.490 1842.110 946.670 ;
        RECT 1840.930 767.090 1842.110 768.270 ;
        RECT 1840.930 765.490 1842.110 766.670 ;
        RECT 1840.930 587.090 1842.110 588.270 ;
        RECT 1840.930 585.490 1842.110 586.670 ;
        RECT 1840.930 407.090 1842.110 408.270 ;
        RECT 1840.930 405.490 1842.110 406.670 ;
        RECT 1840.930 227.090 1842.110 228.270 ;
        RECT 1840.930 225.490 1842.110 226.670 ;
        RECT 1840.930 47.090 1842.110 48.270 ;
        RECT 1840.930 45.490 1842.110 46.670 ;
        RECT 1840.930 -21.310 1842.110 -20.130 ;
        RECT 1840.930 -22.910 1842.110 -21.730 ;
        RECT 2020.930 3541.410 2022.110 3542.590 ;
        RECT 2020.930 3539.810 2022.110 3540.990 ;
        RECT 2020.930 3467.090 2022.110 3468.270 ;
        RECT 2020.930 3465.490 2022.110 3466.670 ;
        RECT 2020.930 3287.090 2022.110 3288.270 ;
        RECT 2020.930 3285.490 2022.110 3286.670 ;
        RECT 2020.930 3107.090 2022.110 3108.270 ;
        RECT 2020.930 3105.490 2022.110 3106.670 ;
        RECT 2020.930 2927.090 2022.110 2928.270 ;
        RECT 2020.930 2925.490 2022.110 2926.670 ;
        RECT 2020.930 2747.090 2022.110 2748.270 ;
        RECT 2020.930 2745.490 2022.110 2746.670 ;
        RECT 2020.930 2567.090 2022.110 2568.270 ;
        RECT 2020.930 2565.490 2022.110 2566.670 ;
        RECT 2020.930 2387.090 2022.110 2388.270 ;
        RECT 2020.930 2385.490 2022.110 2386.670 ;
        RECT 2020.930 2207.090 2022.110 2208.270 ;
        RECT 2020.930 2205.490 2022.110 2206.670 ;
        RECT 2020.930 2027.090 2022.110 2028.270 ;
        RECT 2020.930 2025.490 2022.110 2026.670 ;
        RECT 2020.930 1847.090 2022.110 1848.270 ;
        RECT 2020.930 1845.490 2022.110 1846.670 ;
        RECT 2020.930 1667.090 2022.110 1668.270 ;
        RECT 2020.930 1665.490 2022.110 1666.670 ;
        RECT 2020.930 1487.090 2022.110 1488.270 ;
        RECT 2020.930 1485.490 2022.110 1486.670 ;
        RECT 2020.930 1307.090 2022.110 1308.270 ;
        RECT 2020.930 1305.490 2022.110 1306.670 ;
        RECT 2020.930 1127.090 2022.110 1128.270 ;
        RECT 2020.930 1125.490 2022.110 1126.670 ;
        RECT 2020.930 947.090 2022.110 948.270 ;
        RECT 2020.930 945.490 2022.110 946.670 ;
        RECT 2020.930 767.090 2022.110 768.270 ;
        RECT 2020.930 765.490 2022.110 766.670 ;
        RECT 2020.930 587.090 2022.110 588.270 ;
        RECT 2020.930 585.490 2022.110 586.670 ;
        RECT 2020.930 407.090 2022.110 408.270 ;
        RECT 2020.930 405.490 2022.110 406.670 ;
        RECT 2020.930 227.090 2022.110 228.270 ;
        RECT 2020.930 225.490 2022.110 226.670 ;
        RECT 2020.930 47.090 2022.110 48.270 ;
        RECT 2020.930 45.490 2022.110 46.670 ;
        RECT 2020.930 -21.310 2022.110 -20.130 ;
        RECT 2020.930 -22.910 2022.110 -21.730 ;
        RECT 2200.930 3541.410 2202.110 3542.590 ;
        RECT 2200.930 3539.810 2202.110 3540.990 ;
        RECT 2200.930 3467.090 2202.110 3468.270 ;
        RECT 2200.930 3465.490 2202.110 3466.670 ;
        RECT 2200.930 3287.090 2202.110 3288.270 ;
        RECT 2200.930 3285.490 2202.110 3286.670 ;
        RECT 2200.930 3107.090 2202.110 3108.270 ;
        RECT 2200.930 3105.490 2202.110 3106.670 ;
        RECT 2200.930 2927.090 2202.110 2928.270 ;
        RECT 2200.930 2925.490 2202.110 2926.670 ;
        RECT 2200.930 2747.090 2202.110 2748.270 ;
        RECT 2200.930 2745.490 2202.110 2746.670 ;
        RECT 2200.930 2567.090 2202.110 2568.270 ;
        RECT 2200.930 2565.490 2202.110 2566.670 ;
        RECT 2200.930 2387.090 2202.110 2388.270 ;
        RECT 2200.930 2385.490 2202.110 2386.670 ;
        RECT 2200.930 2207.090 2202.110 2208.270 ;
        RECT 2200.930 2205.490 2202.110 2206.670 ;
        RECT 2200.930 2027.090 2202.110 2028.270 ;
        RECT 2200.930 2025.490 2202.110 2026.670 ;
        RECT 2200.930 1847.090 2202.110 1848.270 ;
        RECT 2200.930 1845.490 2202.110 1846.670 ;
        RECT 2200.930 1667.090 2202.110 1668.270 ;
        RECT 2200.930 1665.490 2202.110 1666.670 ;
        RECT 2200.930 1487.090 2202.110 1488.270 ;
        RECT 2200.930 1485.490 2202.110 1486.670 ;
        RECT 2200.930 1307.090 2202.110 1308.270 ;
        RECT 2200.930 1305.490 2202.110 1306.670 ;
        RECT 2200.930 1127.090 2202.110 1128.270 ;
        RECT 2200.930 1125.490 2202.110 1126.670 ;
        RECT 2200.930 947.090 2202.110 948.270 ;
        RECT 2200.930 945.490 2202.110 946.670 ;
        RECT 2200.930 767.090 2202.110 768.270 ;
        RECT 2200.930 765.490 2202.110 766.670 ;
        RECT 2200.930 587.090 2202.110 588.270 ;
        RECT 2200.930 585.490 2202.110 586.670 ;
        RECT 2200.930 407.090 2202.110 408.270 ;
        RECT 2200.930 405.490 2202.110 406.670 ;
        RECT 2200.930 227.090 2202.110 228.270 ;
        RECT 2200.930 225.490 2202.110 226.670 ;
        RECT 2200.930 47.090 2202.110 48.270 ;
        RECT 2200.930 45.490 2202.110 46.670 ;
        RECT 2200.930 -21.310 2202.110 -20.130 ;
        RECT 2200.930 -22.910 2202.110 -21.730 ;
        RECT 2380.930 3541.410 2382.110 3542.590 ;
        RECT 2380.930 3539.810 2382.110 3540.990 ;
        RECT 2380.930 3467.090 2382.110 3468.270 ;
        RECT 2380.930 3465.490 2382.110 3466.670 ;
        RECT 2380.930 3287.090 2382.110 3288.270 ;
        RECT 2380.930 3285.490 2382.110 3286.670 ;
        RECT 2380.930 3107.090 2382.110 3108.270 ;
        RECT 2380.930 3105.490 2382.110 3106.670 ;
        RECT 2380.930 2927.090 2382.110 2928.270 ;
        RECT 2380.930 2925.490 2382.110 2926.670 ;
        RECT 2380.930 2747.090 2382.110 2748.270 ;
        RECT 2380.930 2745.490 2382.110 2746.670 ;
        RECT 2380.930 2567.090 2382.110 2568.270 ;
        RECT 2380.930 2565.490 2382.110 2566.670 ;
        RECT 2380.930 2387.090 2382.110 2388.270 ;
        RECT 2380.930 2385.490 2382.110 2386.670 ;
        RECT 2380.930 2207.090 2382.110 2208.270 ;
        RECT 2380.930 2205.490 2382.110 2206.670 ;
        RECT 2380.930 2027.090 2382.110 2028.270 ;
        RECT 2380.930 2025.490 2382.110 2026.670 ;
        RECT 2380.930 1847.090 2382.110 1848.270 ;
        RECT 2380.930 1845.490 2382.110 1846.670 ;
        RECT 2380.930 1667.090 2382.110 1668.270 ;
        RECT 2380.930 1665.490 2382.110 1666.670 ;
        RECT 2380.930 1487.090 2382.110 1488.270 ;
        RECT 2380.930 1485.490 2382.110 1486.670 ;
        RECT 2380.930 1307.090 2382.110 1308.270 ;
        RECT 2380.930 1305.490 2382.110 1306.670 ;
        RECT 2380.930 1127.090 2382.110 1128.270 ;
        RECT 2380.930 1125.490 2382.110 1126.670 ;
        RECT 2380.930 947.090 2382.110 948.270 ;
        RECT 2380.930 945.490 2382.110 946.670 ;
        RECT 2380.930 767.090 2382.110 768.270 ;
        RECT 2380.930 765.490 2382.110 766.670 ;
        RECT 2380.930 587.090 2382.110 588.270 ;
        RECT 2380.930 585.490 2382.110 586.670 ;
        RECT 2380.930 407.090 2382.110 408.270 ;
        RECT 2380.930 405.490 2382.110 406.670 ;
        RECT 2380.930 227.090 2382.110 228.270 ;
        RECT 2380.930 225.490 2382.110 226.670 ;
        RECT 2380.930 47.090 2382.110 48.270 ;
        RECT 2380.930 45.490 2382.110 46.670 ;
        RECT 2380.930 -21.310 2382.110 -20.130 ;
        RECT 2380.930 -22.910 2382.110 -21.730 ;
        RECT 2560.930 3541.410 2562.110 3542.590 ;
        RECT 2560.930 3539.810 2562.110 3540.990 ;
        RECT 2560.930 3467.090 2562.110 3468.270 ;
        RECT 2560.930 3465.490 2562.110 3466.670 ;
        RECT 2560.930 3287.090 2562.110 3288.270 ;
        RECT 2560.930 3285.490 2562.110 3286.670 ;
        RECT 2560.930 3107.090 2562.110 3108.270 ;
        RECT 2560.930 3105.490 2562.110 3106.670 ;
        RECT 2560.930 2927.090 2562.110 2928.270 ;
        RECT 2560.930 2925.490 2562.110 2926.670 ;
        RECT 2560.930 2747.090 2562.110 2748.270 ;
        RECT 2560.930 2745.490 2562.110 2746.670 ;
        RECT 2560.930 2567.090 2562.110 2568.270 ;
        RECT 2560.930 2565.490 2562.110 2566.670 ;
        RECT 2560.930 2387.090 2562.110 2388.270 ;
        RECT 2560.930 2385.490 2562.110 2386.670 ;
        RECT 2560.930 2207.090 2562.110 2208.270 ;
        RECT 2560.930 2205.490 2562.110 2206.670 ;
        RECT 2560.930 2027.090 2562.110 2028.270 ;
        RECT 2560.930 2025.490 2562.110 2026.670 ;
        RECT 2560.930 1847.090 2562.110 1848.270 ;
        RECT 2560.930 1845.490 2562.110 1846.670 ;
        RECT 2560.930 1667.090 2562.110 1668.270 ;
        RECT 2560.930 1665.490 2562.110 1666.670 ;
        RECT 2560.930 1487.090 2562.110 1488.270 ;
        RECT 2560.930 1485.490 2562.110 1486.670 ;
        RECT 2560.930 1307.090 2562.110 1308.270 ;
        RECT 2560.930 1305.490 2562.110 1306.670 ;
        RECT 2560.930 1127.090 2562.110 1128.270 ;
        RECT 2560.930 1125.490 2562.110 1126.670 ;
        RECT 2560.930 947.090 2562.110 948.270 ;
        RECT 2560.930 945.490 2562.110 946.670 ;
        RECT 2560.930 767.090 2562.110 768.270 ;
        RECT 2560.930 765.490 2562.110 766.670 ;
        RECT 2560.930 587.090 2562.110 588.270 ;
        RECT 2560.930 585.490 2562.110 586.670 ;
        RECT 2560.930 407.090 2562.110 408.270 ;
        RECT 2560.930 405.490 2562.110 406.670 ;
        RECT 2560.930 227.090 2562.110 228.270 ;
        RECT 2560.930 225.490 2562.110 226.670 ;
        RECT 2560.930 47.090 2562.110 48.270 ;
        RECT 2560.930 45.490 2562.110 46.670 ;
        RECT 2560.930 -21.310 2562.110 -20.130 ;
        RECT 2560.930 -22.910 2562.110 -21.730 ;
        RECT 2740.930 3541.410 2742.110 3542.590 ;
        RECT 2740.930 3539.810 2742.110 3540.990 ;
        RECT 2740.930 3467.090 2742.110 3468.270 ;
        RECT 2740.930 3465.490 2742.110 3466.670 ;
        RECT 2740.930 3287.090 2742.110 3288.270 ;
        RECT 2740.930 3285.490 2742.110 3286.670 ;
        RECT 2740.930 3107.090 2742.110 3108.270 ;
        RECT 2740.930 3105.490 2742.110 3106.670 ;
        RECT 2740.930 2927.090 2742.110 2928.270 ;
        RECT 2740.930 2925.490 2742.110 2926.670 ;
        RECT 2740.930 2747.090 2742.110 2748.270 ;
        RECT 2740.930 2745.490 2742.110 2746.670 ;
        RECT 2740.930 2567.090 2742.110 2568.270 ;
        RECT 2740.930 2565.490 2742.110 2566.670 ;
        RECT 2740.930 2387.090 2742.110 2388.270 ;
        RECT 2740.930 2385.490 2742.110 2386.670 ;
        RECT 2740.930 2207.090 2742.110 2208.270 ;
        RECT 2740.930 2205.490 2742.110 2206.670 ;
        RECT 2740.930 2027.090 2742.110 2028.270 ;
        RECT 2740.930 2025.490 2742.110 2026.670 ;
        RECT 2740.930 1847.090 2742.110 1848.270 ;
        RECT 2740.930 1845.490 2742.110 1846.670 ;
        RECT 2740.930 1667.090 2742.110 1668.270 ;
        RECT 2740.930 1665.490 2742.110 1666.670 ;
        RECT 2740.930 1487.090 2742.110 1488.270 ;
        RECT 2740.930 1485.490 2742.110 1486.670 ;
        RECT 2740.930 1307.090 2742.110 1308.270 ;
        RECT 2740.930 1305.490 2742.110 1306.670 ;
        RECT 2740.930 1127.090 2742.110 1128.270 ;
        RECT 2740.930 1125.490 2742.110 1126.670 ;
        RECT 2740.930 947.090 2742.110 948.270 ;
        RECT 2740.930 945.490 2742.110 946.670 ;
        RECT 2740.930 767.090 2742.110 768.270 ;
        RECT 2740.930 765.490 2742.110 766.670 ;
        RECT 2740.930 587.090 2742.110 588.270 ;
        RECT 2740.930 585.490 2742.110 586.670 ;
        RECT 2740.930 407.090 2742.110 408.270 ;
        RECT 2740.930 405.490 2742.110 406.670 ;
        RECT 2740.930 227.090 2742.110 228.270 ;
        RECT 2740.930 225.490 2742.110 226.670 ;
        RECT 2740.930 47.090 2742.110 48.270 ;
        RECT 2740.930 45.490 2742.110 46.670 ;
        RECT 2740.930 -21.310 2742.110 -20.130 ;
        RECT 2740.930 -22.910 2742.110 -21.730 ;
        RECT 2945.910 3541.410 2947.090 3542.590 ;
        RECT 2945.910 3539.810 2947.090 3540.990 ;
        RECT 2945.910 3467.090 2947.090 3468.270 ;
        RECT 2945.910 3465.490 2947.090 3466.670 ;
        RECT 2945.910 3287.090 2947.090 3288.270 ;
        RECT 2945.910 3285.490 2947.090 3286.670 ;
        RECT 2945.910 3107.090 2947.090 3108.270 ;
        RECT 2945.910 3105.490 2947.090 3106.670 ;
        RECT 2945.910 2927.090 2947.090 2928.270 ;
        RECT 2945.910 2925.490 2947.090 2926.670 ;
        RECT 2945.910 2747.090 2947.090 2748.270 ;
        RECT 2945.910 2745.490 2947.090 2746.670 ;
        RECT 2945.910 2567.090 2947.090 2568.270 ;
        RECT 2945.910 2565.490 2947.090 2566.670 ;
        RECT 2945.910 2387.090 2947.090 2388.270 ;
        RECT 2945.910 2385.490 2947.090 2386.670 ;
        RECT 2945.910 2207.090 2947.090 2208.270 ;
        RECT 2945.910 2205.490 2947.090 2206.670 ;
        RECT 2945.910 2027.090 2947.090 2028.270 ;
        RECT 2945.910 2025.490 2947.090 2026.670 ;
        RECT 2945.910 1847.090 2947.090 1848.270 ;
        RECT 2945.910 1845.490 2947.090 1846.670 ;
        RECT 2945.910 1667.090 2947.090 1668.270 ;
        RECT 2945.910 1665.490 2947.090 1666.670 ;
        RECT 2945.910 1487.090 2947.090 1488.270 ;
        RECT 2945.910 1485.490 2947.090 1486.670 ;
        RECT 2945.910 1307.090 2947.090 1308.270 ;
        RECT 2945.910 1305.490 2947.090 1306.670 ;
        RECT 2945.910 1127.090 2947.090 1128.270 ;
        RECT 2945.910 1125.490 2947.090 1126.670 ;
        RECT 2945.910 947.090 2947.090 948.270 ;
        RECT 2945.910 945.490 2947.090 946.670 ;
        RECT 2945.910 767.090 2947.090 768.270 ;
        RECT 2945.910 765.490 2947.090 766.670 ;
        RECT 2945.910 587.090 2947.090 588.270 ;
        RECT 2945.910 585.490 2947.090 586.670 ;
        RECT 2945.910 407.090 2947.090 408.270 ;
        RECT 2945.910 405.490 2947.090 406.670 ;
        RECT 2945.910 227.090 2947.090 228.270 ;
        RECT 2945.910 225.490 2947.090 226.670 ;
        RECT 2945.910 47.090 2947.090 48.270 ;
        RECT 2945.910 45.490 2947.090 46.670 ;
        RECT 2945.910 -21.310 2947.090 -20.130 ;
        RECT 2945.910 -22.910 2947.090 -21.730 ;
      LAYER met5 ;
        RECT -28.380 3542.700 -25.380 3542.710 ;
        RECT 40.020 3542.700 43.020 3542.710 ;
        RECT 220.020 3542.700 223.020 3542.710 ;
        RECT 400.020 3542.700 403.020 3542.710 ;
        RECT 580.020 3542.700 583.020 3542.710 ;
        RECT 760.020 3542.700 763.020 3542.710 ;
        RECT 940.020 3542.700 943.020 3542.710 ;
        RECT 1120.020 3542.700 1123.020 3542.710 ;
        RECT 1300.020 3542.700 1303.020 3542.710 ;
        RECT 1480.020 3542.700 1483.020 3542.710 ;
        RECT 1660.020 3542.700 1663.020 3542.710 ;
        RECT 1840.020 3542.700 1843.020 3542.710 ;
        RECT 2020.020 3542.700 2023.020 3542.710 ;
        RECT 2200.020 3542.700 2203.020 3542.710 ;
        RECT 2380.020 3542.700 2383.020 3542.710 ;
        RECT 2560.020 3542.700 2563.020 3542.710 ;
        RECT 2740.020 3542.700 2743.020 3542.710 ;
        RECT 2945.000 3542.700 2948.000 3542.710 ;
        RECT -28.380 3539.700 2948.000 3542.700 ;
        RECT -28.380 3539.690 -25.380 3539.700 ;
        RECT 40.020 3539.690 43.020 3539.700 ;
        RECT 220.020 3539.690 223.020 3539.700 ;
        RECT 400.020 3539.690 403.020 3539.700 ;
        RECT 580.020 3539.690 583.020 3539.700 ;
        RECT 760.020 3539.690 763.020 3539.700 ;
        RECT 940.020 3539.690 943.020 3539.700 ;
        RECT 1120.020 3539.690 1123.020 3539.700 ;
        RECT 1300.020 3539.690 1303.020 3539.700 ;
        RECT 1480.020 3539.690 1483.020 3539.700 ;
        RECT 1660.020 3539.690 1663.020 3539.700 ;
        RECT 1840.020 3539.690 1843.020 3539.700 ;
        RECT 2020.020 3539.690 2023.020 3539.700 ;
        RECT 2200.020 3539.690 2203.020 3539.700 ;
        RECT 2380.020 3539.690 2383.020 3539.700 ;
        RECT 2560.020 3539.690 2563.020 3539.700 ;
        RECT 2740.020 3539.690 2743.020 3539.700 ;
        RECT 2945.000 3539.690 2948.000 3539.700 ;
        RECT -28.380 3468.380 -25.380 3468.390 ;
        RECT 40.020 3468.380 43.020 3468.390 ;
        RECT 220.020 3468.380 223.020 3468.390 ;
        RECT 400.020 3468.380 403.020 3468.390 ;
        RECT 580.020 3468.380 583.020 3468.390 ;
        RECT 760.020 3468.380 763.020 3468.390 ;
        RECT 940.020 3468.380 943.020 3468.390 ;
        RECT 1120.020 3468.380 1123.020 3468.390 ;
        RECT 1300.020 3468.380 1303.020 3468.390 ;
        RECT 1480.020 3468.380 1483.020 3468.390 ;
        RECT 1660.020 3468.380 1663.020 3468.390 ;
        RECT 1840.020 3468.380 1843.020 3468.390 ;
        RECT 2020.020 3468.380 2023.020 3468.390 ;
        RECT 2200.020 3468.380 2203.020 3468.390 ;
        RECT 2380.020 3468.380 2383.020 3468.390 ;
        RECT 2560.020 3468.380 2563.020 3468.390 ;
        RECT 2740.020 3468.380 2743.020 3468.390 ;
        RECT 2945.000 3468.380 2948.000 3468.390 ;
        RECT -32.980 3465.380 2952.600 3468.380 ;
        RECT -28.380 3465.370 -25.380 3465.380 ;
        RECT 40.020 3465.370 43.020 3465.380 ;
        RECT 220.020 3465.370 223.020 3465.380 ;
        RECT 400.020 3465.370 403.020 3465.380 ;
        RECT 580.020 3465.370 583.020 3465.380 ;
        RECT 760.020 3465.370 763.020 3465.380 ;
        RECT 940.020 3465.370 943.020 3465.380 ;
        RECT 1120.020 3465.370 1123.020 3465.380 ;
        RECT 1300.020 3465.370 1303.020 3465.380 ;
        RECT 1480.020 3465.370 1483.020 3465.380 ;
        RECT 1660.020 3465.370 1663.020 3465.380 ;
        RECT 1840.020 3465.370 1843.020 3465.380 ;
        RECT 2020.020 3465.370 2023.020 3465.380 ;
        RECT 2200.020 3465.370 2203.020 3465.380 ;
        RECT 2380.020 3465.370 2383.020 3465.380 ;
        RECT 2560.020 3465.370 2563.020 3465.380 ;
        RECT 2740.020 3465.370 2743.020 3465.380 ;
        RECT 2945.000 3465.370 2948.000 3465.380 ;
        RECT -28.380 3288.380 -25.380 3288.390 ;
        RECT 40.020 3288.380 43.020 3288.390 ;
        RECT 220.020 3288.380 223.020 3288.390 ;
        RECT 400.020 3288.380 403.020 3288.390 ;
        RECT 580.020 3288.380 583.020 3288.390 ;
        RECT 760.020 3288.380 763.020 3288.390 ;
        RECT 940.020 3288.380 943.020 3288.390 ;
        RECT 1120.020 3288.380 1123.020 3288.390 ;
        RECT 1300.020 3288.380 1303.020 3288.390 ;
        RECT 1480.020 3288.380 1483.020 3288.390 ;
        RECT 1660.020 3288.380 1663.020 3288.390 ;
        RECT 1840.020 3288.380 1843.020 3288.390 ;
        RECT 2020.020 3288.380 2023.020 3288.390 ;
        RECT 2200.020 3288.380 2203.020 3288.390 ;
        RECT 2380.020 3288.380 2383.020 3288.390 ;
        RECT 2560.020 3288.380 2563.020 3288.390 ;
        RECT 2740.020 3288.380 2743.020 3288.390 ;
        RECT 2945.000 3288.380 2948.000 3288.390 ;
        RECT -32.980 3285.380 2952.600 3288.380 ;
        RECT -28.380 3285.370 -25.380 3285.380 ;
        RECT 40.020 3285.370 43.020 3285.380 ;
        RECT 220.020 3285.370 223.020 3285.380 ;
        RECT 400.020 3285.370 403.020 3285.380 ;
        RECT 580.020 3285.370 583.020 3285.380 ;
        RECT 760.020 3285.370 763.020 3285.380 ;
        RECT 940.020 3285.370 943.020 3285.380 ;
        RECT 1120.020 3285.370 1123.020 3285.380 ;
        RECT 1300.020 3285.370 1303.020 3285.380 ;
        RECT 1480.020 3285.370 1483.020 3285.380 ;
        RECT 1660.020 3285.370 1663.020 3285.380 ;
        RECT 1840.020 3285.370 1843.020 3285.380 ;
        RECT 2020.020 3285.370 2023.020 3285.380 ;
        RECT 2200.020 3285.370 2203.020 3285.380 ;
        RECT 2380.020 3285.370 2383.020 3285.380 ;
        RECT 2560.020 3285.370 2563.020 3285.380 ;
        RECT 2740.020 3285.370 2743.020 3285.380 ;
        RECT 2945.000 3285.370 2948.000 3285.380 ;
        RECT -28.380 3108.380 -25.380 3108.390 ;
        RECT 40.020 3108.380 43.020 3108.390 ;
        RECT 220.020 3108.380 223.020 3108.390 ;
        RECT 400.020 3108.380 403.020 3108.390 ;
        RECT 580.020 3108.380 583.020 3108.390 ;
        RECT 760.020 3108.380 763.020 3108.390 ;
        RECT 940.020 3108.380 943.020 3108.390 ;
        RECT 1120.020 3108.380 1123.020 3108.390 ;
        RECT 1300.020 3108.380 1303.020 3108.390 ;
        RECT 1480.020 3108.380 1483.020 3108.390 ;
        RECT 1660.020 3108.380 1663.020 3108.390 ;
        RECT 1840.020 3108.380 1843.020 3108.390 ;
        RECT 2020.020 3108.380 2023.020 3108.390 ;
        RECT 2200.020 3108.380 2203.020 3108.390 ;
        RECT 2380.020 3108.380 2383.020 3108.390 ;
        RECT 2560.020 3108.380 2563.020 3108.390 ;
        RECT 2740.020 3108.380 2743.020 3108.390 ;
        RECT 2945.000 3108.380 2948.000 3108.390 ;
        RECT -32.980 3105.380 2952.600 3108.380 ;
        RECT -28.380 3105.370 -25.380 3105.380 ;
        RECT 40.020 3105.370 43.020 3105.380 ;
        RECT 220.020 3105.370 223.020 3105.380 ;
        RECT 400.020 3105.370 403.020 3105.380 ;
        RECT 580.020 3105.370 583.020 3105.380 ;
        RECT 760.020 3105.370 763.020 3105.380 ;
        RECT 940.020 3105.370 943.020 3105.380 ;
        RECT 1120.020 3105.370 1123.020 3105.380 ;
        RECT 1300.020 3105.370 1303.020 3105.380 ;
        RECT 1480.020 3105.370 1483.020 3105.380 ;
        RECT 1660.020 3105.370 1663.020 3105.380 ;
        RECT 1840.020 3105.370 1843.020 3105.380 ;
        RECT 2020.020 3105.370 2023.020 3105.380 ;
        RECT 2200.020 3105.370 2203.020 3105.380 ;
        RECT 2380.020 3105.370 2383.020 3105.380 ;
        RECT 2560.020 3105.370 2563.020 3105.380 ;
        RECT 2740.020 3105.370 2743.020 3105.380 ;
        RECT 2945.000 3105.370 2948.000 3105.380 ;
        RECT -28.380 2928.380 -25.380 2928.390 ;
        RECT 40.020 2928.380 43.020 2928.390 ;
        RECT 220.020 2928.380 223.020 2928.390 ;
        RECT 400.020 2928.380 403.020 2928.390 ;
        RECT 580.020 2928.380 583.020 2928.390 ;
        RECT 760.020 2928.380 763.020 2928.390 ;
        RECT 940.020 2928.380 943.020 2928.390 ;
        RECT 1120.020 2928.380 1123.020 2928.390 ;
        RECT 1300.020 2928.380 1303.020 2928.390 ;
        RECT 1480.020 2928.380 1483.020 2928.390 ;
        RECT 1660.020 2928.380 1663.020 2928.390 ;
        RECT 1840.020 2928.380 1843.020 2928.390 ;
        RECT 2020.020 2928.380 2023.020 2928.390 ;
        RECT 2200.020 2928.380 2203.020 2928.390 ;
        RECT 2380.020 2928.380 2383.020 2928.390 ;
        RECT 2560.020 2928.380 2563.020 2928.390 ;
        RECT 2740.020 2928.380 2743.020 2928.390 ;
        RECT 2945.000 2928.380 2948.000 2928.390 ;
        RECT -32.980 2925.380 2952.600 2928.380 ;
        RECT -28.380 2925.370 -25.380 2925.380 ;
        RECT 40.020 2925.370 43.020 2925.380 ;
        RECT 220.020 2925.370 223.020 2925.380 ;
        RECT 400.020 2925.370 403.020 2925.380 ;
        RECT 580.020 2925.370 583.020 2925.380 ;
        RECT 760.020 2925.370 763.020 2925.380 ;
        RECT 940.020 2925.370 943.020 2925.380 ;
        RECT 1120.020 2925.370 1123.020 2925.380 ;
        RECT 1300.020 2925.370 1303.020 2925.380 ;
        RECT 1480.020 2925.370 1483.020 2925.380 ;
        RECT 1660.020 2925.370 1663.020 2925.380 ;
        RECT 1840.020 2925.370 1843.020 2925.380 ;
        RECT 2020.020 2925.370 2023.020 2925.380 ;
        RECT 2200.020 2925.370 2203.020 2925.380 ;
        RECT 2380.020 2925.370 2383.020 2925.380 ;
        RECT 2560.020 2925.370 2563.020 2925.380 ;
        RECT 2740.020 2925.370 2743.020 2925.380 ;
        RECT 2945.000 2925.370 2948.000 2925.380 ;
        RECT -28.380 2748.380 -25.380 2748.390 ;
        RECT 40.020 2748.380 43.020 2748.390 ;
        RECT 220.020 2748.380 223.020 2748.390 ;
        RECT 400.020 2748.380 403.020 2748.390 ;
        RECT 580.020 2748.380 583.020 2748.390 ;
        RECT 760.020 2748.380 763.020 2748.390 ;
        RECT 940.020 2748.380 943.020 2748.390 ;
        RECT 1120.020 2748.380 1123.020 2748.390 ;
        RECT 1300.020 2748.380 1303.020 2748.390 ;
        RECT 1480.020 2748.380 1483.020 2748.390 ;
        RECT 1660.020 2748.380 1663.020 2748.390 ;
        RECT 1840.020 2748.380 1843.020 2748.390 ;
        RECT 2020.020 2748.380 2023.020 2748.390 ;
        RECT 2200.020 2748.380 2203.020 2748.390 ;
        RECT 2380.020 2748.380 2383.020 2748.390 ;
        RECT 2560.020 2748.380 2563.020 2748.390 ;
        RECT 2740.020 2748.380 2743.020 2748.390 ;
        RECT 2945.000 2748.380 2948.000 2748.390 ;
        RECT -32.980 2745.380 2952.600 2748.380 ;
        RECT -28.380 2745.370 -25.380 2745.380 ;
        RECT 40.020 2745.370 43.020 2745.380 ;
        RECT 220.020 2745.370 223.020 2745.380 ;
        RECT 400.020 2745.370 403.020 2745.380 ;
        RECT 580.020 2745.370 583.020 2745.380 ;
        RECT 760.020 2745.370 763.020 2745.380 ;
        RECT 940.020 2745.370 943.020 2745.380 ;
        RECT 1120.020 2745.370 1123.020 2745.380 ;
        RECT 1300.020 2745.370 1303.020 2745.380 ;
        RECT 1480.020 2745.370 1483.020 2745.380 ;
        RECT 1660.020 2745.370 1663.020 2745.380 ;
        RECT 1840.020 2745.370 1843.020 2745.380 ;
        RECT 2020.020 2745.370 2023.020 2745.380 ;
        RECT 2200.020 2745.370 2203.020 2745.380 ;
        RECT 2380.020 2745.370 2383.020 2745.380 ;
        RECT 2560.020 2745.370 2563.020 2745.380 ;
        RECT 2740.020 2745.370 2743.020 2745.380 ;
        RECT 2945.000 2745.370 2948.000 2745.380 ;
        RECT -28.380 2568.380 -25.380 2568.390 ;
        RECT 40.020 2568.380 43.020 2568.390 ;
        RECT 220.020 2568.380 223.020 2568.390 ;
        RECT 400.020 2568.380 403.020 2568.390 ;
        RECT 580.020 2568.380 583.020 2568.390 ;
        RECT 760.020 2568.380 763.020 2568.390 ;
        RECT 940.020 2568.380 943.020 2568.390 ;
        RECT 1120.020 2568.380 1123.020 2568.390 ;
        RECT 1300.020 2568.380 1303.020 2568.390 ;
        RECT 1480.020 2568.380 1483.020 2568.390 ;
        RECT 1660.020 2568.380 1663.020 2568.390 ;
        RECT 1840.020 2568.380 1843.020 2568.390 ;
        RECT 2020.020 2568.380 2023.020 2568.390 ;
        RECT 2200.020 2568.380 2203.020 2568.390 ;
        RECT 2380.020 2568.380 2383.020 2568.390 ;
        RECT 2560.020 2568.380 2563.020 2568.390 ;
        RECT 2740.020 2568.380 2743.020 2568.390 ;
        RECT 2945.000 2568.380 2948.000 2568.390 ;
        RECT -32.980 2565.380 2952.600 2568.380 ;
        RECT -28.380 2565.370 -25.380 2565.380 ;
        RECT 40.020 2565.370 43.020 2565.380 ;
        RECT 220.020 2565.370 223.020 2565.380 ;
        RECT 400.020 2565.370 403.020 2565.380 ;
        RECT 580.020 2565.370 583.020 2565.380 ;
        RECT 760.020 2565.370 763.020 2565.380 ;
        RECT 940.020 2565.370 943.020 2565.380 ;
        RECT 1120.020 2565.370 1123.020 2565.380 ;
        RECT 1300.020 2565.370 1303.020 2565.380 ;
        RECT 1480.020 2565.370 1483.020 2565.380 ;
        RECT 1660.020 2565.370 1663.020 2565.380 ;
        RECT 1840.020 2565.370 1843.020 2565.380 ;
        RECT 2020.020 2565.370 2023.020 2565.380 ;
        RECT 2200.020 2565.370 2203.020 2565.380 ;
        RECT 2380.020 2565.370 2383.020 2565.380 ;
        RECT 2560.020 2565.370 2563.020 2565.380 ;
        RECT 2740.020 2565.370 2743.020 2565.380 ;
        RECT 2945.000 2565.370 2948.000 2565.380 ;
        RECT -28.380 2388.380 -25.380 2388.390 ;
        RECT 40.020 2388.380 43.020 2388.390 ;
        RECT 220.020 2388.380 223.020 2388.390 ;
        RECT 400.020 2388.380 403.020 2388.390 ;
        RECT 580.020 2388.380 583.020 2388.390 ;
        RECT 760.020 2388.380 763.020 2388.390 ;
        RECT 940.020 2388.380 943.020 2388.390 ;
        RECT 1120.020 2388.380 1123.020 2388.390 ;
        RECT 1300.020 2388.380 1303.020 2388.390 ;
        RECT 1480.020 2388.380 1483.020 2388.390 ;
        RECT 1660.020 2388.380 1663.020 2388.390 ;
        RECT 1840.020 2388.380 1843.020 2388.390 ;
        RECT 2020.020 2388.380 2023.020 2388.390 ;
        RECT 2200.020 2388.380 2203.020 2388.390 ;
        RECT 2380.020 2388.380 2383.020 2388.390 ;
        RECT 2560.020 2388.380 2563.020 2388.390 ;
        RECT 2740.020 2388.380 2743.020 2388.390 ;
        RECT 2945.000 2388.380 2948.000 2388.390 ;
        RECT -32.980 2385.380 2952.600 2388.380 ;
        RECT -28.380 2385.370 -25.380 2385.380 ;
        RECT 40.020 2385.370 43.020 2385.380 ;
        RECT 220.020 2385.370 223.020 2385.380 ;
        RECT 400.020 2385.370 403.020 2385.380 ;
        RECT 580.020 2385.370 583.020 2385.380 ;
        RECT 760.020 2385.370 763.020 2385.380 ;
        RECT 940.020 2385.370 943.020 2385.380 ;
        RECT 1120.020 2385.370 1123.020 2385.380 ;
        RECT 1300.020 2385.370 1303.020 2385.380 ;
        RECT 1480.020 2385.370 1483.020 2385.380 ;
        RECT 1660.020 2385.370 1663.020 2385.380 ;
        RECT 1840.020 2385.370 1843.020 2385.380 ;
        RECT 2020.020 2385.370 2023.020 2385.380 ;
        RECT 2200.020 2385.370 2203.020 2385.380 ;
        RECT 2380.020 2385.370 2383.020 2385.380 ;
        RECT 2560.020 2385.370 2563.020 2385.380 ;
        RECT 2740.020 2385.370 2743.020 2385.380 ;
        RECT 2945.000 2385.370 2948.000 2385.380 ;
        RECT -28.380 2208.380 -25.380 2208.390 ;
        RECT 40.020 2208.380 43.020 2208.390 ;
        RECT 220.020 2208.380 223.020 2208.390 ;
        RECT 400.020 2208.380 403.020 2208.390 ;
        RECT 580.020 2208.380 583.020 2208.390 ;
        RECT 760.020 2208.380 763.020 2208.390 ;
        RECT 940.020 2208.380 943.020 2208.390 ;
        RECT 1120.020 2208.380 1123.020 2208.390 ;
        RECT 1300.020 2208.380 1303.020 2208.390 ;
        RECT 1480.020 2208.380 1483.020 2208.390 ;
        RECT 1660.020 2208.380 1663.020 2208.390 ;
        RECT 1840.020 2208.380 1843.020 2208.390 ;
        RECT 2020.020 2208.380 2023.020 2208.390 ;
        RECT 2200.020 2208.380 2203.020 2208.390 ;
        RECT 2380.020 2208.380 2383.020 2208.390 ;
        RECT 2560.020 2208.380 2563.020 2208.390 ;
        RECT 2740.020 2208.380 2743.020 2208.390 ;
        RECT 2945.000 2208.380 2948.000 2208.390 ;
        RECT -32.980 2205.380 2952.600 2208.380 ;
        RECT -28.380 2205.370 -25.380 2205.380 ;
        RECT 40.020 2205.370 43.020 2205.380 ;
        RECT 220.020 2205.370 223.020 2205.380 ;
        RECT 400.020 2205.370 403.020 2205.380 ;
        RECT 580.020 2205.370 583.020 2205.380 ;
        RECT 760.020 2205.370 763.020 2205.380 ;
        RECT 940.020 2205.370 943.020 2205.380 ;
        RECT 1120.020 2205.370 1123.020 2205.380 ;
        RECT 1300.020 2205.370 1303.020 2205.380 ;
        RECT 1480.020 2205.370 1483.020 2205.380 ;
        RECT 1660.020 2205.370 1663.020 2205.380 ;
        RECT 1840.020 2205.370 1843.020 2205.380 ;
        RECT 2020.020 2205.370 2023.020 2205.380 ;
        RECT 2200.020 2205.370 2203.020 2205.380 ;
        RECT 2380.020 2205.370 2383.020 2205.380 ;
        RECT 2560.020 2205.370 2563.020 2205.380 ;
        RECT 2740.020 2205.370 2743.020 2205.380 ;
        RECT 2945.000 2205.370 2948.000 2205.380 ;
        RECT -28.380 2028.380 -25.380 2028.390 ;
        RECT 40.020 2028.380 43.020 2028.390 ;
        RECT 220.020 2028.380 223.020 2028.390 ;
        RECT 400.020 2028.380 403.020 2028.390 ;
        RECT 580.020 2028.380 583.020 2028.390 ;
        RECT 760.020 2028.380 763.020 2028.390 ;
        RECT 940.020 2028.380 943.020 2028.390 ;
        RECT 1120.020 2028.380 1123.020 2028.390 ;
        RECT 1300.020 2028.380 1303.020 2028.390 ;
        RECT 1480.020 2028.380 1483.020 2028.390 ;
        RECT 1660.020 2028.380 1663.020 2028.390 ;
        RECT 1840.020 2028.380 1843.020 2028.390 ;
        RECT 2020.020 2028.380 2023.020 2028.390 ;
        RECT 2200.020 2028.380 2203.020 2028.390 ;
        RECT 2380.020 2028.380 2383.020 2028.390 ;
        RECT 2560.020 2028.380 2563.020 2028.390 ;
        RECT 2740.020 2028.380 2743.020 2028.390 ;
        RECT 2945.000 2028.380 2948.000 2028.390 ;
        RECT -32.980 2025.380 2952.600 2028.380 ;
        RECT -28.380 2025.370 -25.380 2025.380 ;
        RECT 40.020 2025.370 43.020 2025.380 ;
        RECT 220.020 2025.370 223.020 2025.380 ;
        RECT 400.020 2025.370 403.020 2025.380 ;
        RECT 580.020 2025.370 583.020 2025.380 ;
        RECT 760.020 2025.370 763.020 2025.380 ;
        RECT 940.020 2025.370 943.020 2025.380 ;
        RECT 1120.020 2025.370 1123.020 2025.380 ;
        RECT 1300.020 2025.370 1303.020 2025.380 ;
        RECT 1480.020 2025.370 1483.020 2025.380 ;
        RECT 1660.020 2025.370 1663.020 2025.380 ;
        RECT 1840.020 2025.370 1843.020 2025.380 ;
        RECT 2020.020 2025.370 2023.020 2025.380 ;
        RECT 2200.020 2025.370 2203.020 2025.380 ;
        RECT 2380.020 2025.370 2383.020 2025.380 ;
        RECT 2560.020 2025.370 2563.020 2025.380 ;
        RECT 2740.020 2025.370 2743.020 2025.380 ;
        RECT 2945.000 2025.370 2948.000 2025.380 ;
        RECT -28.380 1848.380 -25.380 1848.390 ;
        RECT 40.020 1848.380 43.020 1848.390 ;
        RECT 220.020 1848.380 223.020 1848.390 ;
        RECT 400.020 1848.380 403.020 1848.390 ;
        RECT 580.020 1848.380 583.020 1848.390 ;
        RECT 760.020 1848.380 763.020 1848.390 ;
        RECT 940.020 1848.380 943.020 1848.390 ;
        RECT 1120.020 1848.380 1123.020 1848.390 ;
        RECT 1300.020 1848.380 1303.020 1848.390 ;
        RECT 1480.020 1848.380 1483.020 1848.390 ;
        RECT 1660.020 1848.380 1663.020 1848.390 ;
        RECT 1840.020 1848.380 1843.020 1848.390 ;
        RECT 2020.020 1848.380 2023.020 1848.390 ;
        RECT 2200.020 1848.380 2203.020 1848.390 ;
        RECT 2380.020 1848.380 2383.020 1848.390 ;
        RECT 2560.020 1848.380 2563.020 1848.390 ;
        RECT 2740.020 1848.380 2743.020 1848.390 ;
        RECT 2945.000 1848.380 2948.000 1848.390 ;
        RECT -32.980 1845.380 2952.600 1848.380 ;
        RECT -28.380 1845.370 -25.380 1845.380 ;
        RECT 40.020 1845.370 43.020 1845.380 ;
        RECT 220.020 1845.370 223.020 1845.380 ;
        RECT 400.020 1845.370 403.020 1845.380 ;
        RECT 580.020 1845.370 583.020 1845.380 ;
        RECT 760.020 1845.370 763.020 1845.380 ;
        RECT 940.020 1845.370 943.020 1845.380 ;
        RECT 1120.020 1845.370 1123.020 1845.380 ;
        RECT 1300.020 1845.370 1303.020 1845.380 ;
        RECT 1480.020 1845.370 1483.020 1845.380 ;
        RECT 1660.020 1845.370 1663.020 1845.380 ;
        RECT 1840.020 1845.370 1843.020 1845.380 ;
        RECT 2020.020 1845.370 2023.020 1845.380 ;
        RECT 2200.020 1845.370 2203.020 1845.380 ;
        RECT 2380.020 1845.370 2383.020 1845.380 ;
        RECT 2560.020 1845.370 2563.020 1845.380 ;
        RECT 2740.020 1845.370 2743.020 1845.380 ;
        RECT 2945.000 1845.370 2948.000 1845.380 ;
        RECT -28.380 1668.380 -25.380 1668.390 ;
        RECT 40.020 1668.380 43.020 1668.390 ;
        RECT 220.020 1668.380 223.020 1668.390 ;
        RECT 400.020 1668.380 403.020 1668.390 ;
        RECT 580.020 1668.380 583.020 1668.390 ;
        RECT 760.020 1668.380 763.020 1668.390 ;
        RECT 940.020 1668.380 943.020 1668.390 ;
        RECT 1120.020 1668.380 1123.020 1668.390 ;
        RECT 1300.020 1668.380 1303.020 1668.390 ;
        RECT 1480.020 1668.380 1483.020 1668.390 ;
        RECT 1660.020 1668.380 1663.020 1668.390 ;
        RECT 1840.020 1668.380 1843.020 1668.390 ;
        RECT 2020.020 1668.380 2023.020 1668.390 ;
        RECT 2200.020 1668.380 2203.020 1668.390 ;
        RECT 2380.020 1668.380 2383.020 1668.390 ;
        RECT 2560.020 1668.380 2563.020 1668.390 ;
        RECT 2740.020 1668.380 2743.020 1668.390 ;
        RECT 2945.000 1668.380 2948.000 1668.390 ;
        RECT -32.980 1665.380 2952.600 1668.380 ;
        RECT -28.380 1665.370 -25.380 1665.380 ;
        RECT 40.020 1665.370 43.020 1665.380 ;
        RECT 220.020 1665.370 223.020 1665.380 ;
        RECT 400.020 1665.370 403.020 1665.380 ;
        RECT 580.020 1665.370 583.020 1665.380 ;
        RECT 760.020 1665.370 763.020 1665.380 ;
        RECT 940.020 1665.370 943.020 1665.380 ;
        RECT 1120.020 1665.370 1123.020 1665.380 ;
        RECT 1300.020 1665.370 1303.020 1665.380 ;
        RECT 1480.020 1665.370 1483.020 1665.380 ;
        RECT 1660.020 1665.370 1663.020 1665.380 ;
        RECT 1840.020 1665.370 1843.020 1665.380 ;
        RECT 2020.020 1665.370 2023.020 1665.380 ;
        RECT 2200.020 1665.370 2203.020 1665.380 ;
        RECT 2380.020 1665.370 2383.020 1665.380 ;
        RECT 2560.020 1665.370 2563.020 1665.380 ;
        RECT 2740.020 1665.370 2743.020 1665.380 ;
        RECT 2945.000 1665.370 2948.000 1665.380 ;
        RECT -28.380 1488.380 -25.380 1488.390 ;
        RECT 40.020 1488.380 43.020 1488.390 ;
        RECT 220.020 1488.380 223.020 1488.390 ;
        RECT 400.020 1488.380 403.020 1488.390 ;
        RECT 580.020 1488.380 583.020 1488.390 ;
        RECT 760.020 1488.380 763.020 1488.390 ;
        RECT 940.020 1488.380 943.020 1488.390 ;
        RECT 1120.020 1488.380 1123.020 1488.390 ;
        RECT 1300.020 1488.380 1303.020 1488.390 ;
        RECT 1480.020 1488.380 1483.020 1488.390 ;
        RECT 1660.020 1488.380 1663.020 1488.390 ;
        RECT 1840.020 1488.380 1843.020 1488.390 ;
        RECT 2020.020 1488.380 2023.020 1488.390 ;
        RECT 2200.020 1488.380 2203.020 1488.390 ;
        RECT 2380.020 1488.380 2383.020 1488.390 ;
        RECT 2560.020 1488.380 2563.020 1488.390 ;
        RECT 2740.020 1488.380 2743.020 1488.390 ;
        RECT 2945.000 1488.380 2948.000 1488.390 ;
        RECT -32.980 1485.380 2952.600 1488.380 ;
        RECT -28.380 1485.370 -25.380 1485.380 ;
        RECT 40.020 1485.370 43.020 1485.380 ;
        RECT 220.020 1485.370 223.020 1485.380 ;
        RECT 400.020 1485.370 403.020 1485.380 ;
        RECT 580.020 1485.370 583.020 1485.380 ;
        RECT 760.020 1485.370 763.020 1485.380 ;
        RECT 940.020 1485.370 943.020 1485.380 ;
        RECT 1120.020 1485.370 1123.020 1485.380 ;
        RECT 1300.020 1485.370 1303.020 1485.380 ;
        RECT 1480.020 1485.370 1483.020 1485.380 ;
        RECT 1660.020 1485.370 1663.020 1485.380 ;
        RECT 1840.020 1485.370 1843.020 1485.380 ;
        RECT 2020.020 1485.370 2023.020 1485.380 ;
        RECT 2200.020 1485.370 2203.020 1485.380 ;
        RECT 2380.020 1485.370 2383.020 1485.380 ;
        RECT 2560.020 1485.370 2563.020 1485.380 ;
        RECT 2740.020 1485.370 2743.020 1485.380 ;
        RECT 2945.000 1485.370 2948.000 1485.380 ;
        RECT -28.380 1308.380 -25.380 1308.390 ;
        RECT 40.020 1308.380 43.020 1308.390 ;
        RECT 220.020 1308.380 223.020 1308.390 ;
        RECT 400.020 1308.380 403.020 1308.390 ;
        RECT 580.020 1308.380 583.020 1308.390 ;
        RECT 760.020 1308.380 763.020 1308.390 ;
        RECT 940.020 1308.380 943.020 1308.390 ;
        RECT 1120.020 1308.380 1123.020 1308.390 ;
        RECT 1300.020 1308.380 1303.020 1308.390 ;
        RECT 1480.020 1308.380 1483.020 1308.390 ;
        RECT 1660.020 1308.380 1663.020 1308.390 ;
        RECT 1840.020 1308.380 1843.020 1308.390 ;
        RECT 2020.020 1308.380 2023.020 1308.390 ;
        RECT 2200.020 1308.380 2203.020 1308.390 ;
        RECT 2380.020 1308.380 2383.020 1308.390 ;
        RECT 2560.020 1308.380 2563.020 1308.390 ;
        RECT 2740.020 1308.380 2743.020 1308.390 ;
        RECT 2945.000 1308.380 2948.000 1308.390 ;
        RECT -32.980 1305.380 2952.600 1308.380 ;
        RECT -28.380 1305.370 -25.380 1305.380 ;
        RECT 40.020 1305.370 43.020 1305.380 ;
        RECT 220.020 1305.370 223.020 1305.380 ;
        RECT 400.020 1305.370 403.020 1305.380 ;
        RECT 580.020 1305.370 583.020 1305.380 ;
        RECT 760.020 1305.370 763.020 1305.380 ;
        RECT 940.020 1305.370 943.020 1305.380 ;
        RECT 1120.020 1305.370 1123.020 1305.380 ;
        RECT 1300.020 1305.370 1303.020 1305.380 ;
        RECT 1480.020 1305.370 1483.020 1305.380 ;
        RECT 1660.020 1305.370 1663.020 1305.380 ;
        RECT 1840.020 1305.370 1843.020 1305.380 ;
        RECT 2020.020 1305.370 2023.020 1305.380 ;
        RECT 2200.020 1305.370 2203.020 1305.380 ;
        RECT 2380.020 1305.370 2383.020 1305.380 ;
        RECT 2560.020 1305.370 2563.020 1305.380 ;
        RECT 2740.020 1305.370 2743.020 1305.380 ;
        RECT 2945.000 1305.370 2948.000 1305.380 ;
        RECT -28.380 1128.380 -25.380 1128.390 ;
        RECT 40.020 1128.380 43.020 1128.390 ;
        RECT 220.020 1128.380 223.020 1128.390 ;
        RECT 400.020 1128.380 403.020 1128.390 ;
        RECT 580.020 1128.380 583.020 1128.390 ;
        RECT 760.020 1128.380 763.020 1128.390 ;
        RECT 940.020 1128.380 943.020 1128.390 ;
        RECT 1120.020 1128.380 1123.020 1128.390 ;
        RECT 1300.020 1128.380 1303.020 1128.390 ;
        RECT 1480.020 1128.380 1483.020 1128.390 ;
        RECT 1660.020 1128.380 1663.020 1128.390 ;
        RECT 1840.020 1128.380 1843.020 1128.390 ;
        RECT 2020.020 1128.380 2023.020 1128.390 ;
        RECT 2200.020 1128.380 2203.020 1128.390 ;
        RECT 2380.020 1128.380 2383.020 1128.390 ;
        RECT 2560.020 1128.380 2563.020 1128.390 ;
        RECT 2740.020 1128.380 2743.020 1128.390 ;
        RECT 2945.000 1128.380 2948.000 1128.390 ;
        RECT -32.980 1125.380 2952.600 1128.380 ;
        RECT -28.380 1125.370 -25.380 1125.380 ;
        RECT 40.020 1125.370 43.020 1125.380 ;
        RECT 220.020 1125.370 223.020 1125.380 ;
        RECT 400.020 1125.370 403.020 1125.380 ;
        RECT 580.020 1125.370 583.020 1125.380 ;
        RECT 760.020 1125.370 763.020 1125.380 ;
        RECT 940.020 1125.370 943.020 1125.380 ;
        RECT 1120.020 1125.370 1123.020 1125.380 ;
        RECT 1300.020 1125.370 1303.020 1125.380 ;
        RECT 1480.020 1125.370 1483.020 1125.380 ;
        RECT 1660.020 1125.370 1663.020 1125.380 ;
        RECT 1840.020 1125.370 1843.020 1125.380 ;
        RECT 2020.020 1125.370 2023.020 1125.380 ;
        RECT 2200.020 1125.370 2203.020 1125.380 ;
        RECT 2380.020 1125.370 2383.020 1125.380 ;
        RECT 2560.020 1125.370 2563.020 1125.380 ;
        RECT 2740.020 1125.370 2743.020 1125.380 ;
        RECT 2945.000 1125.370 2948.000 1125.380 ;
        RECT -28.380 948.380 -25.380 948.390 ;
        RECT 40.020 948.380 43.020 948.390 ;
        RECT 220.020 948.380 223.020 948.390 ;
        RECT 400.020 948.380 403.020 948.390 ;
        RECT 580.020 948.380 583.020 948.390 ;
        RECT 760.020 948.380 763.020 948.390 ;
        RECT 940.020 948.380 943.020 948.390 ;
        RECT 1120.020 948.380 1123.020 948.390 ;
        RECT 1300.020 948.380 1303.020 948.390 ;
        RECT 1480.020 948.380 1483.020 948.390 ;
        RECT 1660.020 948.380 1663.020 948.390 ;
        RECT 1840.020 948.380 1843.020 948.390 ;
        RECT 2020.020 948.380 2023.020 948.390 ;
        RECT 2200.020 948.380 2203.020 948.390 ;
        RECT 2380.020 948.380 2383.020 948.390 ;
        RECT 2560.020 948.380 2563.020 948.390 ;
        RECT 2740.020 948.380 2743.020 948.390 ;
        RECT 2945.000 948.380 2948.000 948.390 ;
        RECT -32.980 945.380 2952.600 948.380 ;
        RECT -28.380 945.370 -25.380 945.380 ;
        RECT 40.020 945.370 43.020 945.380 ;
        RECT 220.020 945.370 223.020 945.380 ;
        RECT 400.020 945.370 403.020 945.380 ;
        RECT 580.020 945.370 583.020 945.380 ;
        RECT 760.020 945.370 763.020 945.380 ;
        RECT 940.020 945.370 943.020 945.380 ;
        RECT 1120.020 945.370 1123.020 945.380 ;
        RECT 1300.020 945.370 1303.020 945.380 ;
        RECT 1480.020 945.370 1483.020 945.380 ;
        RECT 1660.020 945.370 1663.020 945.380 ;
        RECT 1840.020 945.370 1843.020 945.380 ;
        RECT 2020.020 945.370 2023.020 945.380 ;
        RECT 2200.020 945.370 2203.020 945.380 ;
        RECT 2380.020 945.370 2383.020 945.380 ;
        RECT 2560.020 945.370 2563.020 945.380 ;
        RECT 2740.020 945.370 2743.020 945.380 ;
        RECT 2945.000 945.370 2948.000 945.380 ;
        RECT -28.380 768.380 -25.380 768.390 ;
        RECT 40.020 768.380 43.020 768.390 ;
        RECT 220.020 768.380 223.020 768.390 ;
        RECT 400.020 768.380 403.020 768.390 ;
        RECT 580.020 768.380 583.020 768.390 ;
        RECT 760.020 768.380 763.020 768.390 ;
        RECT 940.020 768.380 943.020 768.390 ;
        RECT 1120.020 768.380 1123.020 768.390 ;
        RECT 1300.020 768.380 1303.020 768.390 ;
        RECT 1480.020 768.380 1483.020 768.390 ;
        RECT 1660.020 768.380 1663.020 768.390 ;
        RECT 1840.020 768.380 1843.020 768.390 ;
        RECT 2020.020 768.380 2023.020 768.390 ;
        RECT 2200.020 768.380 2203.020 768.390 ;
        RECT 2380.020 768.380 2383.020 768.390 ;
        RECT 2560.020 768.380 2563.020 768.390 ;
        RECT 2740.020 768.380 2743.020 768.390 ;
        RECT 2945.000 768.380 2948.000 768.390 ;
        RECT -32.980 765.380 2952.600 768.380 ;
        RECT -28.380 765.370 -25.380 765.380 ;
        RECT 40.020 765.370 43.020 765.380 ;
        RECT 220.020 765.370 223.020 765.380 ;
        RECT 400.020 765.370 403.020 765.380 ;
        RECT 580.020 765.370 583.020 765.380 ;
        RECT 760.020 765.370 763.020 765.380 ;
        RECT 940.020 765.370 943.020 765.380 ;
        RECT 1120.020 765.370 1123.020 765.380 ;
        RECT 1300.020 765.370 1303.020 765.380 ;
        RECT 1480.020 765.370 1483.020 765.380 ;
        RECT 1660.020 765.370 1663.020 765.380 ;
        RECT 1840.020 765.370 1843.020 765.380 ;
        RECT 2020.020 765.370 2023.020 765.380 ;
        RECT 2200.020 765.370 2203.020 765.380 ;
        RECT 2380.020 765.370 2383.020 765.380 ;
        RECT 2560.020 765.370 2563.020 765.380 ;
        RECT 2740.020 765.370 2743.020 765.380 ;
        RECT 2945.000 765.370 2948.000 765.380 ;
        RECT -28.380 588.380 -25.380 588.390 ;
        RECT 40.020 588.380 43.020 588.390 ;
        RECT 220.020 588.380 223.020 588.390 ;
        RECT 400.020 588.380 403.020 588.390 ;
        RECT 580.020 588.380 583.020 588.390 ;
        RECT 760.020 588.380 763.020 588.390 ;
        RECT 940.020 588.380 943.020 588.390 ;
        RECT 1120.020 588.380 1123.020 588.390 ;
        RECT 1300.020 588.380 1303.020 588.390 ;
        RECT 1480.020 588.380 1483.020 588.390 ;
        RECT 1660.020 588.380 1663.020 588.390 ;
        RECT 1840.020 588.380 1843.020 588.390 ;
        RECT 2020.020 588.380 2023.020 588.390 ;
        RECT 2200.020 588.380 2203.020 588.390 ;
        RECT 2380.020 588.380 2383.020 588.390 ;
        RECT 2560.020 588.380 2563.020 588.390 ;
        RECT 2740.020 588.380 2743.020 588.390 ;
        RECT 2945.000 588.380 2948.000 588.390 ;
        RECT -32.980 585.380 2952.600 588.380 ;
        RECT -28.380 585.370 -25.380 585.380 ;
        RECT 40.020 585.370 43.020 585.380 ;
        RECT 220.020 585.370 223.020 585.380 ;
        RECT 400.020 585.370 403.020 585.380 ;
        RECT 580.020 585.370 583.020 585.380 ;
        RECT 760.020 585.370 763.020 585.380 ;
        RECT 940.020 585.370 943.020 585.380 ;
        RECT 1120.020 585.370 1123.020 585.380 ;
        RECT 1300.020 585.370 1303.020 585.380 ;
        RECT 1480.020 585.370 1483.020 585.380 ;
        RECT 1660.020 585.370 1663.020 585.380 ;
        RECT 1840.020 585.370 1843.020 585.380 ;
        RECT 2020.020 585.370 2023.020 585.380 ;
        RECT 2200.020 585.370 2203.020 585.380 ;
        RECT 2380.020 585.370 2383.020 585.380 ;
        RECT 2560.020 585.370 2563.020 585.380 ;
        RECT 2740.020 585.370 2743.020 585.380 ;
        RECT 2945.000 585.370 2948.000 585.380 ;
        RECT -28.380 408.380 -25.380 408.390 ;
        RECT 40.020 408.380 43.020 408.390 ;
        RECT 220.020 408.380 223.020 408.390 ;
        RECT 400.020 408.380 403.020 408.390 ;
        RECT 580.020 408.380 583.020 408.390 ;
        RECT 760.020 408.380 763.020 408.390 ;
        RECT 940.020 408.380 943.020 408.390 ;
        RECT 1120.020 408.380 1123.020 408.390 ;
        RECT 1300.020 408.380 1303.020 408.390 ;
        RECT 1480.020 408.380 1483.020 408.390 ;
        RECT 1660.020 408.380 1663.020 408.390 ;
        RECT 1840.020 408.380 1843.020 408.390 ;
        RECT 2020.020 408.380 2023.020 408.390 ;
        RECT 2200.020 408.380 2203.020 408.390 ;
        RECT 2380.020 408.380 2383.020 408.390 ;
        RECT 2560.020 408.380 2563.020 408.390 ;
        RECT 2740.020 408.380 2743.020 408.390 ;
        RECT 2945.000 408.380 2948.000 408.390 ;
        RECT -32.980 405.380 2952.600 408.380 ;
        RECT -28.380 405.370 -25.380 405.380 ;
        RECT 40.020 405.370 43.020 405.380 ;
        RECT 220.020 405.370 223.020 405.380 ;
        RECT 400.020 405.370 403.020 405.380 ;
        RECT 580.020 405.370 583.020 405.380 ;
        RECT 760.020 405.370 763.020 405.380 ;
        RECT 940.020 405.370 943.020 405.380 ;
        RECT 1120.020 405.370 1123.020 405.380 ;
        RECT 1300.020 405.370 1303.020 405.380 ;
        RECT 1480.020 405.370 1483.020 405.380 ;
        RECT 1660.020 405.370 1663.020 405.380 ;
        RECT 1840.020 405.370 1843.020 405.380 ;
        RECT 2020.020 405.370 2023.020 405.380 ;
        RECT 2200.020 405.370 2203.020 405.380 ;
        RECT 2380.020 405.370 2383.020 405.380 ;
        RECT 2560.020 405.370 2563.020 405.380 ;
        RECT 2740.020 405.370 2743.020 405.380 ;
        RECT 2945.000 405.370 2948.000 405.380 ;
        RECT -28.380 228.380 -25.380 228.390 ;
        RECT 40.020 228.380 43.020 228.390 ;
        RECT 220.020 228.380 223.020 228.390 ;
        RECT 400.020 228.380 403.020 228.390 ;
        RECT 580.020 228.380 583.020 228.390 ;
        RECT 760.020 228.380 763.020 228.390 ;
        RECT 940.020 228.380 943.020 228.390 ;
        RECT 1120.020 228.380 1123.020 228.390 ;
        RECT 1300.020 228.380 1303.020 228.390 ;
        RECT 1480.020 228.380 1483.020 228.390 ;
        RECT 1660.020 228.380 1663.020 228.390 ;
        RECT 1840.020 228.380 1843.020 228.390 ;
        RECT 2020.020 228.380 2023.020 228.390 ;
        RECT 2200.020 228.380 2203.020 228.390 ;
        RECT 2380.020 228.380 2383.020 228.390 ;
        RECT 2560.020 228.380 2563.020 228.390 ;
        RECT 2740.020 228.380 2743.020 228.390 ;
        RECT 2945.000 228.380 2948.000 228.390 ;
        RECT -32.980 225.380 2952.600 228.380 ;
        RECT -28.380 225.370 -25.380 225.380 ;
        RECT 40.020 225.370 43.020 225.380 ;
        RECT 220.020 225.370 223.020 225.380 ;
        RECT 400.020 225.370 403.020 225.380 ;
        RECT 580.020 225.370 583.020 225.380 ;
        RECT 760.020 225.370 763.020 225.380 ;
        RECT 940.020 225.370 943.020 225.380 ;
        RECT 1120.020 225.370 1123.020 225.380 ;
        RECT 1300.020 225.370 1303.020 225.380 ;
        RECT 1480.020 225.370 1483.020 225.380 ;
        RECT 1660.020 225.370 1663.020 225.380 ;
        RECT 1840.020 225.370 1843.020 225.380 ;
        RECT 2020.020 225.370 2023.020 225.380 ;
        RECT 2200.020 225.370 2203.020 225.380 ;
        RECT 2380.020 225.370 2383.020 225.380 ;
        RECT 2560.020 225.370 2563.020 225.380 ;
        RECT 2740.020 225.370 2743.020 225.380 ;
        RECT 2945.000 225.370 2948.000 225.380 ;
        RECT -28.380 48.380 -25.380 48.390 ;
        RECT 40.020 48.380 43.020 48.390 ;
        RECT 220.020 48.380 223.020 48.390 ;
        RECT 400.020 48.380 403.020 48.390 ;
        RECT 580.020 48.380 583.020 48.390 ;
        RECT 760.020 48.380 763.020 48.390 ;
        RECT 940.020 48.380 943.020 48.390 ;
        RECT 1120.020 48.380 1123.020 48.390 ;
        RECT 1300.020 48.380 1303.020 48.390 ;
        RECT 1480.020 48.380 1483.020 48.390 ;
        RECT 1660.020 48.380 1663.020 48.390 ;
        RECT 1840.020 48.380 1843.020 48.390 ;
        RECT 2020.020 48.380 2023.020 48.390 ;
        RECT 2200.020 48.380 2203.020 48.390 ;
        RECT 2380.020 48.380 2383.020 48.390 ;
        RECT 2560.020 48.380 2563.020 48.390 ;
        RECT 2740.020 48.380 2743.020 48.390 ;
        RECT 2945.000 48.380 2948.000 48.390 ;
        RECT -32.980 45.380 2952.600 48.380 ;
        RECT -28.380 45.370 -25.380 45.380 ;
        RECT 40.020 45.370 43.020 45.380 ;
        RECT 220.020 45.370 223.020 45.380 ;
        RECT 400.020 45.370 403.020 45.380 ;
        RECT 580.020 45.370 583.020 45.380 ;
        RECT 760.020 45.370 763.020 45.380 ;
        RECT 940.020 45.370 943.020 45.380 ;
        RECT 1120.020 45.370 1123.020 45.380 ;
        RECT 1300.020 45.370 1303.020 45.380 ;
        RECT 1480.020 45.370 1483.020 45.380 ;
        RECT 1660.020 45.370 1663.020 45.380 ;
        RECT 1840.020 45.370 1843.020 45.380 ;
        RECT 2020.020 45.370 2023.020 45.380 ;
        RECT 2200.020 45.370 2203.020 45.380 ;
        RECT 2380.020 45.370 2383.020 45.380 ;
        RECT 2560.020 45.370 2563.020 45.380 ;
        RECT 2740.020 45.370 2743.020 45.380 ;
        RECT 2945.000 45.370 2948.000 45.380 ;
        RECT -28.380 -20.020 -25.380 -20.010 ;
        RECT 40.020 -20.020 43.020 -20.010 ;
        RECT 220.020 -20.020 223.020 -20.010 ;
        RECT 400.020 -20.020 403.020 -20.010 ;
        RECT 580.020 -20.020 583.020 -20.010 ;
        RECT 760.020 -20.020 763.020 -20.010 ;
        RECT 940.020 -20.020 943.020 -20.010 ;
        RECT 1120.020 -20.020 1123.020 -20.010 ;
        RECT 1300.020 -20.020 1303.020 -20.010 ;
        RECT 1480.020 -20.020 1483.020 -20.010 ;
        RECT 1660.020 -20.020 1663.020 -20.010 ;
        RECT 1840.020 -20.020 1843.020 -20.010 ;
        RECT 2020.020 -20.020 2023.020 -20.010 ;
        RECT 2200.020 -20.020 2203.020 -20.010 ;
        RECT 2380.020 -20.020 2383.020 -20.010 ;
        RECT 2560.020 -20.020 2563.020 -20.010 ;
        RECT 2740.020 -20.020 2743.020 -20.010 ;
        RECT 2945.000 -20.020 2948.000 -20.010 ;
        RECT -28.380 -23.020 2948.000 -20.020 ;
        RECT -28.380 -23.030 -25.380 -23.020 ;
        RECT 40.020 -23.030 43.020 -23.020 ;
        RECT 220.020 -23.030 223.020 -23.020 ;
        RECT 400.020 -23.030 403.020 -23.020 ;
        RECT 580.020 -23.030 583.020 -23.020 ;
        RECT 760.020 -23.030 763.020 -23.020 ;
        RECT 940.020 -23.030 943.020 -23.020 ;
        RECT 1120.020 -23.030 1123.020 -23.020 ;
        RECT 1300.020 -23.030 1303.020 -23.020 ;
        RECT 1480.020 -23.030 1483.020 -23.020 ;
        RECT 1660.020 -23.030 1663.020 -23.020 ;
        RECT 1840.020 -23.030 1843.020 -23.020 ;
        RECT 2020.020 -23.030 2023.020 -23.020 ;
        RECT 2200.020 -23.030 2203.020 -23.020 ;
        RECT 2380.020 -23.030 2383.020 -23.020 ;
        RECT 2560.020 -23.030 2563.020 -23.020 ;
        RECT 2740.020 -23.030 2743.020 -23.020 ;
        RECT 2945.000 -23.030 2948.000 -23.020 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -32.980 -27.620 -29.980 3547.300 ;
        RECT 130.020 -27.620 133.020 3547.300 ;
        RECT 310.020 -27.620 313.020 3547.300 ;
        RECT 490.020 -27.620 493.020 3547.300 ;
        RECT 670.020 -27.620 673.020 3547.300 ;
        RECT 850.020 -27.620 853.020 3547.300 ;
        RECT 1030.020 -27.620 1033.020 3547.300 ;
        RECT 1210.020 -27.620 1213.020 3547.300 ;
        RECT 1390.020 -27.620 1393.020 3547.300 ;
        RECT 1570.020 -27.620 1573.020 3547.300 ;
        RECT 1750.020 -27.620 1753.020 3547.300 ;
        RECT 1930.020 -27.620 1933.020 3547.300 ;
        RECT 2110.020 -27.620 2113.020 3547.300 ;
        RECT 2290.020 -27.620 2293.020 3547.300 ;
        RECT 2470.020 -27.620 2473.020 3547.300 ;
        RECT 2650.020 -27.620 2653.020 3547.300 ;
        RECT 2830.020 -27.620 2833.020 3547.300 ;
        RECT 2949.600 -27.620 2952.600 3547.300 ;
      LAYER via4 ;
        RECT -32.070 3546.010 -30.890 3547.190 ;
        RECT -32.070 3544.410 -30.890 3545.590 ;
        RECT -32.070 3377.090 -30.890 3378.270 ;
        RECT -32.070 3375.490 -30.890 3376.670 ;
        RECT -32.070 3197.090 -30.890 3198.270 ;
        RECT -32.070 3195.490 -30.890 3196.670 ;
        RECT -32.070 3017.090 -30.890 3018.270 ;
        RECT -32.070 3015.490 -30.890 3016.670 ;
        RECT -32.070 2837.090 -30.890 2838.270 ;
        RECT -32.070 2835.490 -30.890 2836.670 ;
        RECT -32.070 2657.090 -30.890 2658.270 ;
        RECT -32.070 2655.490 -30.890 2656.670 ;
        RECT -32.070 2477.090 -30.890 2478.270 ;
        RECT -32.070 2475.490 -30.890 2476.670 ;
        RECT -32.070 2297.090 -30.890 2298.270 ;
        RECT -32.070 2295.490 -30.890 2296.670 ;
        RECT -32.070 2117.090 -30.890 2118.270 ;
        RECT -32.070 2115.490 -30.890 2116.670 ;
        RECT -32.070 1937.090 -30.890 1938.270 ;
        RECT -32.070 1935.490 -30.890 1936.670 ;
        RECT -32.070 1757.090 -30.890 1758.270 ;
        RECT -32.070 1755.490 -30.890 1756.670 ;
        RECT -32.070 1577.090 -30.890 1578.270 ;
        RECT -32.070 1575.490 -30.890 1576.670 ;
        RECT -32.070 1397.090 -30.890 1398.270 ;
        RECT -32.070 1395.490 -30.890 1396.670 ;
        RECT -32.070 1217.090 -30.890 1218.270 ;
        RECT -32.070 1215.490 -30.890 1216.670 ;
        RECT -32.070 1037.090 -30.890 1038.270 ;
        RECT -32.070 1035.490 -30.890 1036.670 ;
        RECT -32.070 857.090 -30.890 858.270 ;
        RECT -32.070 855.490 -30.890 856.670 ;
        RECT -32.070 677.090 -30.890 678.270 ;
        RECT -32.070 675.490 -30.890 676.670 ;
        RECT -32.070 497.090 -30.890 498.270 ;
        RECT -32.070 495.490 -30.890 496.670 ;
        RECT -32.070 317.090 -30.890 318.270 ;
        RECT -32.070 315.490 -30.890 316.670 ;
        RECT -32.070 137.090 -30.890 138.270 ;
        RECT -32.070 135.490 -30.890 136.670 ;
        RECT -32.070 -25.910 -30.890 -24.730 ;
        RECT -32.070 -27.510 -30.890 -26.330 ;
        RECT 130.930 3546.010 132.110 3547.190 ;
        RECT 130.930 3544.410 132.110 3545.590 ;
        RECT 130.930 3377.090 132.110 3378.270 ;
        RECT 130.930 3375.490 132.110 3376.670 ;
        RECT 130.930 3197.090 132.110 3198.270 ;
        RECT 130.930 3195.490 132.110 3196.670 ;
        RECT 130.930 3017.090 132.110 3018.270 ;
        RECT 130.930 3015.490 132.110 3016.670 ;
        RECT 130.930 2837.090 132.110 2838.270 ;
        RECT 130.930 2835.490 132.110 2836.670 ;
        RECT 130.930 2657.090 132.110 2658.270 ;
        RECT 130.930 2655.490 132.110 2656.670 ;
        RECT 130.930 2477.090 132.110 2478.270 ;
        RECT 130.930 2475.490 132.110 2476.670 ;
        RECT 130.930 2297.090 132.110 2298.270 ;
        RECT 130.930 2295.490 132.110 2296.670 ;
        RECT 130.930 2117.090 132.110 2118.270 ;
        RECT 130.930 2115.490 132.110 2116.670 ;
        RECT 130.930 1937.090 132.110 1938.270 ;
        RECT 130.930 1935.490 132.110 1936.670 ;
        RECT 130.930 1757.090 132.110 1758.270 ;
        RECT 130.930 1755.490 132.110 1756.670 ;
        RECT 130.930 1577.090 132.110 1578.270 ;
        RECT 130.930 1575.490 132.110 1576.670 ;
        RECT 130.930 1397.090 132.110 1398.270 ;
        RECT 130.930 1395.490 132.110 1396.670 ;
        RECT 130.930 1217.090 132.110 1218.270 ;
        RECT 130.930 1215.490 132.110 1216.670 ;
        RECT 130.930 1037.090 132.110 1038.270 ;
        RECT 130.930 1035.490 132.110 1036.670 ;
        RECT 130.930 857.090 132.110 858.270 ;
        RECT 130.930 855.490 132.110 856.670 ;
        RECT 130.930 677.090 132.110 678.270 ;
        RECT 130.930 675.490 132.110 676.670 ;
        RECT 130.930 497.090 132.110 498.270 ;
        RECT 130.930 495.490 132.110 496.670 ;
        RECT 130.930 317.090 132.110 318.270 ;
        RECT 130.930 315.490 132.110 316.670 ;
        RECT 130.930 137.090 132.110 138.270 ;
        RECT 130.930 135.490 132.110 136.670 ;
        RECT 130.930 -25.910 132.110 -24.730 ;
        RECT 130.930 -27.510 132.110 -26.330 ;
        RECT 310.930 3546.010 312.110 3547.190 ;
        RECT 310.930 3544.410 312.110 3545.590 ;
        RECT 310.930 3377.090 312.110 3378.270 ;
        RECT 310.930 3375.490 312.110 3376.670 ;
        RECT 310.930 3197.090 312.110 3198.270 ;
        RECT 310.930 3195.490 312.110 3196.670 ;
        RECT 310.930 3017.090 312.110 3018.270 ;
        RECT 310.930 3015.490 312.110 3016.670 ;
        RECT 310.930 2837.090 312.110 2838.270 ;
        RECT 310.930 2835.490 312.110 2836.670 ;
        RECT 310.930 2657.090 312.110 2658.270 ;
        RECT 310.930 2655.490 312.110 2656.670 ;
        RECT 310.930 2477.090 312.110 2478.270 ;
        RECT 310.930 2475.490 312.110 2476.670 ;
        RECT 310.930 2297.090 312.110 2298.270 ;
        RECT 310.930 2295.490 312.110 2296.670 ;
        RECT 310.930 2117.090 312.110 2118.270 ;
        RECT 310.930 2115.490 312.110 2116.670 ;
        RECT 310.930 1937.090 312.110 1938.270 ;
        RECT 310.930 1935.490 312.110 1936.670 ;
        RECT 310.930 1757.090 312.110 1758.270 ;
        RECT 310.930 1755.490 312.110 1756.670 ;
        RECT 310.930 1577.090 312.110 1578.270 ;
        RECT 310.930 1575.490 312.110 1576.670 ;
        RECT 310.930 1397.090 312.110 1398.270 ;
        RECT 310.930 1395.490 312.110 1396.670 ;
        RECT 310.930 1217.090 312.110 1218.270 ;
        RECT 310.930 1215.490 312.110 1216.670 ;
        RECT 310.930 1037.090 312.110 1038.270 ;
        RECT 310.930 1035.490 312.110 1036.670 ;
        RECT 310.930 857.090 312.110 858.270 ;
        RECT 310.930 855.490 312.110 856.670 ;
        RECT 310.930 677.090 312.110 678.270 ;
        RECT 310.930 675.490 312.110 676.670 ;
        RECT 310.930 497.090 312.110 498.270 ;
        RECT 310.930 495.490 312.110 496.670 ;
        RECT 310.930 317.090 312.110 318.270 ;
        RECT 310.930 315.490 312.110 316.670 ;
        RECT 310.930 137.090 312.110 138.270 ;
        RECT 310.930 135.490 312.110 136.670 ;
        RECT 310.930 -25.910 312.110 -24.730 ;
        RECT 310.930 -27.510 312.110 -26.330 ;
        RECT 490.930 3546.010 492.110 3547.190 ;
        RECT 490.930 3544.410 492.110 3545.590 ;
        RECT 490.930 3377.090 492.110 3378.270 ;
        RECT 490.930 3375.490 492.110 3376.670 ;
        RECT 490.930 3197.090 492.110 3198.270 ;
        RECT 490.930 3195.490 492.110 3196.670 ;
        RECT 490.930 3017.090 492.110 3018.270 ;
        RECT 490.930 3015.490 492.110 3016.670 ;
        RECT 490.930 2837.090 492.110 2838.270 ;
        RECT 490.930 2835.490 492.110 2836.670 ;
        RECT 490.930 2657.090 492.110 2658.270 ;
        RECT 490.930 2655.490 492.110 2656.670 ;
        RECT 490.930 2477.090 492.110 2478.270 ;
        RECT 490.930 2475.490 492.110 2476.670 ;
        RECT 490.930 2297.090 492.110 2298.270 ;
        RECT 490.930 2295.490 492.110 2296.670 ;
        RECT 490.930 2117.090 492.110 2118.270 ;
        RECT 490.930 2115.490 492.110 2116.670 ;
        RECT 490.930 1937.090 492.110 1938.270 ;
        RECT 490.930 1935.490 492.110 1936.670 ;
        RECT 490.930 1757.090 492.110 1758.270 ;
        RECT 490.930 1755.490 492.110 1756.670 ;
        RECT 490.930 1577.090 492.110 1578.270 ;
        RECT 490.930 1575.490 492.110 1576.670 ;
        RECT 490.930 1397.090 492.110 1398.270 ;
        RECT 490.930 1395.490 492.110 1396.670 ;
        RECT 490.930 1217.090 492.110 1218.270 ;
        RECT 490.930 1215.490 492.110 1216.670 ;
        RECT 490.930 1037.090 492.110 1038.270 ;
        RECT 490.930 1035.490 492.110 1036.670 ;
        RECT 490.930 857.090 492.110 858.270 ;
        RECT 490.930 855.490 492.110 856.670 ;
        RECT 490.930 677.090 492.110 678.270 ;
        RECT 490.930 675.490 492.110 676.670 ;
        RECT 490.930 497.090 492.110 498.270 ;
        RECT 490.930 495.490 492.110 496.670 ;
        RECT 490.930 317.090 492.110 318.270 ;
        RECT 490.930 315.490 492.110 316.670 ;
        RECT 490.930 137.090 492.110 138.270 ;
        RECT 490.930 135.490 492.110 136.670 ;
        RECT 490.930 -25.910 492.110 -24.730 ;
        RECT 490.930 -27.510 492.110 -26.330 ;
        RECT 670.930 3546.010 672.110 3547.190 ;
        RECT 670.930 3544.410 672.110 3545.590 ;
        RECT 670.930 3377.090 672.110 3378.270 ;
        RECT 670.930 3375.490 672.110 3376.670 ;
        RECT 670.930 3197.090 672.110 3198.270 ;
        RECT 670.930 3195.490 672.110 3196.670 ;
        RECT 670.930 3017.090 672.110 3018.270 ;
        RECT 670.930 3015.490 672.110 3016.670 ;
        RECT 670.930 2837.090 672.110 2838.270 ;
        RECT 670.930 2835.490 672.110 2836.670 ;
        RECT 670.930 2657.090 672.110 2658.270 ;
        RECT 670.930 2655.490 672.110 2656.670 ;
        RECT 670.930 2477.090 672.110 2478.270 ;
        RECT 670.930 2475.490 672.110 2476.670 ;
        RECT 670.930 2297.090 672.110 2298.270 ;
        RECT 670.930 2295.490 672.110 2296.670 ;
        RECT 670.930 2117.090 672.110 2118.270 ;
        RECT 670.930 2115.490 672.110 2116.670 ;
        RECT 670.930 1937.090 672.110 1938.270 ;
        RECT 670.930 1935.490 672.110 1936.670 ;
        RECT 670.930 1757.090 672.110 1758.270 ;
        RECT 670.930 1755.490 672.110 1756.670 ;
        RECT 670.930 1577.090 672.110 1578.270 ;
        RECT 670.930 1575.490 672.110 1576.670 ;
        RECT 670.930 1397.090 672.110 1398.270 ;
        RECT 670.930 1395.490 672.110 1396.670 ;
        RECT 670.930 1217.090 672.110 1218.270 ;
        RECT 670.930 1215.490 672.110 1216.670 ;
        RECT 670.930 1037.090 672.110 1038.270 ;
        RECT 670.930 1035.490 672.110 1036.670 ;
        RECT 670.930 857.090 672.110 858.270 ;
        RECT 670.930 855.490 672.110 856.670 ;
        RECT 670.930 677.090 672.110 678.270 ;
        RECT 670.930 675.490 672.110 676.670 ;
        RECT 670.930 497.090 672.110 498.270 ;
        RECT 670.930 495.490 672.110 496.670 ;
        RECT 670.930 317.090 672.110 318.270 ;
        RECT 670.930 315.490 672.110 316.670 ;
        RECT 670.930 137.090 672.110 138.270 ;
        RECT 670.930 135.490 672.110 136.670 ;
        RECT 670.930 -25.910 672.110 -24.730 ;
        RECT 670.930 -27.510 672.110 -26.330 ;
        RECT 850.930 3546.010 852.110 3547.190 ;
        RECT 850.930 3544.410 852.110 3545.590 ;
        RECT 850.930 3377.090 852.110 3378.270 ;
        RECT 850.930 3375.490 852.110 3376.670 ;
        RECT 850.930 3197.090 852.110 3198.270 ;
        RECT 850.930 3195.490 852.110 3196.670 ;
        RECT 850.930 3017.090 852.110 3018.270 ;
        RECT 850.930 3015.490 852.110 3016.670 ;
        RECT 850.930 2837.090 852.110 2838.270 ;
        RECT 850.930 2835.490 852.110 2836.670 ;
        RECT 850.930 2657.090 852.110 2658.270 ;
        RECT 850.930 2655.490 852.110 2656.670 ;
        RECT 850.930 2477.090 852.110 2478.270 ;
        RECT 850.930 2475.490 852.110 2476.670 ;
        RECT 850.930 2297.090 852.110 2298.270 ;
        RECT 850.930 2295.490 852.110 2296.670 ;
        RECT 850.930 2117.090 852.110 2118.270 ;
        RECT 850.930 2115.490 852.110 2116.670 ;
        RECT 850.930 1937.090 852.110 1938.270 ;
        RECT 850.930 1935.490 852.110 1936.670 ;
        RECT 850.930 1757.090 852.110 1758.270 ;
        RECT 850.930 1755.490 852.110 1756.670 ;
        RECT 850.930 1577.090 852.110 1578.270 ;
        RECT 850.930 1575.490 852.110 1576.670 ;
        RECT 850.930 1397.090 852.110 1398.270 ;
        RECT 850.930 1395.490 852.110 1396.670 ;
        RECT 850.930 1217.090 852.110 1218.270 ;
        RECT 850.930 1215.490 852.110 1216.670 ;
        RECT 850.930 1037.090 852.110 1038.270 ;
        RECT 850.930 1035.490 852.110 1036.670 ;
        RECT 850.930 857.090 852.110 858.270 ;
        RECT 850.930 855.490 852.110 856.670 ;
        RECT 850.930 677.090 852.110 678.270 ;
        RECT 850.930 675.490 852.110 676.670 ;
        RECT 850.930 497.090 852.110 498.270 ;
        RECT 850.930 495.490 852.110 496.670 ;
        RECT 850.930 317.090 852.110 318.270 ;
        RECT 850.930 315.490 852.110 316.670 ;
        RECT 850.930 137.090 852.110 138.270 ;
        RECT 850.930 135.490 852.110 136.670 ;
        RECT 850.930 -25.910 852.110 -24.730 ;
        RECT 850.930 -27.510 852.110 -26.330 ;
        RECT 1030.930 3546.010 1032.110 3547.190 ;
        RECT 1030.930 3544.410 1032.110 3545.590 ;
        RECT 1030.930 3377.090 1032.110 3378.270 ;
        RECT 1030.930 3375.490 1032.110 3376.670 ;
        RECT 1030.930 3197.090 1032.110 3198.270 ;
        RECT 1030.930 3195.490 1032.110 3196.670 ;
        RECT 1030.930 3017.090 1032.110 3018.270 ;
        RECT 1030.930 3015.490 1032.110 3016.670 ;
        RECT 1030.930 2837.090 1032.110 2838.270 ;
        RECT 1030.930 2835.490 1032.110 2836.670 ;
        RECT 1030.930 2657.090 1032.110 2658.270 ;
        RECT 1030.930 2655.490 1032.110 2656.670 ;
        RECT 1030.930 2477.090 1032.110 2478.270 ;
        RECT 1030.930 2475.490 1032.110 2476.670 ;
        RECT 1030.930 2297.090 1032.110 2298.270 ;
        RECT 1030.930 2295.490 1032.110 2296.670 ;
        RECT 1030.930 2117.090 1032.110 2118.270 ;
        RECT 1030.930 2115.490 1032.110 2116.670 ;
        RECT 1030.930 1937.090 1032.110 1938.270 ;
        RECT 1030.930 1935.490 1032.110 1936.670 ;
        RECT 1030.930 1757.090 1032.110 1758.270 ;
        RECT 1030.930 1755.490 1032.110 1756.670 ;
        RECT 1030.930 1577.090 1032.110 1578.270 ;
        RECT 1030.930 1575.490 1032.110 1576.670 ;
        RECT 1030.930 1397.090 1032.110 1398.270 ;
        RECT 1030.930 1395.490 1032.110 1396.670 ;
        RECT 1030.930 1217.090 1032.110 1218.270 ;
        RECT 1030.930 1215.490 1032.110 1216.670 ;
        RECT 1030.930 1037.090 1032.110 1038.270 ;
        RECT 1030.930 1035.490 1032.110 1036.670 ;
        RECT 1030.930 857.090 1032.110 858.270 ;
        RECT 1030.930 855.490 1032.110 856.670 ;
        RECT 1030.930 677.090 1032.110 678.270 ;
        RECT 1030.930 675.490 1032.110 676.670 ;
        RECT 1030.930 497.090 1032.110 498.270 ;
        RECT 1030.930 495.490 1032.110 496.670 ;
        RECT 1030.930 317.090 1032.110 318.270 ;
        RECT 1030.930 315.490 1032.110 316.670 ;
        RECT 1030.930 137.090 1032.110 138.270 ;
        RECT 1030.930 135.490 1032.110 136.670 ;
        RECT 1030.930 -25.910 1032.110 -24.730 ;
        RECT 1030.930 -27.510 1032.110 -26.330 ;
        RECT 1210.930 3546.010 1212.110 3547.190 ;
        RECT 1210.930 3544.410 1212.110 3545.590 ;
        RECT 1210.930 3377.090 1212.110 3378.270 ;
        RECT 1210.930 3375.490 1212.110 3376.670 ;
        RECT 1210.930 3197.090 1212.110 3198.270 ;
        RECT 1210.930 3195.490 1212.110 3196.670 ;
        RECT 1210.930 3017.090 1212.110 3018.270 ;
        RECT 1210.930 3015.490 1212.110 3016.670 ;
        RECT 1210.930 2837.090 1212.110 2838.270 ;
        RECT 1210.930 2835.490 1212.110 2836.670 ;
        RECT 1210.930 2657.090 1212.110 2658.270 ;
        RECT 1210.930 2655.490 1212.110 2656.670 ;
        RECT 1210.930 2477.090 1212.110 2478.270 ;
        RECT 1210.930 2475.490 1212.110 2476.670 ;
        RECT 1210.930 2297.090 1212.110 2298.270 ;
        RECT 1210.930 2295.490 1212.110 2296.670 ;
        RECT 1210.930 2117.090 1212.110 2118.270 ;
        RECT 1210.930 2115.490 1212.110 2116.670 ;
        RECT 1210.930 1937.090 1212.110 1938.270 ;
        RECT 1210.930 1935.490 1212.110 1936.670 ;
        RECT 1210.930 1757.090 1212.110 1758.270 ;
        RECT 1210.930 1755.490 1212.110 1756.670 ;
        RECT 1210.930 1577.090 1212.110 1578.270 ;
        RECT 1210.930 1575.490 1212.110 1576.670 ;
        RECT 1210.930 1397.090 1212.110 1398.270 ;
        RECT 1210.930 1395.490 1212.110 1396.670 ;
        RECT 1210.930 1217.090 1212.110 1218.270 ;
        RECT 1210.930 1215.490 1212.110 1216.670 ;
        RECT 1210.930 1037.090 1212.110 1038.270 ;
        RECT 1210.930 1035.490 1212.110 1036.670 ;
        RECT 1210.930 857.090 1212.110 858.270 ;
        RECT 1210.930 855.490 1212.110 856.670 ;
        RECT 1210.930 677.090 1212.110 678.270 ;
        RECT 1210.930 675.490 1212.110 676.670 ;
        RECT 1210.930 497.090 1212.110 498.270 ;
        RECT 1210.930 495.490 1212.110 496.670 ;
        RECT 1210.930 317.090 1212.110 318.270 ;
        RECT 1210.930 315.490 1212.110 316.670 ;
        RECT 1210.930 137.090 1212.110 138.270 ;
        RECT 1210.930 135.490 1212.110 136.670 ;
        RECT 1210.930 -25.910 1212.110 -24.730 ;
        RECT 1210.930 -27.510 1212.110 -26.330 ;
        RECT 1390.930 3546.010 1392.110 3547.190 ;
        RECT 1390.930 3544.410 1392.110 3545.590 ;
        RECT 1390.930 3377.090 1392.110 3378.270 ;
        RECT 1390.930 3375.490 1392.110 3376.670 ;
        RECT 1390.930 3197.090 1392.110 3198.270 ;
        RECT 1390.930 3195.490 1392.110 3196.670 ;
        RECT 1390.930 3017.090 1392.110 3018.270 ;
        RECT 1390.930 3015.490 1392.110 3016.670 ;
        RECT 1390.930 2837.090 1392.110 2838.270 ;
        RECT 1390.930 2835.490 1392.110 2836.670 ;
        RECT 1390.930 2657.090 1392.110 2658.270 ;
        RECT 1390.930 2655.490 1392.110 2656.670 ;
        RECT 1390.930 2477.090 1392.110 2478.270 ;
        RECT 1390.930 2475.490 1392.110 2476.670 ;
        RECT 1390.930 2297.090 1392.110 2298.270 ;
        RECT 1390.930 2295.490 1392.110 2296.670 ;
        RECT 1390.930 2117.090 1392.110 2118.270 ;
        RECT 1390.930 2115.490 1392.110 2116.670 ;
        RECT 1390.930 1937.090 1392.110 1938.270 ;
        RECT 1390.930 1935.490 1392.110 1936.670 ;
        RECT 1390.930 1757.090 1392.110 1758.270 ;
        RECT 1390.930 1755.490 1392.110 1756.670 ;
        RECT 1390.930 1577.090 1392.110 1578.270 ;
        RECT 1390.930 1575.490 1392.110 1576.670 ;
        RECT 1390.930 1397.090 1392.110 1398.270 ;
        RECT 1390.930 1395.490 1392.110 1396.670 ;
        RECT 1390.930 1217.090 1392.110 1218.270 ;
        RECT 1390.930 1215.490 1392.110 1216.670 ;
        RECT 1390.930 1037.090 1392.110 1038.270 ;
        RECT 1390.930 1035.490 1392.110 1036.670 ;
        RECT 1390.930 857.090 1392.110 858.270 ;
        RECT 1390.930 855.490 1392.110 856.670 ;
        RECT 1390.930 677.090 1392.110 678.270 ;
        RECT 1390.930 675.490 1392.110 676.670 ;
        RECT 1390.930 497.090 1392.110 498.270 ;
        RECT 1390.930 495.490 1392.110 496.670 ;
        RECT 1390.930 317.090 1392.110 318.270 ;
        RECT 1390.930 315.490 1392.110 316.670 ;
        RECT 1390.930 137.090 1392.110 138.270 ;
        RECT 1390.930 135.490 1392.110 136.670 ;
        RECT 1390.930 -25.910 1392.110 -24.730 ;
        RECT 1390.930 -27.510 1392.110 -26.330 ;
        RECT 1570.930 3546.010 1572.110 3547.190 ;
        RECT 1570.930 3544.410 1572.110 3545.590 ;
        RECT 1570.930 3377.090 1572.110 3378.270 ;
        RECT 1570.930 3375.490 1572.110 3376.670 ;
        RECT 1570.930 3197.090 1572.110 3198.270 ;
        RECT 1570.930 3195.490 1572.110 3196.670 ;
        RECT 1570.930 3017.090 1572.110 3018.270 ;
        RECT 1570.930 3015.490 1572.110 3016.670 ;
        RECT 1570.930 2837.090 1572.110 2838.270 ;
        RECT 1570.930 2835.490 1572.110 2836.670 ;
        RECT 1570.930 2657.090 1572.110 2658.270 ;
        RECT 1570.930 2655.490 1572.110 2656.670 ;
        RECT 1570.930 2477.090 1572.110 2478.270 ;
        RECT 1570.930 2475.490 1572.110 2476.670 ;
        RECT 1570.930 2297.090 1572.110 2298.270 ;
        RECT 1570.930 2295.490 1572.110 2296.670 ;
        RECT 1570.930 2117.090 1572.110 2118.270 ;
        RECT 1570.930 2115.490 1572.110 2116.670 ;
        RECT 1570.930 1937.090 1572.110 1938.270 ;
        RECT 1570.930 1935.490 1572.110 1936.670 ;
        RECT 1570.930 1757.090 1572.110 1758.270 ;
        RECT 1570.930 1755.490 1572.110 1756.670 ;
        RECT 1570.930 1577.090 1572.110 1578.270 ;
        RECT 1570.930 1575.490 1572.110 1576.670 ;
        RECT 1570.930 1397.090 1572.110 1398.270 ;
        RECT 1570.930 1395.490 1572.110 1396.670 ;
        RECT 1570.930 1217.090 1572.110 1218.270 ;
        RECT 1570.930 1215.490 1572.110 1216.670 ;
        RECT 1570.930 1037.090 1572.110 1038.270 ;
        RECT 1570.930 1035.490 1572.110 1036.670 ;
        RECT 1570.930 857.090 1572.110 858.270 ;
        RECT 1570.930 855.490 1572.110 856.670 ;
        RECT 1570.930 677.090 1572.110 678.270 ;
        RECT 1570.930 675.490 1572.110 676.670 ;
        RECT 1570.930 497.090 1572.110 498.270 ;
        RECT 1570.930 495.490 1572.110 496.670 ;
        RECT 1570.930 317.090 1572.110 318.270 ;
        RECT 1570.930 315.490 1572.110 316.670 ;
        RECT 1570.930 137.090 1572.110 138.270 ;
        RECT 1570.930 135.490 1572.110 136.670 ;
        RECT 1570.930 -25.910 1572.110 -24.730 ;
        RECT 1570.930 -27.510 1572.110 -26.330 ;
        RECT 1750.930 3546.010 1752.110 3547.190 ;
        RECT 1750.930 3544.410 1752.110 3545.590 ;
        RECT 1750.930 3377.090 1752.110 3378.270 ;
        RECT 1750.930 3375.490 1752.110 3376.670 ;
        RECT 1750.930 3197.090 1752.110 3198.270 ;
        RECT 1750.930 3195.490 1752.110 3196.670 ;
        RECT 1750.930 3017.090 1752.110 3018.270 ;
        RECT 1750.930 3015.490 1752.110 3016.670 ;
        RECT 1750.930 2837.090 1752.110 2838.270 ;
        RECT 1750.930 2835.490 1752.110 2836.670 ;
        RECT 1750.930 2657.090 1752.110 2658.270 ;
        RECT 1750.930 2655.490 1752.110 2656.670 ;
        RECT 1750.930 2477.090 1752.110 2478.270 ;
        RECT 1750.930 2475.490 1752.110 2476.670 ;
        RECT 1750.930 2297.090 1752.110 2298.270 ;
        RECT 1750.930 2295.490 1752.110 2296.670 ;
        RECT 1750.930 2117.090 1752.110 2118.270 ;
        RECT 1750.930 2115.490 1752.110 2116.670 ;
        RECT 1750.930 1937.090 1752.110 1938.270 ;
        RECT 1750.930 1935.490 1752.110 1936.670 ;
        RECT 1750.930 1757.090 1752.110 1758.270 ;
        RECT 1750.930 1755.490 1752.110 1756.670 ;
        RECT 1750.930 1577.090 1752.110 1578.270 ;
        RECT 1750.930 1575.490 1752.110 1576.670 ;
        RECT 1750.930 1397.090 1752.110 1398.270 ;
        RECT 1750.930 1395.490 1752.110 1396.670 ;
        RECT 1750.930 1217.090 1752.110 1218.270 ;
        RECT 1750.930 1215.490 1752.110 1216.670 ;
        RECT 1750.930 1037.090 1752.110 1038.270 ;
        RECT 1750.930 1035.490 1752.110 1036.670 ;
        RECT 1750.930 857.090 1752.110 858.270 ;
        RECT 1750.930 855.490 1752.110 856.670 ;
        RECT 1750.930 677.090 1752.110 678.270 ;
        RECT 1750.930 675.490 1752.110 676.670 ;
        RECT 1750.930 497.090 1752.110 498.270 ;
        RECT 1750.930 495.490 1752.110 496.670 ;
        RECT 1750.930 317.090 1752.110 318.270 ;
        RECT 1750.930 315.490 1752.110 316.670 ;
        RECT 1750.930 137.090 1752.110 138.270 ;
        RECT 1750.930 135.490 1752.110 136.670 ;
        RECT 1750.930 -25.910 1752.110 -24.730 ;
        RECT 1750.930 -27.510 1752.110 -26.330 ;
        RECT 1930.930 3546.010 1932.110 3547.190 ;
        RECT 1930.930 3544.410 1932.110 3545.590 ;
        RECT 1930.930 3377.090 1932.110 3378.270 ;
        RECT 1930.930 3375.490 1932.110 3376.670 ;
        RECT 1930.930 3197.090 1932.110 3198.270 ;
        RECT 1930.930 3195.490 1932.110 3196.670 ;
        RECT 1930.930 3017.090 1932.110 3018.270 ;
        RECT 1930.930 3015.490 1932.110 3016.670 ;
        RECT 1930.930 2837.090 1932.110 2838.270 ;
        RECT 1930.930 2835.490 1932.110 2836.670 ;
        RECT 1930.930 2657.090 1932.110 2658.270 ;
        RECT 1930.930 2655.490 1932.110 2656.670 ;
        RECT 1930.930 2477.090 1932.110 2478.270 ;
        RECT 1930.930 2475.490 1932.110 2476.670 ;
        RECT 1930.930 2297.090 1932.110 2298.270 ;
        RECT 1930.930 2295.490 1932.110 2296.670 ;
        RECT 1930.930 2117.090 1932.110 2118.270 ;
        RECT 1930.930 2115.490 1932.110 2116.670 ;
        RECT 1930.930 1937.090 1932.110 1938.270 ;
        RECT 1930.930 1935.490 1932.110 1936.670 ;
        RECT 1930.930 1757.090 1932.110 1758.270 ;
        RECT 1930.930 1755.490 1932.110 1756.670 ;
        RECT 1930.930 1577.090 1932.110 1578.270 ;
        RECT 1930.930 1575.490 1932.110 1576.670 ;
        RECT 1930.930 1397.090 1932.110 1398.270 ;
        RECT 1930.930 1395.490 1932.110 1396.670 ;
        RECT 1930.930 1217.090 1932.110 1218.270 ;
        RECT 1930.930 1215.490 1932.110 1216.670 ;
        RECT 1930.930 1037.090 1932.110 1038.270 ;
        RECT 1930.930 1035.490 1932.110 1036.670 ;
        RECT 1930.930 857.090 1932.110 858.270 ;
        RECT 1930.930 855.490 1932.110 856.670 ;
        RECT 1930.930 677.090 1932.110 678.270 ;
        RECT 1930.930 675.490 1932.110 676.670 ;
        RECT 1930.930 497.090 1932.110 498.270 ;
        RECT 1930.930 495.490 1932.110 496.670 ;
        RECT 1930.930 317.090 1932.110 318.270 ;
        RECT 1930.930 315.490 1932.110 316.670 ;
        RECT 1930.930 137.090 1932.110 138.270 ;
        RECT 1930.930 135.490 1932.110 136.670 ;
        RECT 1930.930 -25.910 1932.110 -24.730 ;
        RECT 1930.930 -27.510 1932.110 -26.330 ;
        RECT 2110.930 3546.010 2112.110 3547.190 ;
        RECT 2110.930 3544.410 2112.110 3545.590 ;
        RECT 2110.930 3377.090 2112.110 3378.270 ;
        RECT 2110.930 3375.490 2112.110 3376.670 ;
        RECT 2110.930 3197.090 2112.110 3198.270 ;
        RECT 2110.930 3195.490 2112.110 3196.670 ;
        RECT 2110.930 3017.090 2112.110 3018.270 ;
        RECT 2110.930 3015.490 2112.110 3016.670 ;
        RECT 2110.930 2837.090 2112.110 2838.270 ;
        RECT 2110.930 2835.490 2112.110 2836.670 ;
        RECT 2110.930 2657.090 2112.110 2658.270 ;
        RECT 2110.930 2655.490 2112.110 2656.670 ;
        RECT 2110.930 2477.090 2112.110 2478.270 ;
        RECT 2110.930 2475.490 2112.110 2476.670 ;
        RECT 2110.930 2297.090 2112.110 2298.270 ;
        RECT 2110.930 2295.490 2112.110 2296.670 ;
        RECT 2110.930 2117.090 2112.110 2118.270 ;
        RECT 2110.930 2115.490 2112.110 2116.670 ;
        RECT 2110.930 1937.090 2112.110 1938.270 ;
        RECT 2110.930 1935.490 2112.110 1936.670 ;
        RECT 2110.930 1757.090 2112.110 1758.270 ;
        RECT 2110.930 1755.490 2112.110 1756.670 ;
        RECT 2110.930 1577.090 2112.110 1578.270 ;
        RECT 2110.930 1575.490 2112.110 1576.670 ;
        RECT 2110.930 1397.090 2112.110 1398.270 ;
        RECT 2110.930 1395.490 2112.110 1396.670 ;
        RECT 2110.930 1217.090 2112.110 1218.270 ;
        RECT 2110.930 1215.490 2112.110 1216.670 ;
        RECT 2110.930 1037.090 2112.110 1038.270 ;
        RECT 2110.930 1035.490 2112.110 1036.670 ;
        RECT 2110.930 857.090 2112.110 858.270 ;
        RECT 2110.930 855.490 2112.110 856.670 ;
        RECT 2110.930 677.090 2112.110 678.270 ;
        RECT 2110.930 675.490 2112.110 676.670 ;
        RECT 2110.930 497.090 2112.110 498.270 ;
        RECT 2110.930 495.490 2112.110 496.670 ;
        RECT 2110.930 317.090 2112.110 318.270 ;
        RECT 2110.930 315.490 2112.110 316.670 ;
        RECT 2110.930 137.090 2112.110 138.270 ;
        RECT 2110.930 135.490 2112.110 136.670 ;
        RECT 2110.930 -25.910 2112.110 -24.730 ;
        RECT 2110.930 -27.510 2112.110 -26.330 ;
        RECT 2290.930 3546.010 2292.110 3547.190 ;
        RECT 2290.930 3544.410 2292.110 3545.590 ;
        RECT 2290.930 3377.090 2292.110 3378.270 ;
        RECT 2290.930 3375.490 2292.110 3376.670 ;
        RECT 2290.930 3197.090 2292.110 3198.270 ;
        RECT 2290.930 3195.490 2292.110 3196.670 ;
        RECT 2290.930 3017.090 2292.110 3018.270 ;
        RECT 2290.930 3015.490 2292.110 3016.670 ;
        RECT 2290.930 2837.090 2292.110 2838.270 ;
        RECT 2290.930 2835.490 2292.110 2836.670 ;
        RECT 2290.930 2657.090 2292.110 2658.270 ;
        RECT 2290.930 2655.490 2292.110 2656.670 ;
        RECT 2290.930 2477.090 2292.110 2478.270 ;
        RECT 2290.930 2475.490 2292.110 2476.670 ;
        RECT 2290.930 2297.090 2292.110 2298.270 ;
        RECT 2290.930 2295.490 2292.110 2296.670 ;
        RECT 2290.930 2117.090 2292.110 2118.270 ;
        RECT 2290.930 2115.490 2292.110 2116.670 ;
        RECT 2290.930 1937.090 2292.110 1938.270 ;
        RECT 2290.930 1935.490 2292.110 1936.670 ;
        RECT 2290.930 1757.090 2292.110 1758.270 ;
        RECT 2290.930 1755.490 2292.110 1756.670 ;
        RECT 2290.930 1577.090 2292.110 1578.270 ;
        RECT 2290.930 1575.490 2292.110 1576.670 ;
        RECT 2290.930 1397.090 2292.110 1398.270 ;
        RECT 2290.930 1395.490 2292.110 1396.670 ;
        RECT 2290.930 1217.090 2292.110 1218.270 ;
        RECT 2290.930 1215.490 2292.110 1216.670 ;
        RECT 2290.930 1037.090 2292.110 1038.270 ;
        RECT 2290.930 1035.490 2292.110 1036.670 ;
        RECT 2290.930 857.090 2292.110 858.270 ;
        RECT 2290.930 855.490 2292.110 856.670 ;
        RECT 2290.930 677.090 2292.110 678.270 ;
        RECT 2290.930 675.490 2292.110 676.670 ;
        RECT 2290.930 497.090 2292.110 498.270 ;
        RECT 2290.930 495.490 2292.110 496.670 ;
        RECT 2290.930 317.090 2292.110 318.270 ;
        RECT 2290.930 315.490 2292.110 316.670 ;
        RECT 2290.930 137.090 2292.110 138.270 ;
        RECT 2290.930 135.490 2292.110 136.670 ;
        RECT 2290.930 -25.910 2292.110 -24.730 ;
        RECT 2290.930 -27.510 2292.110 -26.330 ;
        RECT 2470.930 3546.010 2472.110 3547.190 ;
        RECT 2470.930 3544.410 2472.110 3545.590 ;
        RECT 2470.930 3377.090 2472.110 3378.270 ;
        RECT 2470.930 3375.490 2472.110 3376.670 ;
        RECT 2470.930 3197.090 2472.110 3198.270 ;
        RECT 2470.930 3195.490 2472.110 3196.670 ;
        RECT 2470.930 3017.090 2472.110 3018.270 ;
        RECT 2470.930 3015.490 2472.110 3016.670 ;
        RECT 2470.930 2837.090 2472.110 2838.270 ;
        RECT 2470.930 2835.490 2472.110 2836.670 ;
        RECT 2470.930 2657.090 2472.110 2658.270 ;
        RECT 2470.930 2655.490 2472.110 2656.670 ;
        RECT 2470.930 2477.090 2472.110 2478.270 ;
        RECT 2470.930 2475.490 2472.110 2476.670 ;
        RECT 2470.930 2297.090 2472.110 2298.270 ;
        RECT 2470.930 2295.490 2472.110 2296.670 ;
        RECT 2470.930 2117.090 2472.110 2118.270 ;
        RECT 2470.930 2115.490 2472.110 2116.670 ;
        RECT 2470.930 1937.090 2472.110 1938.270 ;
        RECT 2470.930 1935.490 2472.110 1936.670 ;
        RECT 2470.930 1757.090 2472.110 1758.270 ;
        RECT 2470.930 1755.490 2472.110 1756.670 ;
        RECT 2470.930 1577.090 2472.110 1578.270 ;
        RECT 2470.930 1575.490 2472.110 1576.670 ;
        RECT 2470.930 1397.090 2472.110 1398.270 ;
        RECT 2470.930 1395.490 2472.110 1396.670 ;
        RECT 2470.930 1217.090 2472.110 1218.270 ;
        RECT 2470.930 1215.490 2472.110 1216.670 ;
        RECT 2470.930 1037.090 2472.110 1038.270 ;
        RECT 2470.930 1035.490 2472.110 1036.670 ;
        RECT 2470.930 857.090 2472.110 858.270 ;
        RECT 2470.930 855.490 2472.110 856.670 ;
        RECT 2470.930 677.090 2472.110 678.270 ;
        RECT 2470.930 675.490 2472.110 676.670 ;
        RECT 2470.930 497.090 2472.110 498.270 ;
        RECT 2470.930 495.490 2472.110 496.670 ;
        RECT 2470.930 317.090 2472.110 318.270 ;
        RECT 2470.930 315.490 2472.110 316.670 ;
        RECT 2470.930 137.090 2472.110 138.270 ;
        RECT 2470.930 135.490 2472.110 136.670 ;
        RECT 2470.930 -25.910 2472.110 -24.730 ;
        RECT 2470.930 -27.510 2472.110 -26.330 ;
        RECT 2650.930 3546.010 2652.110 3547.190 ;
        RECT 2650.930 3544.410 2652.110 3545.590 ;
        RECT 2650.930 3377.090 2652.110 3378.270 ;
        RECT 2650.930 3375.490 2652.110 3376.670 ;
        RECT 2650.930 3197.090 2652.110 3198.270 ;
        RECT 2650.930 3195.490 2652.110 3196.670 ;
        RECT 2650.930 3017.090 2652.110 3018.270 ;
        RECT 2650.930 3015.490 2652.110 3016.670 ;
        RECT 2650.930 2837.090 2652.110 2838.270 ;
        RECT 2650.930 2835.490 2652.110 2836.670 ;
        RECT 2650.930 2657.090 2652.110 2658.270 ;
        RECT 2650.930 2655.490 2652.110 2656.670 ;
        RECT 2650.930 2477.090 2652.110 2478.270 ;
        RECT 2650.930 2475.490 2652.110 2476.670 ;
        RECT 2650.930 2297.090 2652.110 2298.270 ;
        RECT 2650.930 2295.490 2652.110 2296.670 ;
        RECT 2650.930 2117.090 2652.110 2118.270 ;
        RECT 2650.930 2115.490 2652.110 2116.670 ;
        RECT 2650.930 1937.090 2652.110 1938.270 ;
        RECT 2650.930 1935.490 2652.110 1936.670 ;
        RECT 2650.930 1757.090 2652.110 1758.270 ;
        RECT 2650.930 1755.490 2652.110 1756.670 ;
        RECT 2650.930 1577.090 2652.110 1578.270 ;
        RECT 2650.930 1575.490 2652.110 1576.670 ;
        RECT 2650.930 1397.090 2652.110 1398.270 ;
        RECT 2650.930 1395.490 2652.110 1396.670 ;
        RECT 2650.930 1217.090 2652.110 1218.270 ;
        RECT 2650.930 1215.490 2652.110 1216.670 ;
        RECT 2650.930 1037.090 2652.110 1038.270 ;
        RECT 2650.930 1035.490 2652.110 1036.670 ;
        RECT 2650.930 857.090 2652.110 858.270 ;
        RECT 2650.930 855.490 2652.110 856.670 ;
        RECT 2650.930 677.090 2652.110 678.270 ;
        RECT 2650.930 675.490 2652.110 676.670 ;
        RECT 2650.930 497.090 2652.110 498.270 ;
        RECT 2650.930 495.490 2652.110 496.670 ;
        RECT 2650.930 317.090 2652.110 318.270 ;
        RECT 2650.930 315.490 2652.110 316.670 ;
        RECT 2650.930 137.090 2652.110 138.270 ;
        RECT 2650.930 135.490 2652.110 136.670 ;
        RECT 2650.930 -25.910 2652.110 -24.730 ;
        RECT 2650.930 -27.510 2652.110 -26.330 ;
        RECT 2830.930 3546.010 2832.110 3547.190 ;
        RECT 2830.930 3544.410 2832.110 3545.590 ;
        RECT 2830.930 3377.090 2832.110 3378.270 ;
        RECT 2830.930 3375.490 2832.110 3376.670 ;
        RECT 2830.930 3197.090 2832.110 3198.270 ;
        RECT 2830.930 3195.490 2832.110 3196.670 ;
        RECT 2830.930 3017.090 2832.110 3018.270 ;
        RECT 2830.930 3015.490 2832.110 3016.670 ;
        RECT 2830.930 2837.090 2832.110 2838.270 ;
        RECT 2830.930 2835.490 2832.110 2836.670 ;
        RECT 2830.930 2657.090 2832.110 2658.270 ;
        RECT 2830.930 2655.490 2832.110 2656.670 ;
        RECT 2830.930 2477.090 2832.110 2478.270 ;
        RECT 2830.930 2475.490 2832.110 2476.670 ;
        RECT 2830.930 2297.090 2832.110 2298.270 ;
        RECT 2830.930 2295.490 2832.110 2296.670 ;
        RECT 2830.930 2117.090 2832.110 2118.270 ;
        RECT 2830.930 2115.490 2832.110 2116.670 ;
        RECT 2830.930 1937.090 2832.110 1938.270 ;
        RECT 2830.930 1935.490 2832.110 1936.670 ;
        RECT 2830.930 1757.090 2832.110 1758.270 ;
        RECT 2830.930 1755.490 2832.110 1756.670 ;
        RECT 2830.930 1577.090 2832.110 1578.270 ;
        RECT 2830.930 1575.490 2832.110 1576.670 ;
        RECT 2830.930 1397.090 2832.110 1398.270 ;
        RECT 2830.930 1395.490 2832.110 1396.670 ;
        RECT 2830.930 1217.090 2832.110 1218.270 ;
        RECT 2830.930 1215.490 2832.110 1216.670 ;
        RECT 2830.930 1037.090 2832.110 1038.270 ;
        RECT 2830.930 1035.490 2832.110 1036.670 ;
        RECT 2830.930 857.090 2832.110 858.270 ;
        RECT 2830.930 855.490 2832.110 856.670 ;
        RECT 2830.930 677.090 2832.110 678.270 ;
        RECT 2830.930 675.490 2832.110 676.670 ;
        RECT 2830.930 497.090 2832.110 498.270 ;
        RECT 2830.930 495.490 2832.110 496.670 ;
        RECT 2830.930 317.090 2832.110 318.270 ;
        RECT 2830.930 315.490 2832.110 316.670 ;
        RECT 2830.930 137.090 2832.110 138.270 ;
        RECT 2830.930 135.490 2832.110 136.670 ;
        RECT 2830.930 -25.910 2832.110 -24.730 ;
        RECT 2830.930 -27.510 2832.110 -26.330 ;
        RECT 2950.510 3546.010 2951.690 3547.190 ;
        RECT 2950.510 3544.410 2951.690 3545.590 ;
        RECT 2950.510 3377.090 2951.690 3378.270 ;
        RECT 2950.510 3375.490 2951.690 3376.670 ;
        RECT 2950.510 3197.090 2951.690 3198.270 ;
        RECT 2950.510 3195.490 2951.690 3196.670 ;
        RECT 2950.510 3017.090 2951.690 3018.270 ;
        RECT 2950.510 3015.490 2951.690 3016.670 ;
        RECT 2950.510 2837.090 2951.690 2838.270 ;
        RECT 2950.510 2835.490 2951.690 2836.670 ;
        RECT 2950.510 2657.090 2951.690 2658.270 ;
        RECT 2950.510 2655.490 2951.690 2656.670 ;
        RECT 2950.510 2477.090 2951.690 2478.270 ;
        RECT 2950.510 2475.490 2951.690 2476.670 ;
        RECT 2950.510 2297.090 2951.690 2298.270 ;
        RECT 2950.510 2295.490 2951.690 2296.670 ;
        RECT 2950.510 2117.090 2951.690 2118.270 ;
        RECT 2950.510 2115.490 2951.690 2116.670 ;
        RECT 2950.510 1937.090 2951.690 1938.270 ;
        RECT 2950.510 1935.490 2951.690 1936.670 ;
        RECT 2950.510 1757.090 2951.690 1758.270 ;
        RECT 2950.510 1755.490 2951.690 1756.670 ;
        RECT 2950.510 1577.090 2951.690 1578.270 ;
        RECT 2950.510 1575.490 2951.690 1576.670 ;
        RECT 2950.510 1397.090 2951.690 1398.270 ;
        RECT 2950.510 1395.490 2951.690 1396.670 ;
        RECT 2950.510 1217.090 2951.690 1218.270 ;
        RECT 2950.510 1215.490 2951.690 1216.670 ;
        RECT 2950.510 1037.090 2951.690 1038.270 ;
        RECT 2950.510 1035.490 2951.690 1036.670 ;
        RECT 2950.510 857.090 2951.690 858.270 ;
        RECT 2950.510 855.490 2951.690 856.670 ;
        RECT 2950.510 677.090 2951.690 678.270 ;
        RECT 2950.510 675.490 2951.690 676.670 ;
        RECT 2950.510 497.090 2951.690 498.270 ;
        RECT 2950.510 495.490 2951.690 496.670 ;
        RECT 2950.510 317.090 2951.690 318.270 ;
        RECT 2950.510 315.490 2951.690 316.670 ;
        RECT 2950.510 137.090 2951.690 138.270 ;
        RECT 2950.510 135.490 2951.690 136.670 ;
        RECT 2950.510 -25.910 2951.690 -24.730 ;
        RECT 2950.510 -27.510 2951.690 -26.330 ;
      LAYER met5 ;
        RECT -32.980 3547.300 -29.980 3547.310 ;
        RECT 130.020 3547.300 133.020 3547.310 ;
        RECT 310.020 3547.300 313.020 3547.310 ;
        RECT 490.020 3547.300 493.020 3547.310 ;
        RECT 670.020 3547.300 673.020 3547.310 ;
        RECT 850.020 3547.300 853.020 3547.310 ;
        RECT 1030.020 3547.300 1033.020 3547.310 ;
        RECT 1210.020 3547.300 1213.020 3547.310 ;
        RECT 1390.020 3547.300 1393.020 3547.310 ;
        RECT 1570.020 3547.300 1573.020 3547.310 ;
        RECT 1750.020 3547.300 1753.020 3547.310 ;
        RECT 1930.020 3547.300 1933.020 3547.310 ;
        RECT 2110.020 3547.300 2113.020 3547.310 ;
        RECT 2290.020 3547.300 2293.020 3547.310 ;
        RECT 2470.020 3547.300 2473.020 3547.310 ;
        RECT 2650.020 3547.300 2653.020 3547.310 ;
        RECT 2830.020 3547.300 2833.020 3547.310 ;
        RECT 2949.600 3547.300 2952.600 3547.310 ;
        RECT -32.980 3544.300 2952.600 3547.300 ;
        RECT -32.980 3544.290 -29.980 3544.300 ;
        RECT 130.020 3544.290 133.020 3544.300 ;
        RECT 310.020 3544.290 313.020 3544.300 ;
        RECT 490.020 3544.290 493.020 3544.300 ;
        RECT 670.020 3544.290 673.020 3544.300 ;
        RECT 850.020 3544.290 853.020 3544.300 ;
        RECT 1030.020 3544.290 1033.020 3544.300 ;
        RECT 1210.020 3544.290 1213.020 3544.300 ;
        RECT 1390.020 3544.290 1393.020 3544.300 ;
        RECT 1570.020 3544.290 1573.020 3544.300 ;
        RECT 1750.020 3544.290 1753.020 3544.300 ;
        RECT 1930.020 3544.290 1933.020 3544.300 ;
        RECT 2110.020 3544.290 2113.020 3544.300 ;
        RECT 2290.020 3544.290 2293.020 3544.300 ;
        RECT 2470.020 3544.290 2473.020 3544.300 ;
        RECT 2650.020 3544.290 2653.020 3544.300 ;
        RECT 2830.020 3544.290 2833.020 3544.300 ;
        RECT 2949.600 3544.290 2952.600 3544.300 ;
        RECT -32.980 3378.380 -29.980 3378.390 ;
        RECT 130.020 3378.380 133.020 3378.390 ;
        RECT 310.020 3378.380 313.020 3378.390 ;
        RECT 490.020 3378.380 493.020 3378.390 ;
        RECT 670.020 3378.380 673.020 3378.390 ;
        RECT 850.020 3378.380 853.020 3378.390 ;
        RECT 1030.020 3378.380 1033.020 3378.390 ;
        RECT 1210.020 3378.380 1213.020 3378.390 ;
        RECT 1390.020 3378.380 1393.020 3378.390 ;
        RECT 1570.020 3378.380 1573.020 3378.390 ;
        RECT 1750.020 3378.380 1753.020 3378.390 ;
        RECT 1930.020 3378.380 1933.020 3378.390 ;
        RECT 2110.020 3378.380 2113.020 3378.390 ;
        RECT 2290.020 3378.380 2293.020 3378.390 ;
        RECT 2470.020 3378.380 2473.020 3378.390 ;
        RECT 2650.020 3378.380 2653.020 3378.390 ;
        RECT 2830.020 3378.380 2833.020 3378.390 ;
        RECT 2949.600 3378.380 2952.600 3378.390 ;
        RECT -32.980 3375.380 2952.600 3378.380 ;
        RECT -32.980 3375.370 -29.980 3375.380 ;
        RECT 130.020 3375.370 133.020 3375.380 ;
        RECT 310.020 3375.370 313.020 3375.380 ;
        RECT 490.020 3375.370 493.020 3375.380 ;
        RECT 670.020 3375.370 673.020 3375.380 ;
        RECT 850.020 3375.370 853.020 3375.380 ;
        RECT 1030.020 3375.370 1033.020 3375.380 ;
        RECT 1210.020 3375.370 1213.020 3375.380 ;
        RECT 1390.020 3375.370 1393.020 3375.380 ;
        RECT 1570.020 3375.370 1573.020 3375.380 ;
        RECT 1750.020 3375.370 1753.020 3375.380 ;
        RECT 1930.020 3375.370 1933.020 3375.380 ;
        RECT 2110.020 3375.370 2113.020 3375.380 ;
        RECT 2290.020 3375.370 2293.020 3375.380 ;
        RECT 2470.020 3375.370 2473.020 3375.380 ;
        RECT 2650.020 3375.370 2653.020 3375.380 ;
        RECT 2830.020 3375.370 2833.020 3375.380 ;
        RECT 2949.600 3375.370 2952.600 3375.380 ;
        RECT -32.980 3198.380 -29.980 3198.390 ;
        RECT 130.020 3198.380 133.020 3198.390 ;
        RECT 310.020 3198.380 313.020 3198.390 ;
        RECT 490.020 3198.380 493.020 3198.390 ;
        RECT 670.020 3198.380 673.020 3198.390 ;
        RECT 850.020 3198.380 853.020 3198.390 ;
        RECT 1030.020 3198.380 1033.020 3198.390 ;
        RECT 1210.020 3198.380 1213.020 3198.390 ;
        RECT 1390.020 3198.380 1393.020 3198.390 ;
        RECT 1570.020 3198.380 1573.020 3198.390 ;
        RECT 1750.020 3198.380 1753.020 3198.390 ;
        RECT 1930.020 3198.380 1933.020 3198.390 ;
        RECT 2110.020 3198.380 2113.020 3198.390 ;
        RECT 2290.020 3198.380 2293.020 3198.390 ;
        RECT 2470.020 3198.380 2473.020 3198.390 ;
        RECT 2650.020 3198.380 2653.020 3198.390 ;
        RECT 2830.020 3198.380 2833.020 3198.390 ;
        RECT 2949.600 3198.380 2952.600 3198.390 ;
        RECT -32.980 3195.380 2952.600 3198.380 ;
        RECT -32.980 3195.370 -29.980 3195.380 ;
        RECT 130.020 3195.370 133.020 3195.380 ;
        RECT 310.020 3195.370 313.020 3195.380 ;
        RECT 490.020 3195.370 493.020 3195.380 ;
        RECT 670.020 3195.370 673.020 3195.380 ;
        RECT 850.020 3195.370 853.020 3195.380 ;
        RECT 1030.020 3195.370 1033.020 3195.380 ;
        RECT 1210.020 3195.370 1213.020 3195.380 ;
        RECT 1390.020 3195.370 1393.020 3195.380 ;
        RECT 1570.020 3195.370 1573.020 3195.380 ;
        RECT 1750.020 3195.370 1753.020 3195.380 ;
        RECT 1930.020 3195.370 1933.020 3195.380 ;
        RECT 2110.020 3195.370 2113.020 3195.380 ;
        RECT 2290.020 3195.370 2293.020 3195.380 ;
        RECT 2470.020 3195.370 2473.020 3195.380 ;
        RECT 2650.020 3195.370 2653.020 3195.380 ;
        RECT 2830.020 3195.370 2833.020 3195.380 ;
        RECT 2949.600 3195.370 2952.600 3195.380 ;
        RECT -32.980 3018.380 -29.980 3018.390 ;
        RECT 130.020 3018.380 133.020 3018.390 ;
        RECT 310.020 3018.380 313.020 3018.390 ;
        RECT 490.020 3018.380 493.020 3018.390 ;
        RECT 670.020 3018.380 673.020 3018.390 ;
        RECT 850.020 3018.380 853.020 3018.390 ;
        RECT 1030.020 3018.380 1033.020 3018.390 ;
        RECT 1210.020 3018.380 1213.020 3018.390 ;
        RECT 1390.020 3018.380 1393.020 3018.390 ;
        RECT 1570.020 3018.380 1573.020 3018.390 ;
        RECT 1750.020 3018.380 1753.020 3018.390 ;
        RECT 1930.020 3018.380 1933.020 3018.390 ;
        RECT 2110.020 3018.380 2113.020 3018.390 ;
        RECT 2290.020 3018.380 2293.020 3018.390 ;
        RECT 2470.020 3018.380 2473.020 3018.390 ;
        RECT 2650.020 3018.380 2653.020 3018.390 ;
        RECT 2830.020 3018.380 2833.020 3018.390 ;
        RECT 2949.600 3018.380 2952.600 3018.390 ;
        RECT -32.980 3015.380 2952.600 3018.380 ;
        RECT -32.980 3015.370 -29.980 3015.380 ;
        RECT 130.020 3015.370 133.020 3015.380 ;
        RECT 310.020 3015.370 313.020 3015.380 ;
        RECT 490.020 3015.370 493.020 3015.380 ;
        RECT 670.020 3015.370 673.020 3015.380 ;
        RECT 850.020 3015.370 853.020 3015.380 ;
        RECT 1030.020 3015.370 1033.020 3015.380 ;
        RECT 1210.020 3015.370 1213.020 3015.380 ;
        RECT 1390.020 3015.370 1393.020 3015.380 ;
        RECT 1570.020 3015.370 1573.020 3015.380 ;
        RECT 1750.020 3015.370 1753.020 3015.380 ;
        RECT 1930.020 3015.370 1933.020 3015.380 ;
        RECT 2110.020 3015.370 2113.020 3015.380 ;
        RECT 2290.020 3015.370 2293.020 3015.380 ;
        RECT 2470.020 3015.370 2473.020 3015.380 ;
        RECT 2650.020 3015.370 2653.020 3015.380 ;
        RECT 2830.020 3015.370 2833.020 3015.380 ;
        RECT 2949.600 3015.370 2952.600 3015.380 ;
        RECT -32.980 2838.380 -29.980 2838.390 ;
        RECT 130.020 2838.380 133.020 2838.390 ;
        RECT 310.020 2838.380 313.020 2838.390 ;
        RECT 490.020 2838.380 493.020 2838.390 ;
        RECT 670.020 2838.380 673.020 2838.390 ;
        RECT 850.020 2838.380 853.020 2838.390 ;
        RECT 1030.020 2838.380 1033.020 2838.390 ;
        RECT 1210.020 2838.380 1213.020 2838.390 ;
        RECT 1390.020 2838.380 1393.020 2838.390 ;
        RECT 1570.020 2838.380 1573.020 2838.390 ;
        RECT 1750.020 2838.380 1753.020 2838.390 ;
        RECT 1930.020 2838.380 1933.020 2838.390 ;
        RECT 2110.020 2838.380 2113.020 2838.390 ;
        RECT 2290.020 2838.380 2293.020 2838.390 ;
        RECT 2470.020 2838.380 2473.020 2838.390 ;
        RECT 2650.020 2838.380 2653.020 2838.390 ;
        RECT 2830.020 2838.380 2833.020 2838.390 ;
        RECT 2949.600 2838.380 2952.600 2838.390 ;
        RECT -32.980 2835.380 2952.600 2838.380 ;
        RECT -32.980 2835.370 -29.980 2835.380 ;
        RECT 130.020 2835.370 133.020 2835.380 ;
        RECT 310.020 2835.370 313.020 2835.380 ;
        RECT 490.020 2835.370 493.020 2835.380 ;
        RECT 670.020 2835.370 673.020 2835.380 ;
        RECT 850.020 2835.370 853.020 2835.380 ;
        RECT 1030.020 2835.370 1033.020 2835.380 ;
        RECT 1210.020 2835.370 1213.020 2835.380 ;
        RECT 1390.020 2835.370 1393.020 2835.380 ;
        RECT 1570.020 2835.370 1573.020 2835.380 ;
        RECT 1750.020 2835.370 1753.020 2835.380 ;
        RECT 1930.020 2835.370 1933.020 2835.380 ;
        RECT 2110.020 2835.370 2113.020 2835.380 ;
        RECT 2290.020 2835.370 2293.020 2835.380 ;
        RECT 2470.020 2835.370 2473.020 2835.380 ;
        RECT 2650.020 2835.370 2653.020 2835.380 ;
        RECT 2830.020 2835.370 2833.020 2835.380 ;
        RECT 2949.600 2835.370 2952.600 2835.380 ;
        RECT -32.980 2658.380 -29.980 2658.390 ;
        RECT 130.020 2658.380 133.020 2658.390 ;
        RECT 310.020 2658.380 313.020 2658.390 ;
        RECT 490.020 2658.380 493.020 2658.390 ;
        RECT 670.020 2658.380 673.020 2658.390 ;
        RECT 850.020 2658.380 853.020 2658.390 ;
        RECT 1030.020 2658.380 1033.020 2658.390 ;
        RECT 1210.020 2658.380 1213.020 2658.390 ;
        RECT 1390.020 2658.380 1393.020 2658.390 ;
        RECT 1570.020 2658.380 1573.020 2658.390 ;
        RECT 1750.020 2658.380 1753.020 2658.390 ;
        RECT 1930.020 2658.380 1933.020 2658.390 ;
        RECT 2110.020 2658.380 2113.020 2658.390 ;
        RECT 2290.020 2658.380 2293.020 2658.390 ;
        RECT 2470.020 2658.380 2473.020 2658.390 ;
        RECT 2650.020 2658.380 2653.020 2658.390 ;
        RECT 2830.020 2658.380 2833.020 2658.390 ;
        RECT 2949.600 2658.380 2952.600 2658.390 ;
        RECT -32.980 2655.380 2952.600 2658.380 ;
        RECT -32.980 2655.370 -29.980 2655.380 ;
        RECT 130.020 2655.370 133.020 2655.380 ;
        RECT 310.020 2655.370 313.020 2655.380 ;
        RECT 490.020 2655.370 493.020 2655.380 ;
        RECT 670.020 2655.370 673.020 2655.380 ;
        RECT 850.020 2655.370 853.020 2655.380 ;
        RECT 1030.020 2655.370 1033.020 2655.380 ;
        RECT 1210.020 2655.370 1213.020 2655.380 ;
        RECT 1390.020 2655.370 1393.020 2655.380 ;
        RECT 1570.020 2655.370 1573.020 2655.380 ;
        RECT 1750.020 2655.370 1753.020 2655.380 ;
        RECT 1930.020 2655.370 1933.020 2655.380 ;
        RECT 2110.020 2655.370 2113.020 2655.380 ;
        RECT 2290.020 2655.370 2293.020 2655.380 ;
        RECT 2470.020 2655.370 2473.020 2655.380 ;
        RECT 2650.020 2655.370 2653.020 2655.380 ;
        RECT 2830.020 2655.370 2833.020 2655.380 ;
        RECT 2949.600 2655.370 2952.600 2655.380 ;
        RECT -32.980 2478.380 -29.980 2478.390 ;
        RECT 130.020 2478.380 133.020 2478.390 ;
        RECT 310.020 2478.380 313.020 2478.390 ;
        RECT 490.020 2478.380 493.020 2478.390 ;
        RECT 670.020 2478.380 673.020 2478.390 ;
        RECT 850.020 2478.380 853.020 2478.390 ;
        RECT 1030.020 2478.380 1033.020 2478.390 ;
        RECT 1210.020 2478.380 1213.020 2478.390 ;
        RECT 1390.020 2478.380 1393.020 2478.390 ;
        RECT 1570.020 2478.380 1573.020 2478.390 ;
        RECT 1750.020 2478.380 1753.020 2478.390 ;
        RECT 1930.020 2478.380 1933.020 2478.390 ;
        RECT 2110.020 2478.380 2113.020 2478.390 ;
        RECT 2290.020 2478.380 2293.020 2478.390 ;
        RECT 2470.020 2478.380 2473.020 2478.390 ;
        RECT 2650.020 2478.380 2653.020 2478.390 ;
        RECT 2830.020 2478.380 2833.020 2478.390 ;
        RECT 2949.600 2478.380 2952.600 2478.390 ;
        RECT -32.980 2475.380 2952.600 2478.380 ;
        RECT -32.980 2475.370 -29.980 2475.380 ;
        RECT 130.020 2475.370 133.020 2475.380 ;
        RECT 310.020 2475.370 313.020 2475.380 ;
        RECT 490.020 2475.370 493.020 2475.380 ;
        RECT 670.020 2475.370 673.020 2475.380 ;
        RECT 850.020 2475.370 853.020 2475.380 ;
        RECT 1030.020 2475.370 1033.020 2475.380 ;
        RECT 1210.020 2475.370 1213.020 2475.380 ;
        RECT 1390.020 2475.370 1393.020 2475.380 ;
        RECT 1570.020 2475.370 1573.020 2475.380 ;
        RECT 1750.020 2475.370 1753.020 2475.380 ;
        RECT 1930.020 2475.370 1933.020 2475.380 ;
        RECT 2110.020 2475.370 2113.020 2475.380 ;
        RECT 2290.020 2475.370 2293.020 2475.380 ;
        RECT 2470.020 2475.370 2473.020 2475.380 ;
        RECT 2650.020 2475.370 2653.020 2475.380 ;
        RECT 2830.020 2475.370 2833.020 2475.380 ;
        RECT 2949.600 2475.370 2952.600 2475.380 ;
        RECT -32.980 2298.380 -29.980 2298.390 ;
        RECT 130.020 2298.380 133.020 2298.390 ;
        RECT 310.020 2298.380 313.020 2298.390 ;
        RECT 490.020 2298.380 493.020 2298.390 ;
        RECT 670.020 2298.380 673.020 2298.390 ;
        RECT 850.020 2298.380 853.020 2298.390 ;
        RECT 1030.020 2298.380 1033.020 2298.390 ;
        RECT 1210.020 2298.380 1213.020 2298.390 ;
        RECT 1390.020 2298.380 1393.020 2298.390 ;
        RECT 1570.020 2298.380 1573.020 2298.390 ;
        RECT 1750.020 2298.380 1753.020 2298.390 ;
        RECT 1930.020 2298.380 1933.020 2298.390 ;
        RECT 2110.020 2298.380 2113.020 2298.390 ;
        RECT 2290.020 2298.380 2293.020 2298.390 ;
        RECT 2470.020 2298.380 2473.020 2298.390 ;
        RECT 2650.020 2298.380 2653.020 2298.390 ;
        RECT 2830.020 2298.380 2833.020 2298.390 ;
        RECT 2949.600 2298.380 2952.600 2298.390 ;
        RECT -32.980 2295.380 2952.600 2298.380 ;
        RECT -32.980 2295.370 -29.980 2295.380 ;
        RECT 130.020 2295.370 133.020 2295.380 ;
        RECT 310.020 2295.370 313.020 2295.380 ;
        RECT 490.020 2295.370 493.020 2295.380 ;
        RECT 670.020 2295.370 673.020 2295.380 ;
        RECT 850.020 2295.370 853.020 2295.380 ;
        RECT 1030.020 2295.370 1033.020 2295.380 ;
        RECT 1210.020 2295.370 1213.020 2295.380 ;
        RECT 1390.020 2295.370 1393.020 2295.380 ;
        RECT 1570.020 2295.370 1573.020 2295.380 ;
        RECT 1750.020 2295.370 1753.020 2295.380 ;
        RECT 1930.020 2295.370 1933.020 2295.380 ;
        RECT 2110.020 2295.370 2113.020 2295.380 ;
        RECT 2290.020 2295.370 2293.020 2295.380 ;
        RECT 2470.020 2295.370 2473.020 2295.380 ;
        RECT 2650.020 2295.370 2653.020 2295.380 ;
        RECT 2830.020 2295.370 2833.020 2295.380 ;
        RECT 2949.600 2295.370 2952.600 2295.380 ;
        RECT -32.980 2118.380 -29.980 2118.390 ;
        RECT 130.020 2118.380 133.020 2118.390 ;
        RECT 310.020 2118.380 313.020 2118.390 ;
        RECT 490.020 2118.380 493.020 2118.390 ;
        RECT 670.020 2118.380 673.020 2118.390 ;
        RECT 850.020 2118.380 853.020 2118.390 ;
        RECT 1030.020 2118.380 1033.020 2118.390 ;
        RECT 1210.020 2118.380 1213.020 2118.390 ;
        RECT 1390.020 2118.380 1393.020 2118.390 ;
        RECT 1570.020 2118.380 1573.020 2118.390 ;
        RECT 1750.020 2118.380 1753.020 2118.390 ;
        RECT 1930.020 2118.380 1933.020 2118.390 ;
        RECT 2110.020 2118.380 2113.020 2118.390 ;
        RECT 2290.020 2118.380 2293.020 2118.390 ;
        RECT 2470.020 2118.380 2473.020 2118.390 ;
        RECT 2650.020 2118.380 2653.020 2118.390 ;
        RECT 2830.020 2118.380 2833.020 2118.390 ;
        RECT 2949.600 2118.380 2952.600 2118.390 ;
        RECT -32.980 2115.380 2952.600 2118.380 ;
        RECT -32.980 2115.370 -29.980 2115.380 ;
        RECT 130.020 2115.370 133.020 2115.380 ;
        RECT 310.020 2115.370 313.020 2115.380 ;
        RECT 490.020 2115.370 493.020 2115.380 ;
        RECT 670.020 2115.370 673.020 2115.380 ;
        RECT 850.020 2115.370 853.020 2115.380 ;
        RECT 1030.020 2115.370 1033.020 2115.380 ;
        RECT 1210.020 2115.370 1213.020 2115.380 ;
        RECT 1390.020 2115.370 1393.020 2115.380 ;
        RECT 1570.020 2115.370 1573.020 2115.380 ;
        RECT 1750.020 2115.370 1753.020 2115.380 ;
        RECT 1930.020 2115.370 1933.020 2115.380 ;
        RECT 2110.020 2115.370 2113.020 2115.380 ;
        RECT 2290.020 2115.370 2293.020 2115.380 ;
        RECT 2470.020 2115.370 2473.020 2115.380 ;
        RECT 2650.020 2115.370 2653.020 2115.380 ;
        RECT 2830.020 2115.370 2833.020 2115.380 ;
        RECT 2949.600 2115.370 2952.600 2115.380 ;
        RECT -32.980 1938.380 -29.980 1938.390 ;
        RECT 130.020 1938.380 133.020 1938.390 ;
        RECT 310.020 1938.380 313.020 1938.390 ;
        RECT 490.020 1938.380 493.020 1938.390 ;
        RECT 670.020 1938.380 673.020 1938.390 ;
        RECT 850.020 1938.380 853.020 1938.390 ;
        RECT 1030.020 1938.380 1033.020 1938.390 ;
        RECT 1210.020 1938.380 1213.020 1938.390 ;
        RECT 1390.020 1938.380 1393.020 1938.390 ;
        RECT 1570.020 1938.380 1573.020 1938.390 ;
        RECT 1750.020 1938.380 1753.020 1938.390 ;
        RECT 1930.020 1938.380 1933.020 1938.390 ;
        RECT 2110.020 1938.380 2113.020 1938.390 ;
        RECT 2290.020 1938.380 2293.020 1938.390 ;
        RECT 2470.020 1938.380 2473.020 1938.390 ;
        RECT 2650.020 1938.380 2653.020 1938.390 ;
        RECT 2830.020 1938.380 2833.020 1938.390 ;
        RECT 2949.600 1938.380 2952.600 1938.390 ;
        RECT -32.980 1935.380 2952.600 1938.380 ;
        RECT -32.980 1935.370 -29.980 1935.380 ;
        RECT 130.020 1935.370 133.020 1935.380 ;
        RECT 310.020 1935.370 313.020 1935.380 ;
        RECT 490.020 1935.370 493.020 1935.380 ;
        RECT 670.020 1935.370 673.020 1935.380 ;
        RECT 850.020 1935.370 853.020 1935.380 ;
        RECT 1030.020 1935.370 1033.020 1935.380 ;
        RECT 1210.020 1935.370 1213.020 1935.380 ;
        RECT 1390.020 1935.370 1393.020 1935.380 ;
        RECT 1570.020 1935.370 1573.020 1935.380 ;
        RECT 1750.020 1935.370 1753.020 1935.380 ;
        RECT 1930.020 1935.370 1933.020 1935.380 ;
        RECT 2110.020 1935.370 2113.020 1935.380 ;
        RECT 2290.020 1935.370 2293.020 1935.380 ;
        RECT 2470.020 1935.370 2473.020 1935.380 ;
        RECT 2650.020 1935.370 2653.020 1935.380 ;
        RECT 2830.020 1935.370 2833.020 1935.380 ;
        RECT 2949.600 1935.370 2952.600 1935.380 ;
        RECT -32.980 1758.380 -29.980 1758.390 ;
        RECT 130.020 1758.380 133.020 1758.390 ;
        RECT 310.020 1758.380 313.020 1758.390 ;
        RECT 490.020 1758.380 493.020 1758.390 ;
        RECT 670.020 1758.380 673.020 1758.390 ;
        RECT 850.020 1758.380 853.020 1758.390 ;
        RECT 1030.020 1758.380 1033.020 1758.390 ;
        RECT 1210.020 1758.380 1213.020 1758.390 ;
        RECT 1390.020 1758.380 1393.020 1758.390 ;
        RECT 1570.020 1758.380 1573.020 1758.390 ;
        RECT 1750.020 1758.380 1753.020 1758.390 ;
        RECT 1930.020 1758.380 1933.020 1758.390 ;
        RECT 2110.020 1758.380 2113.020 1758.390 ;
        RECT 2290.020 1758.380 2293.020 1758.390 ;
        RECT 2470.020 1758.380 2473.020 1758.390 ;
        RECT 2650.020 1758.380 2653.020 1758.390 ;
        RECT 2830.020 1758.380 2833.020 1758.390 ;
        RECT 2949.600 1758.380 2952.600 1758.390 ;
        RECT -32.980 1755.380 2952.600 1758.380 ;
        RECT -32.980 1755.370 -29.980 1755.380 ;
        RECT 130.020 1755.370 133.020 1755.380 ;
        RECT 310.020 1755.370 313.020 1755.380 ;
        RECT 490.020 1755.370 493.020 1755.380 ;
        RECT 670.020 1755.370 673.020 1755.380 ;
        RECT 850.020 1755.370 853.020 1755.380 ;
        RECT 1030.020 1755.370 1033.020 1755.380 ;
        RECT 1210.020 1755.370 1213.020 1755.380 ;
        RECT 1390.020 1755.370 1393.020 1755.380 ;
        RECT 1570.020 1755.370 1573.020 1755.380 ;
        RECT 1750.020 1755.370 1753.020 1755.380 ;
        RECT 1930.020 1755.370 1933.020 1755.380 ;
        RECT 2110.020 1755.370 2113.020 1755.380 ;
        RECT 2290.020 1755.370 2293.020 1755.380 ;
        RECT 2470.020 1755.370 2473.020 1755.380 ;
        RECT 2650.020 1755.370 2653.020 1755.380 ;
        RECT 2830.020 1755.370 2833.020 1755.380 ;
        RECT 2949.600 1755.370 2952.600 1755.380 ;
        RECT -32.980 1578.380 -29.980 1578.390 ;
        RECT 130.020 1578.380 133.020 1578.390 ;
        RECT 310.020 1578.380 313.020 1578.390 ;
        RECT 490.020 1578.380 493.020 1578.390 ;
        RECT 670.020 1578.380 673.020 1578.390 ;
        RECT 850.020 1578.380 853.020 1578.390 ;
        RECT 1030.020 1578.380 1033.020 1578.390 ;
        RECT 1210.020 1578.380 1213.020 1578.390 ;
        RECT 1390.020 1578.380 1393.020 1578.390 ;
        RECT 1570.020 1578.380 1573.020 1578.390 ;
        RECT 1750.020 1578.380 1753.020 1578.390 ;
        RECT 1930.020 1578.380 1933.020 1578.390 ;
        RECT 2110.020 1578.380 2113.020 1578.390 ;
        RECT 2290.020 1578.380 2293.020 1578.390 ;
        RECT 2470.020 1578.380 2473.020 1578.390 ;
        RECT 2650.020 1578.380 2653.020 1578.390 ;
        RECT 2830.020 1578.380 2833.020 1578.390 ;
        RECT 2949.600 1578.380 2952.600 1578.390 ;
        RECT -32.980 1575.380 2952.600 1578.380 ;
        RECT -32.980 1575.370 -29.980 1575.380 ;
        RECT 130.020 1575.370 133.020 1575.380 ;
        RECT 310.020 1575.370 313.020 1575.380 ;
        RECT 490.020 1575.370 493.020 1575.380 ;
        RECT 670.020 1575.370 673.020 1575.380 ;
        RECT 850.020 1575.370 853.020 1575.380 ;
        RECT 1030.020 1575.370 1033.020 1575.380 ;
        RECT 1210.020 1575.370 1213.020 1575.380 ;
        RECT 1390.020 1575.370 1393.020 1575.380 ;
        RECT 1570.020 1575.370 1573.020 1575.380 ;
        RECT 1750.020 1575.370 1753.020 1575.380 ;
        RECT 1930.020 1575.370 1933.020 1575.380 ;
        RECT 2110.020 1575.370 2113.020 1575.380 ;
        RECT 2290.020 1575.370 2293.020 1575.380 ;
        RECT 2470.020 1575.370 2473.020 1575.380 ;
        RECT 2650.020 1575.370 2653.020 1575.380 ;
        RECT 2830.020 1575.370 2833.020 1575.380 ;
        RECT 2949.600 1575.370 2952.600 1575.380 ;
        RECT -32.980 1398.380 -29.980 1398.390 ;
        RECT 130.020 1398.380 133.020 1398.390 ;
        RECT 310.020 1398.380 313.020 1398.390 ;
        RECT 490.020 1398.380 493.020 1398.390 ;
        RECT 670.020 1398.380 673.020 1398.390 ;
        RECT 850.020 1398.380 853.020 1398.390 ;
        RECT 1030.020 1398.380 1033.020 1398.390 ;
        RECT 1210.020 1398.380 1213.020 1398.390 ;
        RECT 1390.020 1398.380 1393.020 1398.390 ;
        RECT 1570.020 1398.380 1573.020 1398.390 ;
        RECT 1750.020 1398.380 1753.020 1398.390 ;
        RECT 1930.020 1398.380 1933.020 1398.390 ;
        RECT 2110.020 1398.380 2113.020 1398.390 ;
        RECT 2290.020 1398.380 2293.020 1398.390 ;
        RECT 2470.020 1398.380 2473.020 1398.390 ;
        RECT 2650.020 1398.380 2653.020 1398.390 ;
        RECT 2830.020 1398.380 2833.020 1398.390 ;
        RECT 2949.600 1398.380 2952.600 1398.390 ;
        RECT -32.980 1395.380 2952.600 1398.380 ;
        RECT -32.980 1395.370 -29.980 1395.380 ;
        RECT 130.020 1395.370 133.020 1395.380 ;
        RECT 310.020 1395.370 313.020 1395.380 ;
        RECT 490.020 1395.370 493.020 1395.380 ;
        RECT 670.020 1395.370 673.020 1395.380 ;
        RECT 850.020 1395.370 853.020 1395.380 ;
        RECT 1030.020 1395.370 1033.020 1395.380 ;
        RECT 1210.020 1395.370 1213.020 1395.380 ;
        RECT 1390.020 1395.370 1393.020 1395.380 ;
        RECT 1570.020 1395.370 1573.020 1395.380 ;
        RECT 1750.020 1395.370 1753.020 1395.380 ;
        RECT 1930.020 1395.370 1933.020 1395.380 ;
        RECT 2110.020 1395.370 2113.020 1395.380 ;
        RECT 2290.020 1395.370 2293.020 1395.380 ;
        RECT 2470.020 1395.370 2473.020 1395.380 ;
        RECT 2650.020 1395.370 2653.020 1395.380 ;
        RECT 2830.020 1395.370 2833.020 1395.380 ;
        RECT 2949.600 1395.370 2952.600 1395.380 ;
        RECT -32.980 1218.380 -29.980 1218.390 ;
        RECT 130.020 1218.380 133.020 1218.390 ;
        RECT 310.020 1218.380 313.020 1218.390 ;
        RECT 490.020 1218.380 493.020 1218.390 ;
        RECT 670.020 1218.380 673.020 1218.390 ;
        RECT 850.020 1218.380 853.020 1218.390 ;
        RECT 1030.020 1218.380 1033.020 1218.390 ;
        RECT 1210.020 1218.380 1213.020 1218.390 ;
        RECT 1390.020 1218.380 1393.020 1218.390 ;
        RECT 1570.020 1218.380 1573.020 1218.390 ;
        RECT 1750.020 1218.380 1753.020 1218.390 ;
        RECT 1930.020 1218.380 1933.020 1218.390 ;
        RECT 2110.020 1218.380 2113.020 1218.390 ;
        RECT 2290.020 1218.380 2293.020 1218.390 ;
        RECT 2470.020 1218.380 2473.020 1218.390 ;
        RECT 2650.020 1218.380 2653.020 1218.390 ;
        RECT 2830.020 1218.380 2833.020 1218.390 ;
        RECT 2949.600 1218.380 2952.600 1218.390 ;
        RECT -32.980 1215.380 2952.600 1218.380 ;
        RECT -32.980 1215.370 -29.980 1215.380 ;
        RECT 130.020 1215.370 133.020 1215.380 ;
        RECT 310.020 1215.370 313.020 1215.380 ;
        RECT 490.020 1215.370 493.020 1215.380 ;
        RECT 670.020 1215.370 673.020 1215.380 ;
        RECT 850.020 1215.370 853.020 1215.380 ;
        RECT 1030.020 1215.370 1033.020 1215.380 ;
        RECT 1210.020 1215.370 1213.020 1215.380 ;
        RECT 1390.020 1215.370 1393.020 1215.380 ;
        RECT 1570.020 1215.370 1573.020 1215.380 ;
        RECT 1750.020 1215.370 1753.020 1215.380 ;
        RECT 1930.020 1215.370 1933.020 1215.380 ;
        RECT 2110.020 1215.370 2113.020 1215.380 ;
        RECT 2290.020 1215.370 2293.020 1215.380 ;
        RECT 2470.020 1215.370 2473.020 1215.380 ;
        RECT 2650.020 1215.370 2653.020 1215.380 ;
        RECT 2830.020 1215.370 2833.020 1215.380 ;
        RECT 2949.600 1215.370 2952.600 1215.380 ;
        RECT -32.980 1038.380 -29.980 1038.390 ;
        RECT 130.020 1038.380 133.020 1038.390 ;
        RECT 310.020 1038.380 313.020 1038.390 ;
        RECT 490.020 1038.380 493.020 1038.390 ;
        RECT 670.020 1038.380 673.020 1038.390 ;
        RECT 850.020 1038.380 853.020 1038.390 ;
        RECT 1030.020 1038.380 1033.020 1038.390 ;
        RECT 1210.020 1038.380 1213.020 1038.390 ;
        RECT 1390.020 1038.380 1393.020 1038.390 ;
        RECT 1570.020 1038.380 1573.020 1038.390 ;
        RECT 1750.020 1038.380 1753.020 1038.390 ;
        RECT 1930.020 1038.380 1933.020 1038.390 ;
        RECT 2110.020 1038.380 2113.020 1038.390 ;
        RECT 2290.020 1038.380 2293.020 1038.390 ;
        RECT 2470.020 1038.380 2473.020 1038.390 ;
        RECT 2650.020 1038.380 2653.020 1038.390 ;
        RECT 2830.020 1038.380 2833.020 1038.390 ;
        RECT 2949.600 1038.380 2952.600 1038.390 ;
        RECT -32.980 1035.380 2952.600 1038.380 ;
        RECT -32.980 1035.370 -29.980 1035.380 ;
        RECT 130.020 1035.370 133.020 1035.380 ;
        RECT 310.020 1035.370 313.020 1035.380 ;
        RECT 490.020 1035.370 493.020 1035.380 ;
        RECT 670.020 1035.370 673.020 1035.380 ;
        RECT 850.020 1035.370 853.020 1035.380 ;
        RECT 1030.020 1035.370 1033.020 1035.380 ;
        RECT 1210.020 1035.370 1213.020 1035.380 ;
        RECT 1390.020 1035.370 1393.020 1035.380 ;
        RECT 1570.020 1035.370 1573.020 1035.380 ;
        RECT 1750.020 1035.370 1753.020 1035.380 ;
        RECT 1930.020 1035.370 1933.020 1035.380 ;
        RECT 2110.020 1035.370 2113.020 1035.380 ;
        RECT 2290.020 1035.370 2293.020 1035.380 ;
        RECT 2470.020 1035.370 2473.020 1035.380 ;
        RECT 2650.020 1035.370 2653.020 1035.380 ;
        RECT 2830.020 1035.370 2833.020 1035.380 ;
        RECT 2949.600 1035.370 2952.600 1035.380 ;
        RECT -32.980 858.380 -29.980 858.390 ;
        RECT 130.020 858.380 133.020 858.390 ;
        RECT 310.020 858.380 313.020 858.390 ;
        RECT 490.020 858.380 493.020 858.390 ;
        RECT 670.020 858.380 673.020 858.390 ;
        RECT 850.020 858.380 853.020 858.390 ;
        RECT 1030.020 858.380 1033.020 858.390 ;
        RECT 1210.020 858.380 1213.020 858.390 ;
        RECT 1390.020 858.380 1393.020 858.390 ;
        RECT 1570.020 858.380 1573.020 858.390 ;
        RECT 1750.020 858.380 1753.020 858.390 ;
        RECT 1930.020 858.380 1933.020 858.390 ;
        RECT 2110.020 858.380 2113.020 858.390 ;
        RECT 2290.020 858.380 2293.020 858.390 ;
        RECT 2470.020 858.380 2473.020 858.390 ;
        RECT 2650.020 858.380 2653.020 858.390 ;
        RECT 2830.020 858.380 2833.020 858.390 ;
        RECT 2949.600 858.380 2952.600 858.390 ;
        RECT -32.980 855.380 2952.600 858.380 ;
        RECT -32.980 855.370 -29.980 855.380 ;
        RECT 130.020 855.370 133.020 855.380 ;
        RECT 310.020 855.370 313.020 855.380 ;
        RECT 490.020 855.370 493.020 855.380 ;
        RECT 670.020 855.370 673.020 855.380 ;
        RECT 850.020 855.370 853.020 855.380 ;
        RECT 1030.020 855.370 1033.020 855.380 ;
        RECT 1210.020 855.370 1213.020 855.380 ;
        RECT 1390.020 855.370 1393.020 855.380 ;
        RECT 1570.020 855.370 1573.020 855.380 ;
        RECT 1750.020 855.370 1753.020 855.380 ;
        RECT 1930.020 855.370 1933.020 855.380 ;
        RECT 2110.020 855.370 2113.020 855.380 ;
        RECT 2290.020 855.370 2293.020 855.380 ;
        RECT 2470.020 855.370 2473.020 855.380 ;
        RECT 2650.020 855.370 2653.020 855.380 ;
        RECT 2830.020 855.370 2833.020 855.380 ;
        RECT 2949.600 855.370 2952.600 855.380 ;
        RECT -32.980 678.380 -29.980 678.390 ;
        RECT 130.020 678.380 133.020 678.390 ;
        RECT 310.020 678.380 313.020 678.390 ;
        RECT 490.020 678.380 493.020 678.390 ;
        RECT 670.020 678.380 673.020 678.390 ;
        RECT 850.020 678.380 853.020 678.390 ;
        RECT 1030.020 678.380 1033.020 678.390 ;
        RECT 1210.020 678.380 1213.020 678.390 ;
        RECT 1390.020 678.380 1393.020 678.390 ;
        RECT 1570.020 678.380 1573.020 678.390 ;
        RECT 1750.020 678.380 1753.020 678.390 ;
        RECT 1930.020 678.380 1933.020 678.390 ;
        RECT 2110.020 678.380 2113.020 678.390 ;
        RECT 2290.020 678.380 2293.020 678.390 ;
        RECT 2470.020 678.380 2473.020 678.390 ;
        RECT 2650.020 678.380 2653.020 678.390 ;
        RECT 2830.020 678.380 2833.020 678.390 ;
        RECT 2949.600 678.380 2952.600 678.390 ;
        RECT -32.980 675.380 2952.600 678.380 ;
        RECT -32.980 675.370 -29.980 675.380 ;
        RECT 130.020 675.370 133.020 675.380 ;
        RECT 310.020 675.370 313.020 675.380 ;
        RECT 490.020 675.370 493.020 675.380 ;
        RECT 670.020 675.370 673.020 675.380 ;
        RECT 850.020 675.370 853.020 675.380 ;
        RECT 1030.020 675.370 1033.020 675.380 ;
        RECT 1210.020 675.370 1213.020 675.380 ;
        RECT 1390.020 675.370 1393.020 675.380 ;
        RECT 1570.020 675.370 1573.020 675.380 ;
        RECT 1750.020 675.370 1753.020 675.380 ;
        RECT 1930.020 675.370 1933.020 675.380 ;
        RECT 2110.020 675.370 2113.020 675.380 ;
        RECT 2290.020 675.370 2293.020 675.380 ;
        RECT 2470.020 675.370 2473.020 675.380 ;
        RECT 2650.020 675.370 2653.020 675.380 ;
        RECT 2830.020 675.370 2833.020 675.380 ;
        RECT 2949.600 675.370 2952.600 675.380 ;
        RECT -32.980 498.380 -29.980 498.390 ;
        RECT 130.020 498.380 133.020 498.390 ;
        RECT 310.020 498.380 313.020 498.390 ;
        RECT 490.020 498.380 493.020 498.390 ;
        RECT 670.020 498.380 673.020 498.390 ;
        RECT 850.020 498.380 853.020 498.390 ;
        RECT 1030.020 498.380 1033.020 498.390 ;
        RECT 1210.020 498.380 1213.020 498.390 ;
        RECT 1390.020 498.380 1393.020 498.390 ;
        RECT 1570.020 498.380 1573.020 498.390 ;
        RECT 1750.020 498.380 1753.020 498.390 ;
        RECT 1930.020 498.380 1933.020 498.390 ;
        RECT 2110.020 498.380 2113.020 498.390 ;
        RECT 2290.020 498.380 2293.020 498.390 ;
        RECT 2470.020 498.380 2473.020 498.390 ;
        RECT 2650.020 498.380 2653.020 498.390 ;
        RECT 2830.020 498.380 2833.020 498.390 ;
        RECT 2949.600 498.380 2952.600 498.390 ;
        RECT -32.980 495.380 2952.600 498.380 ;
        RECT -32.980 495.370 -29.980 495.380 ;
        RECT 130.020 495.370 133.020 495.380 ;
        RECT 310.020 495.370 313.020 495.380 ;
        RECT 490.020 495.370 493.020 495.380 ;
        RECT 670.020 495.370 673.020 495.380 ;
        RECT 850.020 495.370 853.020 495.380 ;
        RECT 1030.020 495.370 1033.020 495.380 ;
        RECT 1210.020 495.370 1213.020 495.380 ;
        RECT 1390.020 495.370 1393.020 495.380 ;
        RECT 1570.020 495.370 1573.020 495.380 ;
        RECT 1750.020 495.370 1753.020 495.380 ;
        RECT 1930.020 495.370 1933.020 495.380 ;
        RECT 2110.020 495.370 2113.020 495.380 ;
        RECT 2290.020 495.370 2293.020 495.380 ;
        RECT 2470.020 495.370 2473.020 495.380 ;
        RECT 2650.020 495.370 2653.020 495.380 ;
        RECT 2830.020 495.370 2833.020 495.380 ;
        RECT 2949.600 495.370 2952.600 495.380 ;
        RECT -32.980 318.380 -29.980 318.390 ;
        RECT 130.020 318.380 133.020 318.390 ;
        RECT 310.020 318.380 313.020 318.390 ;
        RECT 490.020 318.380 493.020 318.390 ;
        RECT 670.020 318.380 673.020 318.390 ;
        RECT 850.020 318.380 853.020 318.390 ;
        RECT 1030.020 318.380 1033.020 318.390 ;
        RECT 1210.020 318.380 1213.020 318.390 ;
        RECT 1390.020 318.380 1393.020 318.390 ;
        RECT 1570.020 318.380 1573.020 318.390 ;
        RECT 1750.020 318.380 1753.020 318.390 ;
        RECT 1930.020 318.380 1933.020 318.390 ;
        RECT 2110.020 318.380 2113.020 318.390 ;
        RECT 2290.020 318.380 2293.020 318.390 ;
        RECT 2470.020 318.380 2473.020 318.390 ;
        RECT 2650.020 318.380 2653.020 318.390 ;
        RECT 2830.020 318.380 2833.020 318.390 ;
        RECT 2949.600 318.380 2952.600 318.390 ;
        RECT -32.980 315.380 2952.600 318.380 ;
        RECT -32.980 315.370 -29.980 315.380 ;
        RECT 130.020 315.370 133.020 315.380 ;
        RECT 310.020 315.370 313.020 315.380 ;
        RECT 490.020 315.370 493.020 315.380 ;
        RECT 670.020 315.370 673.020 315.380 ;
        RECT 850.020 315.370 853.020 315.380 ;
        RECT 1030.020 315.370 1033.020 315.380 ;
        RECT 1210.020 315.370 1213.020 315.380 ;
        RECT 1390.020 315.370 1393.020 315.380 ;
        RECT 1570.020 315.370 1573.020 315.380 ;
        RECT 1750.020 315.370 1753.020 315.380 ;
        RECT 1930.020 315.370 1933.020 315.380 ;
        RECT 2110.020 315.370 2113.020 315.380 ;
        RECT 2290.020 315.370 2293.020 315.380 ;
        RECT 2470.020 315.370 2473.020 315.380 ;
        RECT 2650.020 315.370 2653.020 315.380 ;
        RECT 2830.020 315.370 2833.020 315.380 ;
        RECT 2949.600 315.370 2952.600 315.380 ;
        RECT -32.980 138.380 -29.980 138.390 ;
        RECT 130.020 138.380 133.020 138.390 ;
        RECT 310.020 138.380 313.020 138.390 ;
        RECT 490.020 138.380 493.020 138.390 ;
        RECT 670.020 138.380 673.020 138.390 ;
        RECT 850.020 138.380 853.020 138.390 ;
        RECT 1030.020 138.380 1033.020 138.390 ;
        RECT 1210.020 138.380 1213.020 138.390 ;
        RECT 1390.020 138.380 1393.020 138.390 ;
        RECT 1570.020 138.380 1573.020 138.390 ;
        RECT 1750.020 138.380 1753.020 138.390 ;
        RECT 1930.020 138.380 1933.020 138.390 ;
        RECT 2110.020 138.380 2113.020 138.390 ;
        RECT 2290.020 138.380 2293.020 138.390 ;
        RECT 2470.020 138.380 2473.020 138.390 ;
        RECT 2650.020 138.380 2653.020 138.390 ;
        RECT 2830.020 138.380 2833.020 138.390 ;
        RECT 2949.600 138.380 2952.600 138.390 ;
        RECT -32.980 135.380 2952.600 138.380 ;
        RECT -32.980 135.370 -29.980 135.380 ;
        RECT 130.020 135.370 133.020 135.380 ;
        RECT 310.020 135.370 313.020 135.380 ;
        RECT 490.020 135.370 493.020 135.380 ;
        RECT 670.020 135.370 673.020 135.380 ;
        RECT 850.020 135.370 853.020 135.380 ;
        RECT 1030.020 135.370 1033.020 135.380 ;
        RECT 1210.020 135.370 1213.020 135.380 ;
        RECT 1390.020 135.370 1393.020 135.380 ;
        RECT 1570.020 135.370 1573.020 135.380 ;
        RECT 1750.020 135.370 1753.020 135.380 ;
        RECT 1930.020 135.370 1933.020 135.380 ;
        RECT 2110.020 135.370 2113.020 135.380 ;
        RECT 2290.020 135.370 2293.020 135.380 ;
        RECT 2470.020 135.370 2473.020 135.380 ;
        RECT 2650.020 135.370 2653.020 135.380 ;
        RECT 2830.020 135.370 2833.020 135.380 ;
        RECT 2949.600 135.370 2952.600 135.380 ;
        RECT -32.980 -24.620 -29.980 -24.610 ;
        RECT 130.020 -24.620 133.020 -24.610 ;
        RECT 310.020 -24.620 313.020 -24.610 ;
        RECT 490.020 -24.620 493.020 -24.610 ;
        RECT 670.020 -24.620 673.020 -24.610 ;
        RECT 850.020 -24.620 853.020 -24.610 ;
        RECT 1030.020 -24.620 1033.020 -24.610 ;
        RECT 1210.020 -24.620 1213.020 -24.610 ;
        RECT 1390.020 -24.620 1393.020 -24.610 ;
        RECT 1570.020 -24.620 1573.020 -24.610 ;
        RECT 1750.020 -24.620 1753.020 -24.610 ;
        RECT 1930.020 -24.620 1933.020 -24.610 ;
        RECT 2110.020 -24.620 2113.020 -24.610 ;
        RECT 2290.020 -24.620 2293.020 -24.610 ;
        RECT 2470.020 -24.620 2473.020 -24.610 ;
        RECT 2650.020 -24.620 2653.020 -24.610 ;
        RECT 2830.020 -24.620 2833.020 -24.610 ;
        RECT 2949.600 -24.620 2952.600 -24.610 ;
        RECT -32.980 -27.620 2952.600 -24.620 ;
        RECT -32.980 -27.630 -29.980 -27.620 ;
        RECT 130.020 -27.630 133.020 -27.620 ;
        RECT 310.020 -27.630 313.020 -27.620 ;
        RECT 490.020 -27.630 493.020 -27.620 ;
        RECT 670.020 -27.630 673.020 -27.620 ;
        RECT 850.020 -27.630 853.020 -27.620 ;
        RECT 1030.020 -27.630 1033.020 -27.620 ;
        RECT 1210.020 -27.630 1213.020 -27.620 ;
        RECT 1390.020 -27.630 1393.020 -27.620 ;
        RECT 1570.020 -27.630 1573.020 -27.620 ;
        RECT 1750.020 -27.630 1753.020 -27.620 ;
        RECT 1930.020 -27.630 1933.020 -27.620 ;
        RECT 2110.020 -27.630 2113.020 -27.620 ;
        RECT 2290.020 -27.630 2293.020 -27.620 ;
        RECT 2470.020 -27.630 2473.020 -27.620 ;
        RECT 2650.020 -27.630 2653.020 -27.620 ;
        RECT 2830.020 -27.630 2833.020 -27.620 ;
        RECT 2949.600 -27.630 2952.600 -27.620 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -37.580 -32.220 -34.580 3551.900 ;
        RECT 58.020 -36.820 61.020 3556.500 ;
        RECT 238.020 -36.820 241.020 3556.500 ;
        RECT 418.020 -36.820 421.020 3556.500 ;
        RECT 598.020 -36.820 601.020 3556.500 ;
        RECT 778.020 -36.820 781.020 3556.500 ;
        RECT 958.020 -36.820 961.020 3556.500 ;
        RECT 1138.020 -36.820 1141.020 3556.500 ;
        RECT 1318.020 -36.820 1321.020 3556.500 ;
        RECT 1498.020 -36.820 1501.020 3556.500 ;
        RECT 1678.020 -36.820 1681.020 3556.500 ;
        RECT 1858.020 -36.820 1861.020 3556.500 ;
        RECT 2038.020 -36.820 2041.020 3556.500 ;
        RECT 2218.020 -36.820 2221.020 3556.500 ;
        RECT 2398.020 -36.820 2401.020 3556.500 ;
        RECT 2578.020 -36.820 2581.020 3556.500 ;
        RECT 2758.020 -36.820 2761.020 3556.500 ;
        RECT 2954.200 -32.220 2957.200 3551.900 ;
      LAYER via4 ;
        RECT -36.670 3550.610 -35.490 3551.790 ;
        RECT -36.670 3549.010 -35.490 3550.190 ;
        RECT -36.670 3485.090 -35.490 3486.270 ;
        RECT -36.670 3483.490 -35.490 3484.670 ;
        RECT -36.670 3305.090 -35.490 3306.270 ;
        RECT -36.670 3303.490 -35.490 3304.670 ;
        RECT -36.670 3125.090 -35.490 3126.270 ;
        RECT -36.670 3123.490 -35.490 3124.670 ;
        RECT -36.670 2945.090 -35.490 2946.270 ;
        RECT -36.670 2943.490 -35.490 2944.670 ;
        RECT -36.670 2765.090 -35.490 2766.270 ;
        RECT -36.670 2763.490 -35.490 2764.670 ;
        RECT -36.670 2585.090 -35.490 2586.270 ;
        RECT -36.670 2583.490 -35.490 2584.670 ;
        RECT -36.670 2405.090 -35.490 2406.270 ;
        RECT -36.670 2403.490 -35.490 2404.670 ;
        RECT -36.670 2225.090 -35.490 2226.270 ;
        RECT -36.670 2223.490 -35.490 2224.670 ;
        RECT -36.670 2045.090 -35.490 2046.270 ;
        RECT -36.670 2043.490 -35.490 2044.670 ;
        RECT -36.670 1865.090 -35.490 1866.270 ;
        RECT -36.670 1863.490 -35.490 1864.670 ;
        RECT -36.670 1685.090 -35.490 1686.270 ;
        RECT -36.670 1683.490 -35.490 1684.670 ;
        RECT -36.670 1505.090 -35.490 1506.270 ;
        RECT -36.670 1503.490 -35.490 1504.670 ;
        RECT -36.670 1325.090 -35.490 1326.270 ;
        RECT -36.670 1323.490 -35.490 1324.670 ;
        RECT -36.670 1145.090 -35.490 1146.270 ;
        RECT -36.670 1143.490 -35.490 1144.670 ;
        RECT -36.670 965.090 -35.490 966.270 ;
        RECT -36.670 963.490 -35.490 964.670 ;
        RECT -36.670 785.090 -35.490 786.270 ;
        RECT -36.670 783.490 -35.490 784.670 ;
        RECT -36.670 605.090 -35.490 606.270 ;
        RECT -36.670 603.490 -35.490 604.670 ;
        RECT -36.670 425.090 -35.490 426.270 ;
        RECT -36.670 423.490 -35.490 424.670 ;
        RECT -36.670 245.090 -35.490 246.270 ;
        RECT -36.670 243.490 -35.490 244.670 ;
        RECT -36.670 65.090 -35.490 66.270 ;
        RECT -36.670 63.490 -35.490 64.670 ;
        RECT -36.670 -30.510 -35.490 -29.330 ;
        RECT -36.670 -32.110 -35.490 -30.930 ;
        RECT 58.930 3550.610 60.110 3551.790 ;
        RECT 58.930 3549.010 60.110 3550.190 ;
        RECT 58.930 3485.090 60.110 3486.270 ;
        RECT 58.930 3483.490 60.110 3484.670 ;
        RECT 58.930 3305.090 60.110 3306.270 ;
        RECT 58.930 3303.490 60.110 3304.670 ;
        RECT 58.930 3125.090 60.110 3126.270 ;
        RECT 58.930 3123.490 60.110 3124.670 ;
        RECT 58.930 2945.090 60.110 2946.270 ;
        RECT 58.930 2943.490 60.110 2944.670 ;
        RECT 58.930 2765.090 60.110 2766.270 ;
        RECT 58.930 2763.490 60.110 2764.670 ;
        RECT 58.930 2585.090 60.110 2586.270 ;
        RECT 58.930 2583.490 60.110 2584.670 ;
        RECT 58.930 2405.090 60.110 2406.270 ;
        RECT 58.930 2403.490 60.110 2404.670 ;
        RECT 58.930 2225.090 60.110 2226.270 ;
        RECT 58.930 2223.490 60.110 2224.670 ;
        RECT 58.930 2045.090 60.110 2046.270 ;
        RECT 58.930 2043.490 60.110 2044.670 ;
        RECT 58.930 1865.090 60.110 1866.270 ;
        RECT 58.930 1863.490 60.110 1864.670 ;
        RECT 58.930 1685.090 60.110 1686.270 ;
        RECT 58.930 1683.490 60.110 1684.670 ;
        RECT 58.930 1505.090 60.110 1506.270 ;
        RECT 58.930 1503.490 60.110 1504.670 ;
        RECT 58.930 1325.090 60.110 1326.270 ;
        RECT 58.930 1323.490 60.110 1324.670 ;
        RECT 58.930 1145.090 60.110 1146.270 ;
        RECT 58.930 1143.490 60.110 1144.670 ;
        RECT 58.930 965.090 60.110 966.270 ;
        RECT 58.930 963.490 60.110 964.670 ;
        RECT 58.930 785.090 60.110 786.270 ;
        RECT 58.930 783.490 60.110 784.670 ;
        RECT 58.930 605.090 60.110 606.270 ;
        RECT 58.930 603.490 60.110 604.670 ;
        RECT 58.930 425.090 60.110 426.270 ;
        RECT 58.930 423.490 60.110 424.670 ;
        RECT 58.930 245.090 60.110 246.270 ;
        RECT 58.930 243.490 60.110 244.670 ;
        RECT 58.930 65.090 60.110 66.270 ;
        RECT 58.930 63.490 60.110 64.670 ;
        RECT 58.930 -30.510 60.110 -29.330 ;
        RECT 58.930 -32.110 60.110 -30.930 ;
        RECT 238.930 3550.610 240.110 3551.790 ;
        RECT 238.930 3549.010 240.110 3550.190 ;
        RECT 238.930 3485.090 240.110 3486.270 ;
        RECT 238.930 3483.490 240.110 3484.670 ;
        RECT 238.930 3305.090 240.110 3306.270 ;
        RECT 238.930 3303.490 240.110 3304.670 ;
        RECT 238.930 3125.090 240.110 3126.270 ;
        RECT 238.930 3123.490 240.110 3124.670 ;
        RECT 238.930 2945.090 240.110 2946.270 ;
        RECT 238.930 2943.490 240.110 2944.670 ;
        RECT 238.930 2765.090 240.110 2766.270 ;
        RECT 238.930 2763.490 240.110 2764.670 ;
        RECT 238.930 2585.090 240.110 2586.270 ;
        RECT 238.930 2583.490 240.110 2584.670 ;
        RECT 238.930 2405.090 240.110 2406.270 ;
        RECT 238.930 2403.490 240.110 2404.670 ;
        RECT 238.930 2225.090 240.110 2226.270 ;
        RECT 238.930 2223.490 240.110 2224.670 ;
        RECT 238.930 2045.090 240.110 2046.270 ;
        RECT 238.930 2043.490 240.110 2044.670 ;
        RECT 238.930 1865.090 240.110 1866.270 ;
        RECT 238.930 1863.490 240.110 1864.670 ;
        RECT 238.930 1685.090 240.110 1686.270 ;
        RECT 238.930 1683.490 240.110 1684.670 ;
        RECT 238.930 1505.090 240.110 1506.270 ;
        RECT 238.930 1503.490 240.110 1504.670 ;
        RECT 238.930 1325.090 240.110 1326.270 ;
        RECT 238.930 1323.490 240.110 1324.670 ;
        RECT 238.930 1145.090 240.110 1146.270 ;
        RECT 238.930 1143.490 240.110 1144.670 ;
        RECT 238.930 965.090 240.110 966.270 ;
        RECT 238.930 963.490 240.110 964.670 ;
        RECT 238.930 785.090 240.110 786.270 ;
        RECT 238.930 783.490 240.110 784.670 ;
        RECT 238.930 605.090 240.110 606.270 ;
        RECT 238.930 603.490 240.110 604.670 ;
        RECT 238.930 425.090 240.110 426.270 ;
        RECT 238.930 423.490 240.110 424.670 ;
        RECT 238.930 245.090 240.110 246.270 ;
        RECT 238.930 243.490 240.110 244.670 ;
        RECT 238.930 65.090 240.110 66.270 ;
        RECT 238.930 63.490 240.110 64.670 ;
        RECT 238.930 -30.510 240.110 -29.330 ;
        RECT 238.930 -32.110 240.110 -30.930 ;
        RECT 418.930 3550.610 420.110 3551.790 ;
        RECT 418.930 3549.010 420.110 3550.190 ;
        RECT 418.930 3485.090 420.110 3486.270 ;
        RECT 418.930 3483.490 420.110 3484.670 ;
        RECT 418.930 3305.090 420.110 3306.270 ;
        RECT 418.930 3303.490 420.110 3304.670 ;
        RECT 418.930 3125.090 420.110 3126.270 ;
        RECT 418.930 3123.490 420.110 3124.670 ;
        RECT 418.930 2945.090 420.110 2946.270 ;
        RECT 418.930 2943.490 420.110 2944.670 ;
        RECT 418.930 2765.090 420.110 2766.270 ;
        RECT 418.930 2763.490 420.110 2764.670 ;
        RECT 418.930 2585.090 420.110 2586.270 ;
        RECT 418.930 2583.490 420.110 2584.670 ;
        RECT 418.930 2405.090 420.110 2406.270 ;
        RECT 418.930 2403.490 420.110 2404.670 ;
        RECT 418.930 2225.090 420.110 2226.270 ;
        RECT 418.930 2223.490 420.110 2224.670 ;
        RECT 418.930 2045.090 420.110 2046.270 ;
        RECT 418.930 2043.490 420.110 2044.670 ;
        RECT 418.930 1865.090 420.110 1866.270 ;
        RECT 418.930 1863.490 420.110 1864.670 ;
        RECT 418.930 1685.090 420.110 1686.270 ;
        RECT 418.930 1683.490 420.110 1684.670 ;
        RECT 418.930 1505.090 420.110 1506.270 ;
        RECT 418.930 1503.490 420.110 1504.670 ;
        RECT 418.930 1325.090 420.110 1326.270 ;
        RECT 418.930 1323.490 420.110 1324.670 ;
        RECT 418.930 1145.090 420.110 1146.270 ;
        RECT 418.930 1143.490 420.110 1144.670 ;
        RECT 418.930 965.090 420.110 966.270 ;
        RECT 418.930 963.490 420.110 964.670 ;
        RECT 418.930 785.090 420.110 786.270 ;
        RECT 418.930 783.490 420.110 784.670 ;
        RECT 418.930 605.090 420.110 606.270 ;
        RECT 418.930 603.490 420.110 604.670 ;
        RECT 418.930 425.090 420.110 426.270 ;
        RECT 418.930 423.490 420.110 424.670 ;
        RECT 418.930 245.090 420.110 246.270 ;
        RECT 418.930 243.490 420.110 244.670 ;
        RECT 418.930 65.090 420.110 66.270 ;
        RECT 418.930 63.490 420.110 64.670 ;
        RECT 418.930 -30.510 420.110 -29.330 ;
        RECT 418.930 -32.110 420.110 -30.930 ;
        RECT 598.930 3550.610 600.110 3551.790 ;
        RECT 598.930 3549.010 600.110 3550.190 ;
        RECT 598.930 3485.090 600.110 3486.270 ;
        RECT 598.930 3483.490 600.110 3484.670 ;
        RECT 598.930 3305.090 600.110 3306.270 ;
        RECT 598.930 3303.490 600.110 3304.670 ;
        RECT 598.930 3125.090 600.110 3126.270 ;
        RECT 598.930 3123.490 600.110 3124.670 ;
        RECT 598.930 2945.090 600.110 2946.270 ;
        RECT 598.930 2943.490 600.110 2944.670 ;
        RECT 598.930 2765.090 600.110 2766.270 ;
        RECT 598.930 2763.490 600.110 2764.670 ;
        RECT 598.930 2585.090 600.110 2586.270 ;
        RECT 598.930 2583.490 600.110 2584.670 ;
        RECT 598.930 2405.090 600.110 2406.270 ;
        RECT 598.930 2403.490 600.110 2404.670 ;
        RECT 598.930 2225.090 600.110 2226.270 ;
        RECT 598.930 2223.490 600.110 2224.670 ;
        RECT 598.930 2045.090 600.110 2046.270 ;
        RECT 598.930 2043.490 600.110 2044.670 ;
        RECT 598.930 1865.090 600.110 1866.270 ;
        RECT 598.930 1863.490 600.110 1864.670 ;
        RECT 598.930 1685.090 600.110 1686.270 ;
        RECT 598.930 1683.490 600.110 1684.670 ;
        RECT 598.930 1505.090 600.110 1506.270 ;
        RECT 598.930 1503.490 600.110 1504.670 ;
        RECT 598.930 1325.090 600.110 1326.270 ;
        RECT 598.930 1323.490 600.110 1324.670 ;
        RECT 598.930 1145.090 600.110 1146.270 ;
        RECT 598.930 1143.490 600.110 1144.670 ;
        RECT 598.930 965.090 600.110 966.270 ;
        RECT 598.930 963.490 600.110 964.670 ;
        RECT 598.930 785.090 600.110 786.270 ;
        RECT 598.930 783.490 600.110 784.670 ;
        RECT 598.930 605.090 600.110 606.270 ;
        RECT 598.930 603.490 600.110 604.670 ;
        RECT 598.930 425.090 600.110 426.270 ;
        RECT 598.930 423.490 600.110 424.670 ;
        RECT 598.930 245.090 600.110 246.270 ;
        RECT 598.930 243.490 600.110 244.670 ;
        RECT 598.930 65.090 600.110 66.270 ;
        RECT 598.930 63.490 600.110 64.670 ;
        RECT 598.930 -30.510 600.110 -29.330 ;
        RECT 598.930 -32.110 600.110 -30.930 ;
        RECT 778.930 3550.610 780.110 3551.790 ;
        RECT 778.930 3549.010 780.110 3550.190 ;
        RECT 778.930 3485.090 780.110 3486.270 ;
        RECT 778.930 3483.490 780.110 3484.670 ;
        RECT 778.930 3305.090 780.110 3306.270 ;
        RECT 778.930 3303.490 780.110 3304.670 ;
        RECT 778.930 3125.090 780.110 3126.270 ;
        RECT 778.930 3123.490 780.110 3124.670 ;
        RECT 778.930 2945.090 780.110 2946.270 ;
        RECT 778.930 2943.490 780.110 2944.670 ;
        RECT 778.930 2765.090 780.110 2766.270 ;
        RECT 778.930 2763.490 780.110 2764.670 ;
        RECT 778.930 2585.090 780.110 2586.270 ;
        RECT 778.930 2583.490 780.110 2584.670 ;
        RECT 778.930 2405.090 780.110 2406.270 ;
        RECT 778.930 2403.490 780.110 2404.670 ;
        RECT 778.930 2225.090 780.110 2226.270 ;
        RECT 778.930 2223.490 780.110 2224.670 ;
        RECT 778.930 2045.090 780.110 2046.270 ;
        RECT 778.930 2043.490 780.110 2044.670 ;
        RECT 778.930 1865.090 780.110 1866.270 ;
        RECT 778.930 1863.490 780.110 1864.670 ;
        RECT 778.930 1685.090 780.110 1686.270 ;
        RECT 778.930 1683.490 780.110 1684.670 ;
        RECT 778.930 1505.090 780.110 1506.270 ;
        RECT 778.930 1503.490 780.110 1504.670 ;
        RECT 778.930 1325.090 780.110 1326.270 ;
        RECT 778.930 1323.490 780.110 1324.670 ;
        RECT 778.930 1145.090 780.110 1146.270 ;
        RECT 778.930 1143.490 780.110 1144.670 ;
        RECT 778.930 965.090 780.110 966.270 ;
        RECT 778.930 963.490 780.110 964.670 ;
        RECT 778.930 785.090 780.110 786.270 ;
        RECT 778.930 783.490 780.110 784.670 ;
        RECT 778.930 605.090 780.110 606.270 ;
        RECT 778.930 603.490 780.110 604.670 ;
        RECT 778.930 425.090 780.110 426.270 ;
        RECT 778.930 423.490 780.110 424.670 ;
        RECT 778.930 245.090 780.110 246.270 ;
        RECT 778.930 243.490 780.110 244.670 ;
        RECT 778.930 65.090 780.110 66.270 ;
        RECT 778.930 63.490 780.110 64.670 ;
        RECT 778.930 -30.510 780.110 -29.330 ;
        RECT 778.930 -32.110 780.110 -30.930 ;
        RECT 958.930 3550.610 960.110 3551.790 ;
        RECT 958.930 3549.010 960.110 3550.190 ;
        RECT 958.930 3485.090 960.110 3486.270 ;
        RECT 958.930 3483.490 960.110 3484.670 ;
        RECT 958.930 3305.090 960.110 3306.270 ;
        RECT 958.930 3303.490 960.110 3304.670 ;
        RECT 958.930 3125.090 960.110 3126.270 ;
        RECT 958.930 3123.490 960.110 3124.670 ;
        RECT 958.930 2945.090 960.110 2946.270 ;
        RECT 958.930 2943.490 960.110 2944.670 ;
        RECT 958.930 2765.090 960.110 2766.270 ;
        RECT 958.930 2763.490 960.110 2764.670 ;
        RECT 958.930 2585.090 960.110 2586.270 ;
        RECT 958.930 2583.490 960.110 2584.670 ;
        RECT 958.930 2405.090 960.110 2406.270 ;
        RECT 958.930 2403.490 960.110 2404.670 ;
        RECT 958.930 2225.090 960.110 2226.270 ;
        RECT 958.930 2223.490 960.110 2224.670 ;
        RECT 958.930 2045.090 960.110 2046.270 ;
        RECT 958.930 2043.490 960.110 2044.670 ;
        RECT 958.930 1865.090 960.110 1866.270 ;
        RECT 958.930 1863.490 960.110 1864.670 ;
        RECT 958.930 1685.090 960.110 1686.270 ;
        RECT 958.930 1683.490 960.110 1684.670 ;
        RECT 958.930 1505.090 960.110 1506.270 ;
        RECT 958.930 1503.490 960.110 1504.670 ;
        RECT 958.930 1325.090 960.110 1326.270 ;
        RECT 958.930 1323.490 960.110 1324.670 ;
        RECT 958.930 1145.090 960.110 1146.270 ;
        RECT 958.930 1143.490 960.110 1144.670 ;
        RECT 958.930 965.090 960.110 966.270 ;
        RECT 958.930 963.490 960.110 964.670 ;
        RECT 958.930 785.090 960.110 786.270 ;
        RECT 958.930 783.490 960.110 784.670 ;
        RECT 958.930 605.090 960.110 606.270 ;
        RECT 958.930 603.490 960.110 604.670 ;
        RECT 958.930 425.090 960.110 426.270 ;
        RECT 958.930 423.490 960.110 424.670 ;
        RECT 958.930 245.090 960.110 246.270 ;
        RECT 958.930 243.490 960.110 244.670 ;
        RECT 958.930 65.090 960.110 66.270 ;
        RECT 958.930 63.490 960.110 64.670 ;
        RECT 958.930 -30.510 960.110 -29.330 ;
        RECT 958.930 -32.110 960.110 -30.930 ;
        RECT 1138.930 3550.610 1140.110 3551.790 ;
        RECT 1138.930 3549.010 1140.110 3550.190 ;
        RECT 1138.930 3485.090 1140.110 3486.270 ;
        RECT 1138.930 3483.490 1140.110 3484.670 ;
        RECT 1138.930 3305.090 1140.110 3306.270 ;
        RECT 1138.930 3303.490 1140.110 3304.670 ;
        RECT 1138.930 3125.090 1140.110 3126.270 ;
        RECT 1138.930 3123.490 1140.110 3124.670 ;
        RECT 1138.930 2945.090 1140.110 2946.270 ;
        RECT 1138.930 2943.490 1140.110 2944.670 ;
        RECT 1138.930 2765.090 1140.110 2766.270 ;
        RECT 1138.930 2763.490 1140.110 2764.670 ;
        RECT 1138.930 2585.090 1140.110 2586.270 ;
        RECT 1138.930 2583.490 1140.110 2584.670 ;
        RECT 1138.930 2405.090 1140.110 2406.270 ;
        RECT 1138.930 2403.490 1140.110 2404.670 ;
        RECT 1138.930 2225.090 1140.110 2226.270 ;
        RECT 1138.930 2223.490 1140.110 2224.670 ;
        RECT 1138.930 2045.090 1140.110 2046.270 ;
        RECT 1138.930 2043.490 1140.110 2044.670 ;
        RECT 1138.930 1865.090 1140.110 1866.270 ;
        RECT 1138.930 1863.490 1140.110 1864.670 ;
        RECT 1138.930 1685.090 1140.110 1686.270 ;
        RECT 1138.930 1683.490 1140.110 1684.670 ;
        RECT 1138.930 1505.090 1140.110 1506.270 ;
        RECT 1138.930 1503.490 1140.110 1504.670 ;
        RECT 1138.930 1325.090 1140.110 1326.270 ;
        RECT 1138.930 1323.490 1140.110 1324.670 ;
        RECT 1138.930 1145.090 1140.110 1146.270 ;
        RECT 1138.930 1143.490 1140.110 1144.670 ;
        RECT 1138.930 965.090 1140.110 966.270 ;
        RECT 1138.930 963.490 1140.110 964.670 ;
        RECT 1138.930 785.090 1140.110 786.270 ;
        RECT 1138.930 783.490 1140.110 784.670 ;
        RECT 1138.930 605.090 1140.110 606.270 ;
        RECT 1138.930 603.490 1140.110 604.670 ;
        RECT 1138.930 425.090 1140.110 426.270 ;
        RECT 1138.930 423.490 1140.110 424.670 ;
        RECT 1138.930 245.090 1140.110 246.270 ;
        RECT 1138.930 243.490 1140.110 244.670 ;
        RECT 1138.930 65.090 1140.110 66.270 ;
        RECT 1138.930 63.490 1140.110 64.670 ;
        RECT 1138.930 -30.510 1140.110 -29.330 ;
        RECT 1138.930 -32.110 1140.110 -30.930 ;
        RECT 1318.930 3550.610 1320.110 3551.790 ;
        RECT 1318.930 3549.010 1320.110 3550.190 ;
        RECT 1318.930 3485.090 1320.110 3486.270 ;
        RECT 1318.930 3483.490 1320.110 3484.670 ;
        RECT 1318.930 3305.090 1320.110 3306.270 ;
        RECT 1318.930 3303.490 1320.110 3304.670 ;
        RECT 1318.930 3125.090 1320.110 3126.270 ;
        RECT 1318.930 3123.490 1320.110 3124.670 ;
        RECT 1318.930 2945.090 1320.110 2946.270 ;
        RECT 1318.930 2943.490 1320.110 2944.670 ;
        RECT 1318.930 2765.090 1320.110 2766.270 ;
        RECT 1318.930 2763.490 1320.110 2764.670 ;
        RECT 1318.930 2585.090 1320.110 2586.270 ;
        RECT 1318.930 2583.490 1320.110 2584.670 ;
        RECT 1318.930 2405.090 1320.110 2406.270 ;
        RECT 1318.930 2403.490 1320.110 2404.670 ;
        RECT 1318.930 2225.090 1320.110 2226.270 ;
        RECT 1318.930 2223.490 1320.110 2224.670 ;
        RECT 1318.930 2045.090 1320.110 2046.270 ;
        RECT 1318.930 2043.490 1320.110 2044.670 ;
        RECT 1318.930 1865.090 1320.110 1866.270 ;
        RECT 1318.930 1863.490 1320.110 1864.670 ;
        RECT 1318.930 1685.090 1320.110 1686.270 ;
        RECT 1318.930 1683.490 1320.110 1684.670 ;
        RECT 1318.930 1505.090 1320.110 1506.270 ;
        RECT 1318.930 1503.490 1320.110 1504.670 ;
        RECT 1318.930 1325.090 1320.110 1326.270 ;
        RECT 1318.930 1323.490 1320.110 1324.670 ;
        RECT 1318.930 1145.090 1320.110 1146.270 ;
        RECT 1318.930 1143.490 1320.110 1144.670 ;
        RECT 1318.930 965.090 1320.110 966.270 ;
        RECT 1318.930 963.490 1320.110 964.670 ;
        RECT 1318.930 785.090 1320.110 786.270 ;
        RECT 1318.930 783.490 1320.110 784.670 ;
        RECT 1318.930 605.090 1320.110 606.270 ;
        RECT 1318.930 603.490 1320.110 604.670 ;
        RECT 1318.930 425.090 1320.110 426.270 ;
        RECT 1318.930 423.490 1320.110 424.670 ;
        RECT 1318.930 245.090 1320.110 246.270 ;
        RECT 1318.930 243.490 1320.110 244.670 ;
        RECT 1318.930 65.090 1320.110 66.270 ;
        RECT 1318.930 63.490 1320.110 64.670 ;
        RECT 1318.930 -30.510 1320.110 -29.330 ;
        RECT 1318.930 -32.110 1320.110 -30.930 ;
        RECT 1498.930 3550.610 1500.110 3551.790 ;
        RECT 1498.930 3549.010 1500.110 3550.190 ;
        RECT 1498.930 3485.090 1500.110 3486.270 ;
        RECT 1498.930 3483.490 1500.110 3484.670 ;
        RECT 1498.930 3305.090 1500.110 3306.270 ;
        RECT 1498.930 3303.490 1500.110 3304.670 ;
        RECT 1498.930 3125.090 1500.110 3126.270 ;
        RECT 1498.930 3123.490 1500.110 3124.670 ;
        RECT 1498.930 2945.090 1500.110 2946.270 ;
        RECT 1498.930 2943.490 1500.110 2944.670 ;
        RECT 1498.930 2765.090 1500.110 2766.270 ;
        RECT 1498.930 2763.490 1500.110 2764.670 ;
        RECT 1498.930 2585.090 1500.110 2586.270 ;
        RECT 1498.930 2583.490 1500.110 2584.670 ;
        RECT 1498.930 2405.090 1500.110 2406.270 ;
        RECT 1498.930 2403.490 1500.110 2404.670 ;
        RECT 1498.930 2225.090 1500.110 2226.270 ;
        RECT 1498.930 2223.490 1500.110 2224.670 ;
        RECT 1498.930 2045.090 1500.110 2046.270 ;
        RECT 1498.930 2043.490 1500.110 2044.670 ;
        RECT 1498.930 1865.090 1500.110 1866.270 ;
        RECT 1498.930 1863.490 1500.110 1864.670 ;
        RECT 1498.930 1685.090 1500.110 1686.270 ;
        RECT 1498.930 1683.490 1500.110 1684.670 ;
        RECT 1498.930 1505.090 1500.110 1506.270 ;
        RECT 1498.930 1503.490 1500.110 1504.670 ;
        RECT 1498.930 1325.090 1500.110 1326.270 ;
        RECT 1498.930 1323.490 1500.110 1324.670 ;
        RECT 1498.930 1145.090 1500.110 1146.270 ;
        RECT 1498.930 1143.490 1500.110 1144.670 ;
        RECT 1498.930 965.090 1500.110 966.270 ;
        RECT 1498.930 963.490 1500.110 964.670 ;
        RECT 1498.930 785.090 1500.110 786.270 ;
        RECT 1498.930 783.490 1500.110 784.670 ;
        RECT 1498.930 605.090 1500.110 606.270 ;
        RECT 1498.930 603.490 1500.110 604.670 ;
        RECT 1498.930 425.090 1500.110 426.270 ;
        RECT 1498.930 423.490 1500.110 424.670 ;
        RECT 1498.930 245.090 1500.110 246.270 ;
        RECT 1498.930 243.490 1500.110 244.670 ;
        RECT 1498.930 65.090 1500.110 66.270 ;
        RECT 1498.930 63.490 1500.110 64.670 ;
        RECT 1498.930 -30.510 1500.110 -29.330 ;
        RECT 1498.930 -32.110 1500.110 -30.930 ;
        RECT 1678.930 3550.610 1680.110 3551.790 ;
        RECT 1678.930 3549.010 1680.110 3550.190 ;
        RECT 1678.930 3485.090 1680.110 3486.270 ;
        RECT 1678.930 3483.490 1680.110 3484.670 ;
        RECT 1678.930 3305.090 1680.110 3306.270 ;
        RECT 1678.930 3303.490 1680.110 3304.670 ;
        RECT 1678.930 3125.090 1680.110 3126.270 ;
        RECT 1678.930 3123.490 1680.110 3124.670 ;
        RECT 1678.930 2945.090 1680.110 2946.270 ;
        RECT 1678.930 2943.490 1680.110 2944.670 ;
        RECT 1678.930 2765.090 1680.110 2766.270 ;
        RECT 1678.930 2763.490 1680.110 2764.670 ;
        RECT 1678.930 2585.090 1680.110 2586.270 ;
        RECT 1678.930 2583.490 1680.110 2584.670 ;
        RECT 1678.930 2405.090 1680.110 2406.270 ;
        RECT 1678.930 2403.490 1680.110 2404.670 ;
        RECT 1678.930 2225.090 1680.110 2226.270 ;
        RECT 1678.930 2223.490 1680.110 2224.670 ;
        RECT 1678.930 2045.090 1680.110 2046.270 ;
        RECT 1678.930 2043.490 1680.110 2044.670 ;
        RECT 1678.930 1865.090 1680.110 1866.270 ;
        RECT 1678.930 1863.490 1680.110 1864.670 ;
        RECT 1678.930 1685.090 1680.110 1686.270 ;
        RECT 1678.930 1683.490 1680.110 1684.670 ;
        RECT 1678.930 1505.090 1680.110 1506.270 ;
        RECT 1678.930 1503.490 1680.110 1504.670 ;
        RECT 1678.930 1325.090 1680.110 1326.270 ;
        RECT 1678.930 1323.490 1680.110 1324.670 ;
        RECT 1678.930 1145.090 1680.110 1146.270 ;
        RECT 1678.930 1143.490 1680.110 1144.670 ;
        RECT 1678.930 965.090 1680.110 966.270 ;
        RECT 1678.930 963.490 1680.110 964.670 ;
        RECT 1678.930 785.090 1680.110 786.270 ;
        RECT 1678.930 783.490 1680.110 784.670 ;
        RECT 1678.930 605.090 1680.110 606.270 ;
        RECT 1678.930 603.490 1680.110 604.670 ;
        RECT 1678.930 425.090 1680.110 426.270 ;
        RECT 1678.930 423.490 1680.110 424.670 ;
        RECT 1678.930 245.090 1680.110 246.270 ;
        RECT 1678.930 243.490 1680.110 244.670 ;
        RECT 1678.930 65.090 1680.110 66.270 ;
        RECT 1678.930 63.490 1680.110 64.670 ;
        RECT 1678.930 -30.510 1680.110 -29.330 ;
        RECT 1678.930 -32.110 1680.110 -30.930 ;
        RECT 1858.930 3550.610 1860.110 3551.790 ;
        RECT 1858.930 3549.010 1860.110 3550.190 ;
        RECT 1858.930 3485.090 1860.110 3486.270 ;
        RECT 1858.930 3483.490 1860.110 3484.670 ;
        RECT 1858.930 3305.090 1860.110 3306.270 ;
        RECT 1858.930 3303.490 1860.110 3304.670 ;
        RECT 1858.930 3125.090 1860.110 3126.270 ;
        RECT 1858.930 3123.490 1860.110 3124.670 ;
        RECT 1858.930 2945.090 1860.110 2946.270 ;
        RECT 1858.930 2943.490 1860.110 2944.670 ;
        RECT 1858.930 2765.090 1860.110 2766.270 ;
        RECT 1858.930 2763.490 1860.110 2764.670 ;
        RECT 1858.930 2585.090 1860.110 2586.270 ;
        RECT 1858.930 2583.490 1860.110 2584.670 ;
        RECT 1858.930 2405.090 1860.110 2406.270 ;
        RECT 1858.930 2403.490 1860.110 2404.670 ;
        RECT 1858.930 2225.090 1860.110 2226.270 ;
        RECT 1858.930 2223.490 1860.110 2224.670 ;
        RECT 1858.930 2045.090 1860.110 2046.270 ;
        RECT 1858.930 2043.490 1860.110 2044.670 ;
        RECT 1858.930 1865.090 1860.110 1866.270 ;
        RECT 1858.930 1863.490 1860.110 1864.670 ;
        RECT 1858.930 1685.090 1860.110 1686.270 ;
        RECT 1858.930 1683.490 1860.110 1684.670 ;
        RECT 1858.930 1505.090 1860.110 1506.270 ;
        RECT 1858.930 1503.490 1860.110 1504.670 ;
        RECT 1858.930 1325.090 1860.110 1326.270 ;
        RECT 1858.930 1323.490 1860.110 1324.670 ;
        RECT 1858.930 1145.090 1860.110 1146.270 ;
        RECT 1858.930 1143.490 1860.110 1144.670 ;
        RECT 1858.930 965.090 1860.110 966.270 ;
        RECT 1858.930 963.490 1860.110 964.670 ;
        RECT 1858.930 785.090 1860.110 786.270 ;
        RECT 1858.930 783.490 1860.110 784.670 ;
        RECT 1858.930 605.090 1860.110 606.270 ;
        RECT 1858.930 603.490 1860.110 604.670 ;
        RECT 1858.930 425.090 1860.110 426.270 ;
        RECT 1858.930 423.490 1860.110 424.670 ;
        RECT 1858.930 245.090 1860.110 246.270 ;
        RECT 1858.930 243.490 1860.110 244.670 ;
        RECT 1858.930 65.090 1860.110 66.270 ;
        RECT 1858.930 63.490 1860.110 64.670 ;
        RECT 1858.930 -30.510 1860.110 -29.330 ;
        RECT 1858.930 -32.110 1860.110 -30.930 ;
        RECT 2038.930 3550.610 2040.110 3551.790 ;
        RECT 2038.930 3549.010 2040.110 3550.190 ;
        RECT 2038.930 3485.090 2040.110 3486.270 ;
        RECT 2038.930 3483.490 2040.110 3484.670 ;
        RECT 2038.930 3305.090 2040.110 3306.270 ;
        RECT 2038.930 3303.490 2040.110 3304.670 ;
        RECT 2038.930 3125.090 2040.110 3126.270 ;
        RECT 2038.930 3123.490 2040.110 3124.670 ;
        RECT 2038.930 2945.090 2040.110 2946.270 ;
        RECT 2038.930 2943.490 2040.110 2944.670 ;
        RECT 2038.930 2765.090 2040.110 2766.270 ;
        RECT 2038.930 2763.490 2040.110 2764.670 ;
        RECT 2038.930 2585.090 2040.110 2586.270 ;
        RECT 2038.930 2583.490 2040.110 2584.670 ;
        RECT 2038.930 2405.090 2040.110 2406.270 ;
        RECT 2038.930 2403.490 2040.110 2404.670 ;
        RECT 2038.930 2225.090 2040.110 2226.270 ;
        RECT 2038.930 2223.490 2040.110 2224.670 ;
        RECT 2038.930 2045.090 2040.110 2046.270 ;
        RECT 2038.930 2043.490 2040.110 2044.670 ;
        RECT 2038.930 1865.090 2040.110 1866.270 ;
        RECT 2038.930 1863.490 2040.110 1864.670 ;
        RECT 2038.930 1685.090 2040.110 1686.270 ;
        RECT 2038.930 1683.490 2040.110 1684.670 ;
        RECT 2038.930 1505.090 2040.110 1506.270 ;
        RECT 2038.930 1503.490 2040.110 1504.670 ;
        RECT 2038.930 1325.090 2040.110 1326.270 ;
        RECT 2038.930 1323.490 2040.110 1324.670 ;
        RECT 2038.930 1145.090 2040.110 1146.270 ;
        RECT 2038.930 1143.490 2040.110 1144.670 ;
        RECT 2038.930 965.090 2040.110 966.270 ;
        RECT 2038.930 963.490 2040.110 964.670 ;
        RECT 2038.930 785.090 2040.110 786.270 ;
        RECT 2038.930 783.490 2040.110 784.670 ;
        RECT 2038.930 605.090 2040.110 606.270 ;
        RECT 2038.930 603.490 2040.110 604.670 ;
        RECT 2038.930 425.090 2040.110 426.270 ;
        RECT 2038.930 423.490 2040.110 424.670 ;
        RECT 2038.930 245.090 2040.110 246.270 ;
        RECT 2038.930 243.490 2040.110 244.670 ;
        RECT 2038.930 65.090 2040.110 66.270 ;
        RECT 2038.930 63.490 2040.110 64.670 ;
        RECT 2038.930 -30.510 2040.110 -29.330 ;
        RECT 2038.930 -32.110 2040.110 -30.930 ;
        RECT 2218.930 3550.610 2220.110 3551.790 ;
        RECT 2218.930 3549.010 2220.110 3550.190 ;
        RECT 2218.930 3485.090 2220.110 3486.270 ;
        RECT 2218.930 3483.490 2220.110 3484.670 ;
        RECT 2218.930 3305.090 2220.110 3306.270 ;
        RECT 2218.930 3303.490 2220.110 3304.670 ;
        RECT 2218.930 3125.090 2220.110 3126.270 ;
        RECT 2218.930 3123.490 2220.110 3124.670 ;
        RECT 2218.930 2945.090 2220.110 2946.270 ;
        RECT 2218.930 2943.490 2220.110 2944.670 ;
        RECT 2218.930 2765.090 2220.110 2766.270 ;
        RECT 2218.930 2763.490 2220.110 2764.670 ;
        RECT 2218.930 2585.090 2220.110 2586.270 ;
        RECT 2218.930 2583.490 2220.110 2584.670 ;
        RECT 2218.930 2405.090 2220.110 2406.270 ;
        RECT 2218.930 2403.490 2220.110 2404.670 ;
        RECT 2218.930 2225.090 2220.110 2226.270 ;
        RECT 2218.930 2223.490 2220.110 2224.670 ;
        RECT 2218.930 2045.090 2220.110 2046.270 ;
        RECT 2218.930 2043.490 2220.110 2044.670 ;
        RECT 2218.930 1865.090 2220.110 1866.270 ;
        RECT 2218.930 1863.490 2220.110 1864.670 ;
        RECT 2218.930 1685.090 2220.110 1686.270 ;
        RECT 2218.930 1683.490 2220.110 1684.670 ;
        RECT 2218.930 1505.090 2220.110 1506.270 ;
        RECT 2218.930 1503.490 2220.110 1504.670 ;
        RECT 2218.930 1325.090 2220.110 1326.270 ;
        RECT 2218.930 1323.490 2220.110 1324.670 ;
        RECT 2218.930 1145.090 2220.110 1146.270 ;
        RECT 2218.930 1143.490 2220.110 1144.670 ;
        RECT 2218.930 965.090 2220.110 966.270 ;
        RECT 2218.930 963.490 2220.110 964.670 ;
        RECT 2218.930 785.090 2220.110 786.270 ;
        RECT 2218.930 783.490 2220.110 784.670 ;
        RECT 2218.930 605.090 2220.110 606.270 ;
        RECT 2218.930 603.490 2220.110 604.670 ;
        RECT 2218.930 425.090 2220.110 426.270 ;
        RECT 2218.930 423.490 2220.110 424.670 ;
        RECT 2218.930 245.090 2220.110 246.270 ;
        RECT 2218.930 243.490 2220.110 244.670 ;
        RECT 2218.930 65.090 2220.110 66.270 ;
        RECT 2218.930 63.490 2220.110 64.670 ;
        RECT 2218.930 -30.510 2220.110 -29.330 ;
        RECT 2218.930 -32.110 2220.110 -30.930 ;
        RECT 2398.930 3550.610 2400.110 3551.790 ;
        RECT 2398.930 3549.010 2400.110 3550.190 ;
        RECT 2398.930 3485.090 2400.110 3486.270 ;
        RECT 2398.930 3483.490 2400.110 3484.670 ;
        RECT 2398.930 3305.090 2400.110 3306.270 ;
        RECT 2398.930 3303.490 2400.110 3304.670 ;
        RECT 2398.930 3125.090 2400.110 3126.270 ;
        RECT 2398.930 3123.490 2400.110 3124.670 ;
        RECT 2398.930 2945.090 2400.110 2946.270 ;
        RECT 2398.930 2943.490 2400.110 2944.670 ;
        RECT 2398.930 2765.090 2400.110 2766.270 ;
        RECT 2398.930 2763.490 2400.110 2764.670 ;
        RECT 2398.930 2585.090 2400.110 2586.270 ;
        RECT 2398.930 2583.490 2400.110 2584.670 ;
        RECT 2398.930 2405.090 2400.110 2406.270 ;
        RECT 2398.930 2403.490 2400.110 2404.670 ;
        RECT 2398.930 2225.090 2400.110 2226.270 ;
        RECT 2398.930 2223.490 2400.110 2224.670 ;
        RECT 2398.930 2045.090 2400.110 2046.270 ;
        RECT 2398.930 2043.490 2400.110 2044.670 ;
        RECT 2398.930 1865.090 2400.110 1866.270 ;
        RECT 2398.930 1863.490 2400.110 1864.670 ;
        RECT 2398.930 1685.090 2400.110 1686.270 ;
        RECT 2398.930 1683.490 2400.110 1684.670 ;
        RECT 2398.930 1505.090 2400.110 1506.270 ;
        RECT 2398.930 1503.490 2400.110 1504.670 ;
        RECT 2398.930 1325.090 2400.110 1326.270 ;
        RECT 2398.930 1323.490 2400.110 1324.670 ;
        RECT 2398.930 1145.090 2400.110 1146.270 ;
        RECT 2398.930 1143.490 2400.110 1144.670 ;
        RECT 2398.930 965.090 2400.110 966.270 ;
        RECT 2398.930 963.490 2400.110 964.670 ;
        RECT 2398.930 785.090 2400.110 786.270 ;
        RECT 2398.930 783.490 2400.110 784.670 ;
        RECT 2398.930 605.090 2400.110 606.270 ;
        RECT 2398.930 603.490 2400.110 604.670 ;
        RECT 2398.930 425.090 2400.110 426.270 ;
        RECT 2398.930 423.490 2400.110 424.670 ;
        RECT 2398.930 245.090 2400.110 246.270 ;
        RECT 2398.930 243.490 2400.110 244.670 ;
        RECT 2398.930 65.090 2400.110 66.270 ;
        RECT 2398.930 63.490 2400.110 64.670 ;
        RECT 2398.930 -30.510 2400.110 -29.330 ;
        RECT 2398.930 -32.110 2400.110 -30.930 ;
        RECT 2578.930 3550.610 2580.110 3551.790 ;
        RECT 2578.930 3549.010 2580.110 3550.190 ;
        RECT 2578.930 3485.090 2580.110 3486.270 ;
        RECT 2578.930 3483.490 2580.110 3484.670 ;
        RECT 2578.930 3305.090 2580.110 3306.270 ;
        RECT 2578.930 3303.490 2580.110 3304.670 ;
        RECT 2578.930 3125.090 2580.110 3126.270 ;
        RECT 2578.930 3123.490 2580.110 3124.670 ;
        RECT 2578.930 2945.090 2580.110 2946.270 ;
        RECT 2578.930 2943.490 2580.110 2944.670 ;
        RECT 2578.930 2765.090 2580.110 2766.270 ;
        RECT 2578.930 2763.490 2580.110 2764.670 ;
        RECT 2578.930 2585.090 2580.110 2586.270 ;
        RECT 2578.930 2583.490 2580.110 2584.670 ;
        RECT 2578.930 2405.090 2580.110 2406.270 ;
        RECT 2578.930 2403.490 2580.110 2404.670 ;
        RECT 2578.930 2225.090 2580.110 2226.270 ;
        RECT 2578.930 2223.490 2580.110 2224.670 ;
        RECT 2578.930 2045.090 2580.110 2046.270 ;
        RECT 2578.930 2043.490 2580.110 2044.670 ;
        RECT 2578.930 1865.090 2580.110 1866.270 ;
        RECT 2578.930 1863.490 2580.110 1864.670 ;
        RECT 2578.930 1685.090 2580.110 1686.270 ;
        RECT 2578.930 1683.490 2580.110 1684.670 ;
        RECT 2578.930 1505.090 2580.110 1506.270 ;
        RECT 2578.930 1503.490 2580.110 1504.670 ;
        RECT 2578.930 1325.090 2580.110 1326.270 ;
        RECT 2578.930 1323.490 2580.110 1324.670 ;
        RECT 2578.930 1145.090 2580.110 1146.270 ;
        RECT 2578.930 1143.490 2580.110 1144.670 ;
        RECT 2578.930 965.090 2580.110 966.270 ;
        RECT 2578.930 963.490 2580.110 964.670 ;
        RECT 2578.930 785.090 2580.110 786.270 ;
        RECT 2578.930 783.490 2580.110 784.670 ;
        RECT 2578.930 605.090 2580.110 606.270 ;
        RECT 2578.930 603.490 2580.110 604.670 ;
        RECT 2578.930 425.090 2580.110 426.270 ;
        RECT 2578.930 423.490 2580.110 424.670 ;
        RECT 2578.930 245.090 2580.110 246.270 ;
        RECT 2578.930 243.490 2580.110 244.670 ;
        RECT 2578.930 65.090 2580.110 66.270 ;
        RECT 2578.930 63.490 2580.110 64.670 ;
        RECT 2578.930 -30.510 2580.110 -29.330 ;
        RECT 2578.930 -32.110 2580.110 -30.930 ;
        RECT 2758.930 3550.610 2760.110 3551.790 ;
        RECT 2758.930 3549.010 2760.110 3550.190 ;
        RECT 2758.930 3485.090 2760.110 3486.270 ;
        RECT 2758.930 3483.490 2760.110 3484.670 ;
        RECT 2758.930 3305.090 2760.110 3306.270 ;
        RECT 2758.930 3303.490 2760.110 3304.670 ;
        RECT 2758.930 3125.090 2760.110 3126.270 ;
        RECT 2758.930 3123.490 2760.110 3124.670 ;
        RECT 2758.930 2945.090 2760.110 2946.270 ;
        RECT 2758.930 2943.490 2760.110 2944.670 ;
        RECT 2758.930 2765.090 2760.110 2766.270 ;
        RECT 2758.930 2763.490 2760.110 2764.670 ;
        RECT 2758.930 2585.090 2760.110 2586.270 ;
        RECT 2758.930 2583.490 2760.110 2584.670 ;
        RECT 2758.930 2405.090 2760.110 2406.270 ;
        RECT 2758.930 2403.490 2760.110 2404.670 ;
        RECT 2758.930 2225.090 2760.110 2226.270 ;
        RECT 2758.930 2223.490 2760.110 2224.670 ;
        RECT 2758.930 2045.090 2760.110 2046.270 ;
        RECT 2758.930 2043.490 2760.110 2044.670 ;
        RECT 2758.930 1865.090 2760.110 1866.270 ;
        RECT 2758.930 1863.490 2760.110 1864.670 ;
        RECT 2758.930 1685.090 2760.110 1686.270 ;
        RECT 2758.930 1683.490 2760.110 1684.670 ;
        RECT 2758.930 1505.090 2760.110 1506.270 ;
        RECT 2758.930 1503.490 2760.110 1504.670 ;
        RECT 2758.930 1325.090 2760.110 1326.270 ;
        RECT 2758.930 1323.490 2760.110 1324.670 ;
        RECT 2758.930 1145.090 2760.110 1146.270 ;
        RECT 2758.930 1143.490 2760.110 1144.670 ;
        RECT 2758.930 965.090 2760.110 966.270 ;
        RECT 2758.930 963.490 2760.110 964.670 ;
        RECT 2758.930 785.090 2760.110 786.270 ;
        RECT 2758.930 783.490 2760.110 784.670 ;
        RECT 2758.930 605.090 2760.110 606.270 ;
        RECT 2758.930 603.490 2760.110 604.670 ;
        RECT 2758.930 425.090 2760.110 426.270 ;
        RECT 2758.930 423.490 2760.110 424.670 ;
        RECT 2758.930 245.090 2760.110 246.270 ;
        RECT 2758.930 243.490 2760.110 244.670 ;
        RECT 2758.930 65.090 2760.110 66.270 ;
        RECT 2758.930 63.490 2760.110 64.670 ;
        RECT 2758.930 -30.510 2760.110 -29.330 ;
        RECT 2758.930 -32.110 2760.110 -30.930 ;
        RECT 2955.110 3550.610 2956.290 3551.790 ;
        RECT 2955.110 3549.010 2956.290 3550.190 ;
        RECT 2955.110 3485.090 2956.290 3486.270 ;
        RECT 2955.110 3483.490 2956.290 3484.670 ;
        RECT 2955.110 3305.090 2956.290 3306.270 ;
        RECT 2955.110 3303.490 2956.290 3304.670 ;
        RECT 2955.110 3125.090 2956.290 3126.270 ;
        RECT 2955.110 3123.490 2956.290 3124.670 ;
        RECT 2955.110 2945.090 2956.290 2946.270 ;
        RECT 2955.110 2943.490 2956.290 2944.670 ;
        RECT 2955.110 2765.090 2956.290 2766.270 ;
        RECT 2955.110 2763.490 2956.290 2764.670 ;
        RECT 2955.110 2585.090 2956.290 2586.270 ;
        RECT 2955.110 2583.490 2956.290 2584.670 ;
        RECT 2955.110 2405.090 2956.290 2406.270 ;
        RECT 2955.110 2403.490 2956.290 2404.670 ;
        RECT 2955.110 2225.090 2956.290 2226.270 ;
        RECT 2955.110 2223.490 2956.290 2224.670 ;
        RECT 2955.110 2045.090 2956.290 2046.270 ;
        RECT 2955.110 2043.490 2956.290 2044.670 ;
        RECT 2955.110 1865.090 2956.290 1866.270 ;
        RECT 2955.110 1863.490 2956.290 1864.670 ;
        RECT 2955.110 1685.090 2956.290 1686.270 ;
        RECT 2955.110 1683.490 2956.290 1684.670 ;
        RECT 2955.110 1505.090 2956.290 1506.270 ;
        RECT 2955.110 1503.490 2956.290 1504.670 ;
        RECT 2955.110 1325.090 2956.290 1326.270 ;
        RECT 2955.110 1323.490 2956.290 1324.670 ;
        RECT 2955.110 1145.090 2956.290 1146.270 ;
        RECT 2955.110 1143.490 2956.290 1144.670 ;
        RECT 2955.110 965.090 2956.290 966.270 ;
        RECT 2955.110 963.490 2956.290 964.670 ;
        RECT 2955.110 785.090 2956.290 786.270 ;
        RECT 2955.110 783.490 2956.290 784.670 ;
        RECT 2955.110 605.090 2956.290 606.270 ;
        RECT 2955.110 603.490 2956.290 604.670 ;
        RECT 2955.110 425.090 2956.290 426.270 ;
        RECT 2955.110 423.490 2956.290 424.670 ;
        RECT 2955.110 245.090 2956.290 246.270 ;
        RECT 2955.110 243.490 2956.290 244.670 ;
        RECT 2955.110 65.090 2956.290 66.270 ;
        RECT 2955.110 63.490 2956.290 64.670 ;
        RECT 2955.110 -30.510 2956.290 -29.330 ;
        RECT 2955.110 -32.110 2956.290 -30.930 ;
      LAYER met5 ;
        RECT -37.580 3551.900 -34.580 3551.910 ;
        RECT 58.020 3551.900 61.020 3551.910 ;
        RECT 238.020 3551.900 241.020 3551.910 ;
        RECT 418.020 3551.900 421.020 3551.910 ;
        RECT 598.020 3551.900 601.020 3551.910 ;
        RECT 778.020 3551.900 781.020 3551.910 ;
        RECT 958.020 3551.900 961.020 3551.910 ;
        RECT 1138.020 3551.900 1141.020 3551.910 ;
        RECT 1318.020 3551.900 1321.020 3551.910 ;
        RECT 1498.020 3551.900 1501.020 3551.910 ;
        RECT 1678.020 3551.900 1681.020 3551.910 ;
        RECT 1858.020 3551.900 1861.020 3551.910 ;
        RECT 2038.020 3551.900 2041.020 3551.910 ;
        RECT 2218.020 3551.900 2221.020 3551.910 ;
        RECT 2398.020 3551.900 2401.020 3551.910 ;
        RECT 2578.020 3551.900 2581.020 3551.910 ;
        RECT 2758.020 3551.900 2761.020 3551.910 ;
        RECT 2954.200 3551.900 2957.200 3551.910 ;
        RECT -37.580 3548.900 2957.200 3551.900 ;
        RECT -37.580 3548.890 -34.580 3548.900 ;
        RECT 58.020 3548.890 61.020 3548.900 ;
        RECT 238.020 3548.890 241.020 3548.900 ;
        RECT 418.020 3548.890 421.020 3548.900 ;
        RECT 598.020 3548.890 601.020 3548.900 ;
        RECT 778.020 3548.890 781.020 3548.900 ;
        RECT 958.020 3548.890 961.020 3548.900 ;
        RECT 1138.020 3548.890 1141.020 3548.900 ;
        RECT 1318.020 3548.890 1321.020 3548.900 ;
        RECT 1498.020 3548.890 1501.020 3548.900 ;
        RECT 1678.020 3548.890 1681.020 3548.900 ;
        RECT 1858.020 3548.890 1861.020 3548.900 ;
        RECT 2038.020 3548.890 2041.020 3548.900 ;
        RECT 2218.020 3548.890 2221.020 3548.900 ;
        RECT 2398.020 3548.890 2401.020 3548.900 ;
        RECT 2578.020 3548.890 2581.020 3548.900 ;
        RECT 2758.020 3548.890 2761.020 3548.900 ;
        RECT 2954.200 3548.890 2957.200 3548.900 ;
        RECT -37.580 3486.380 -34.580 3486.390 ;
        RECT 58.020 3486.380 61.020 3486.390 ;
        RECT 238.020 3486.380 241.020 3486.390 ;
        RECT 418.020 3486.380 421.020 3486.390 ;
        RECT 598.020 3486.380 601.020 3486.390 ;
        RECT 778.020 3486.380 781.020 3486.390 ;
        RECT 958.020 3486.380 961.020 3486.390 ;
        RECT 1138.020 3486.380 1141.020 3486.390 ;
        RECT 1318.020 3486.380 1321.020 3486.390 ;
        RECT 1498.020 3486.380 1501.020 3486.390 ;
        RECT 1678.020 3486.380 1681.020 3486.390 ;
        RECT 1858.020 3486.380 1861.020 3486.390 ;
        RECT 2038.020 3486.380 2041.020 3486.390 ;
        RECT 2218.020 3486.380 2221.020 3486.390 ;
        RECT 2398.020 3486.380 2401.020 3486.390 ;
        RECT 2578.020 3486.380 2581.020 3486.390 ;
        RECT 2758.020 3486.380 2761.020 3486.390 ;
        RECT 2954.200 3486.380 2957.200 3486.390 ;
        RECT -42.180 3483.380 2961.800 3486.380 ;
        RECT -37.580 3483.370 -34.580 3483.380 ;
        RECT 58.020 3483.370 61.020 3483.380 ;
        RECT 238.020 3483.370 241.020 3483.380 ;
        RECT 418.020 3483.370 421.020 3483.380 ;
        RECT 598.020 3483.370 601.020 3483.380 ;
        RECT 778.020 3483.370 781.020 3483.380 ;
        RECT 958.020 3483.370 961.020 3483.380 ;
        RECT 1138.020 3483.370 1141.020 3483.380 ;
        RECT 1318.020 3483.370 1321.020 3483.380 ;
        RECT 1498.020 3483.370 1501.020 3483.380 ;
        RECT 1678.020 3483.370 1681.020 3483.380 ;
        RECT 1858.020 3483.370 1861.020 3483.380 ;
        RECT 2038.020 3483.370 2041.020 3483.380 ;
        RECT 2218.020 3483.370 2221.020 3483.380 ;
        RECT 2398.020 3483.370 2401.020 3483.380 ;
        RECT 2578.020 3483.370 2581.020 3483.380 ;
        RECT 2758.020 3483.370 2761.020 3483.380 ;
        RECT 2954.200 3483.370 2957.200 3483.380 ;
        RECT -37.580 3306.380 -34.580 3306.390 ;
        RECT 58.020 3306.380 61.020 3306.390 ;
        RECT 238.020 3306.380 241.020 3306.390 ;
        RECT 418.020 3306.380 421.020 3306.390 ;
        RECT 598.020 3306.380 601.020 3306.390 ;
        RECT 778.020 3306.380 781.020 3306.390 ;
        RECT 958.020 3306.380 961.020 3306.390 ;
        RECT 1138.020 3306.380 1141.020 3306.390 ;
        RECT 1318.020 3306.380 1321.020 3306.390 ;
        RECT 1498.020 3306.380 1501.020 3306.390 ;
        RECT 1678.020 3306.380 1681.020 3306.390 ;
        RECT 1858.020 3306.380 1861.020 3306.390 ;
        RECT 2038.020 3306.380 2041.020 3306.390 ;
        RECT 2218.020 3306.380 2221.020 3306.390 ;
        RECT 2398.020 3306.380 2401.020 3306.390 ;
        RECT 2578.020 3306.380 2581.020 3306.390 ;
        RECT 2758.020 3306.380 2761.020 3306.390 ;
        RECT 2954.200 3306.380 2957.200 3306.390 ;
        RECT -42.180 3303.380 2961.800 3306.380 ;
        RECT -37.580 3303.370 -34.580 3303.380 ;
        RECT 58.020 3303.370 61.020 3303.380 ;
        RECT 238.020 3303.370 241.020 3303.380 ;
        RECT 418.020 3303.370 421.020 3303.380 ;
        RECT 598.020 3303.370 601.020 3303.380 ;
        RECT 778.020 3303.370 781.020 3303.380 ;
        RECT 958.020 3303.370 961.020 3303.380 ;
        RECT 1138.020 3303.370 1141.020 3303.380 ;
        RECT 1318.020 3303.370 1321.020 3303.380 ;
        RECT 1498.020 3303.370 1501.020 3303.380 ;
        RECT 1678.020 3303.370 1681.020 3303.380 ;
        RECT 1858.020 3303.370 1861.020 3303.380 ;
        RECT 2038.020 3303.370 2041.020 3303.380 ;
        RECT 2218.020 3303.370 2221.020 3303.380 ;
        RECT 2398.020 3303.370 2401.020 3303.380 ;
        RECT 2578.020 3303.370 2581.020 3303.380 ;
        RECT 2758.020 3303.370 2761.020 3303.380 ;
        RECT 2954.200 3303.370 2957.200 3303.380 ;
        RECT -37.580 3126.380 -34.580 3126.390 ;
        RECT 58.020 3126.380 61.020 3126.390 ;
        RECT 238.020 3126.380 241.020 3126.390 ;
        RECT 418.020 3126.380 421.020 3126.390 ;
        RECT 598.020 3126.380 601.020 3126.390 ;
        RECT 778.020 3126.380 781.020 3126.390 ;
        RECT 958.020 3126.380 961.020 3126.390 ;
        RECT 1138.020 3126.380 1141.020 3126.390 ;
        RECT 1318.020 3126.380 1321.020 3126.390 ;
        RECT 1498.020 3126.380 1501.020 3126.390 ;
        RECT 1678.020 3126.380 1681.020 3126.390 ;
        RECT 1858.020 3126.380 1861.020 3126.390 ;
        RECT 2038.020 3126.380 2041.020 3126.390 ;
        RECT 2218.020 3126.380 2221.020 3126.390 ;
        RECT 2398.020 3126.380 2401.020 3126.390 ;
        RECT 2578.020 3126.380 2581.020 3126.390 ;
        RECT 2758.020 3126.380 2761.020 3126.390 ;
        RECT 2954.200 3126.380 2957.200 3126.390 ;
        RECT -42.180 3123.380 2961.800 3126.380 ;
        RECT -37.580 3123.370 -34.580 3123.380 ;
        RECT 58.020 3123.370 61.020 3123.380 ;
        RECT 238.020 3123.370 241.020 3123.380 ;
        RECT 418.020 3123.370 421.020 3123.380 ;
        RECT 598.020 3123.370 601.020 3123.380 ;
        RECT 778.020 3123.370 781.020 3123.380 ;
        RECT 958.020 3123.370 961.020 3123.380 ;
        RECT 1138.020 3123.370 1141.020 3123.380 ;
        RECT 1318.020 3123.370 1321.020 3123.380 ;
        RECT 1498.020 3123.370 1501.020 3123.380 ;
        RECT 1678.020 3123.370 1681.020 3123.380 ;
        RECT 1858.020 3123.370 1861.020 3123.380 ;
        RECT 2038.020 3123.370 2041.020 3123.380 ;
        RECT 2218.020 3123.370 2221.020 3123.380 ;
        RECT 2398.020 3123.370 2401.020 3123.380 ;
        RECT 2578.020 3123.370 2581.020 3123.380 ;
        RECT 2758.020 3123.370 2761.020 3123.380 ;
        RECT 2954.200 3123.370 2957.200 3123.380 ;
        RECT -37.580 2946.380 -34.580 2946.390 ;
        RECT 58.020 2946.380 61.020 2946.390 ;
        RECT 238.020 2946.380 241.020 2946.390 ;
        RECT 418.020 2946.380 421.020 2946.390 ;
        RECT 598.020 2946.380 601.020 2946.390 ;
        RECT 778.020 2946.380 781.020 2946.390 ;
        RECT 958.020 2946.380 961.020 2946.390 ;
        RECT 1138.020 2946.380 1141.020 2946.390 ;
        RECT 1318.020 2946.380 1321.020 2946.390 ;
        RECT 1498.020 2946.380 1501.020 2946.390 ;
        RECT 1678.020 2946.380 1681.020 2946.390 ;
        RECT 1858.020 2946.380 1861.020 2946.390 ;
        RECT 2038.020 2946.380 2041.020 2946.390 ;
        RECT 2218.020 2946.380 2221.020 2946.390 ;
        RECT 2398.020 2946.380 2401.020 2946.390 ;
        RECT 2578.020 2946.380 2581.020 2946.390 ;
        RECT 2758.020 2946.380 2761.020 2946.390 ;
        RECT 2954.200 2946.380 2957.200 2946.390 ;
        RECT -42.180 2943.380 2961.800 2946.380 ;
        RECT -37.580 2943.370 -34.580 2943.380 ;
        RECT 58.020 2943.370 61.020 2943.380 ;
        RECT 238.020 2943.370 241.020 2943.380 ;
        RECT 418.020 2943.370 421.020 2943.380 ;
        RECT 598.020 2943.370 601.020 2943.380 ;
        RECT 778.020 2943.370 781.020 2943.380 ;
        RECT 958.020 2943.370 961.020 2943.380 ;
        RECT 1138.020 2943.370 1141.020 2943.380 ;
        RECT 1318.020 2943.370 1321.020 2943.380 ;
        RECT 1498.020 2943.370 1501.020 2943.380 ;
        RECT 1678.020 2943.370 1681.020 2943.380 ;
        RECT 1858.020 2943.370 1861.020 2943.380 ;
        RECT 2038.020 2943.370 2041.020 2943.380 ;
        RECT 2218.020 2943.370 2221.020 2943.380 ;
        RECT 2398.020 2943.370 2401.020 2943.380 ;
        RECT 2578.020 2943.370 2581.020 2943.380 ;
        RECT 2758.020 2943.370 2761.020 2943.380 ;
        RECT 2954.200 2943.370 2957.200 2943.380 ;
        RECT -37.580 2766.380 -34.580 2766.390 ;
        RECT 58.020 2766.380 61.020 2766.390 ;
        RECT 238.020 2766.380 241.020 2766.390 ;
        RECT 418.020 2766.380 421.020 2766.390 ;
        RECT 598.020 2766.380 601.020 2766.390 ;
        RECT 778.020 2766.380 781.020 2766.390 ;
        RECT 958.020 2766.380 961.020 2766.390 ;
        RECT 1138.020 2766.380 1141.020 2766.390 ;
        RECT 1318.020 2766.380 1321.020 2766.390 ;
        RECT 1498.020 2766.380 1501.020 2766.390 ;
        RECT 1678.020 2766.380 1681.020 2766.390 ;
        RECT 1858.020 2766.380 1861.020 2766.390 ;
        RECT 2038.020 2766.380 2041.020 2766.390 ;
        RECT 2218.020 2766.380 2221.020 2766.390 ;
        RECT 2398.020 2766.380 2401.020 2766.390 ;
        RECT 2578.020 2766.380 2581.020 2766.390 ;
        RECT 2758.020 2766.380 2761.020 2766.390 ;
        RECT 2954.200 2766.380 2957.200 2766.390 ;
        RECT -42.180 2763.380 2961.800 2766.380 ;
        RECT -37.580 2763.370 -34.580 2763.380 ;
        RECT 58.020 2763.370 61.020 2763.380 ;
        RECT 238.020 2763.370 241.020 2763.380 ;
        RECT 418.020 2763.370 421.020 2763.380 ;
        RECT 598.020 2763.370 601.020 2763.380 ;
        RECT 778.020 2763.370 781.020 2763.380 ;
        RECT 958.020 2763.370 961.020 2763.380 ;
        RECT 1138.020 2763.370 1141.020 2763.380 ;
        RECT 1318.020 2763.370 1321.020 2763.380 ;
        RECT 1498.020 2763.370 1501.020 2763.380 ;
        RECT 1678.020 2763.370 1681.020 2763.380 ;
        RECT 1858.020 2763.370 1861.020 2763.380 ;
        RECT 2038.020 2763.370 2041.020 2763.380 ;
        RECT 2218.020 2763.370 2221.020 2763.380 ;
        RECT 2398.020 2763.370 2401.020 2763.380 ;
        RECT 2578.020 2763.370 2581.020 2763.380 ;
        RECT 2758.020 2763.370 2761.020 2763.380 ;
        RECT 2954.200 2763.370 2957.200 2763.380 ;
        RECT -37.580 2586.380 -34.580 2586.390 ;
        RECT 58.020 2586.380 61.020 2586.390 ;
        RECT 238.020 2586.380 241.020 2586.390 ;
        RECT 418.020 2586.380 421.020 2586.390 ;
        RECT 598.020 2586.380 601.020 2586.390 ;
        RECT 778.020 2586.380 781.020 2586.390 ;
        RECT 958.020 2586.380 961.020 2586.390 ;
        RECT 1138.020 2586.380 1141.020 2586.390 ;
        RECT 1318.020 2586.380 1321.020 2586.390 ;
        RECT 1498.020 2586.380 1501.020 2586.390 ;
        RECT 1678.020 2586.380 1681.020 2586.390 ;
        RECT 1858.020 2586.380 1861.020 2586.390 ;
        RECT 2038.020 2586.380 2041.020 2586.390 ;
        RECT 2218.020 2586.380 2221.020 2586.390 ;
        RECT 2398.020 2586.380 2401.020 2586.390 ;
        RECT 2578.020 2586.380 2581.020 2586.390 ;
        RECT 2758.020 2586.380 2761.020 2586.390 ;
        RECT 2954.200 2586.380 2957.200 2586.390 ;
        RECT -42.180 2583.380 2961.800 2586.380 ;
        RECT -37.580 2583.370 -34.580 2583.380 ;
        RECT 58.020 2583.370 61.020 2583.380 ;
        RECT 238.020 2583.370 241.020 2583.380 ;
        RECT 418.020 2583.370 421.020 2583.380 ;
        RECT 598.020 2583.370 601.020 2583.380 ;
        RECT 778.020 2583.370 781.020 2583.380 ;
        RECT 958.020 2583.370 961.020 2583.380 ;
        RECT 1138.020 2583.370 1141.020 2583.380 ;
        RECT 1318.020 2583.370 1321.020 2583.380 ;
        RECT 1498.020 2583.370 1501.020 2583.380 ;
        RECT 1678.020 2583.370 1681.020 2583.380 ;
        RECT 1858.020 2583.370 1861.020 2583.380 ;
        RECT 2038.020 2583.370 2041.020 2583.380 ;
        RECT 2218.020 2583.370 2221.020 2583.380 ;
        RECT 2398.020 2583.370 2401.020 2583.380 ;
        RECT 2578.020 2583.370 2581.020 2583.380 ;
        RECT 2758.020 2583.370 2761.020 2583.380 ;
        RECT 2954.200 2583.370 2957.200 2583.380 ;
        RECT -37.580 2406.380 -34.580 2406.390 ;
        RECT 58.020 2406.380 61.020 2406.390 ;
        RECT 238.020 2406.380 241.020 2406.390 ;
        RECT 418.020 2406.380 421.020 2406.390 ;
        RECT 598.020 2406.380 601.020 2406.390 ;
        RECT 778.020 2406.380 781.020 2406.390 ;
        RECT 958.020 2406.380 961.020 2406.390 ;
        RECT 1138.020 2406.380 1141.020 2406.390 ;
        RECT 1318.020 2406.380 1321.020 2406.390 ;
        RECT 1498.020 2406.380 1501.020 2406.390 ;
        RECT 1678.020 2406.380 1681.020 2406.390 ;
        RECT 1858.020 2406.380 1861.020 2406.390 ;
        RECT 2038.020 2406.380 2041.020 2406.390 ;
        RECT 2218.020 2406.380 2221.020 2406.390 ;
        RECT 2398.020 2406.380 2401.020 2406.390 ;
        RECT 2578.020 2406.380 2581.020 2406.390 ;
        RECT 2758.020 2406.380 2761.020 2406.390 ;
        RECT 2954.200 2406.380 2957.200 2406.390 ;
        RECT -42.180 2403.380 2961.800 2406.380 ;
        RECT -37.580 2403.370 -34.580 2403.380 ;
        RECT 58.020 2403.370 61.020 2403.380 ;
        RECT 238.020 2403.370 241.020 2403.380 ;
        RECT 418.020 2403.370 421.020 2403.380 ;
        RECT 598.020 2403.370 601.020 2403.380 ;
        RECT 778.020 2403.370 781.020 2403.380 ;
        RECT 958.020 2403.370 961.020 2403.380 ;
        RECT 1138.020 2403.370 1141.020 2403.380 ;
        RECT 1318.020 2403.370 1321.020 2403.380 ;
        RECT 1498.020 2403.370 1501.020 2403.380 ;
        RECT 1678.020 2403.370 1681.020 2403.380 ;
        RECT 1858.020 2403.370 1861.020 2403.380 ;
        RECT 2038.020 2403.370 2041.020 2403.380 ;
        RECT 2218.020 2403.370 2221.020 2403.380 ;
        RECT 2398.020 2403.370 2401.020 2403.380 ;
        RECT 2578.020 2403.370 2581.020 2403.380 ;
        RECT 2758.020 2403.370 2761.020 2403.380 ;
        RECT 2954.200 2403.370 2957.200 2403.380 ;
        RECT -37.580 2226.380 -34.580 2226.390 ;
        RECT 58.020 2226.380 61.020 2226.390 ;
        RECT 238.020 2226.380 241.020 2226.390 ;
        RECT 418.020 2226.380 421.020 2226.390 ;
        RECT 598.020 2226.380 601.020 2226.390 ;
        RECT 778.020 2226.380 781.020 2226.390 ;
        RECT 958.020 2226.380 961.020 2226.390 ;
        RECT 1138.020 2226.380 1141.020 2226.390 ;
        RECT 1318.020 2226.380 1321.020 2226.390 ;
        RECT 1498.020 2226.380 1501.020 2226.390 ;
        RECT 1678.020 2226.380 1681.020 2226.390 ;
        RECT 1858.020 2226.380 1861.020 2226.390 ;
        RECT 2038.020 2226.380 2041.020 2226.390 ;
        RECT 2218.020 2226.380 2221.020 2226.390 ;
        RECT 2398.020 2226.380 2401.020 2226.390 ;
        RECT 2578.020 2226.380 2581.020 2226.390 ;
        RECT 2758.020 2226.380 2761.020 2226.390 ;
        RECT 2954.200 2226.380 2957.200 2226.390 ;
        RECT -42.180 2223.380 2961.800 2226.380 ;
        RECT -37.580 2223.370 -34.580 2223.380 ;
        RECT 58.020 2223.370 61.020 2223.380 ;
        RECT 238.020 2223.370 241.020 2223.380 ;
        RECT 418.020 2223.370 421.020 2223.380 ;
        RECT 598.020 2223.370 601.020 2223.380 ;
        RECT 778.020 2223.370 781.020 2223.380 ;
        RECT 958.020 2223.370 961.020 2223.380 ;
        RECT 1138.020 2223.370 1141.020 2223.380 ;
        RECT 1318.020 2223.370 1321.020 2223.380 ;
        RECT 1498.020 2223.370 1501.020 2223.380 ;
        RECT 1678.020 2223.370 1681.020 2223.380 ;
        RECT 1858.020 2223.370 1861.020 2223.380 ;
        RECT 2038.020 2223.370 2041.020 2223.380 ;
        RECT 2218.020 2223.370 2221.020 2223.380 ;
        RECT 2398.020 2223.370 2401.020 2223.380 ;
        RECT 2578.020 2223.370 2581.020 2223.380 ;
        RECT 2758.020 2223.370 2761.020 2223.380 ;
        RECT 2954.200 2223.370 2957.200 2223.380 ;
        RECT -37.580 2046.380 -34.580 2046.390 ;
        RECT 58.020 2046.380 61.020 2046.390 ;
        RECT 238.020 2046.380 241.020 2046.390 ;
        RECT 418.020 2046.380 421.020 2046.390 ;
        RECT 598.020 2046.380 601.020 2046.390 ;
        RECT 778.020 2046.380 781.020 2046.390 ;
        RECT 958.020 2046.380 961.020 2046.390 ;
        RECT 1138.020 2046.380 1141.020 2046.390 ;
        RECT 1318.020 2046.380 1321.020 2046.390 ;
        RECT 1498.020 2046.380 1501.020 2046.390 ;
        RECT 1678.020 2046.380 1681.020 2046.390 ;
        RECT 1858.020 2046.380 1861.020 2046.390 ;
        RECT 2038.020 2046.380 2041.020 2046.390 ;
        RECT 2218.020 2046.380 2221.020 2046.390 ;
        RECT 2398.020 2046.380 2401.020 2046.390 ;
        RECT 2578.020 2046.380 2581.020 2046.390 ;
        RECT 2758.020 2046.380 2761.020 2046.390 ;
        RECT 2954.200 2046.380 2957.200 2046.390 ;
        RECT -42.180 2043.380 2961.800 2046.380 ;
        RECT -37.580 2043.370 -34.580 2043.380 ;
        RECT 58.020 2043.370 61.020 2043.380 ;
        RECT 238.020 2043.370 241.020 2043.380 ;
        RECT 418.020 2043.370 421.020 2043.380 ;
        RECT 598.020 2043.370 601.020 2043.380 ;
        RECT 778.020 2043.370 781.020 2043.380 ;
        RECT 958.020 2043.370 961.020 2043.380 ;
        RECT 1138.020 2043.370 1141.020 2043.380 ;
        RECT 1318.020 2043.370 1321.020 2043.380 ;
        RECT 1498.020 2043.370 1501.020 2043.380 ;
        RECT 1678.020 2043.370 1681.020 2043.380 ;
        RECT 1858.020 2043.370 1861.020 2043.380 ;
        RECT 2038.020 2043.370 2041.020 2043.380 ;
        RECT 2218.020 2043.370 2221.020 2043.380 ;
        RECT 2398.020 2043.370 2401.020 2043.380 ;
        RECT 2578.020 2043.370 2581.020 2043.380 ;
        RECT 2758.020 2043.370 2761.020 2043.380 ;
        RECT 2954.200 2043.370 2957.200 2043.380 ;
        RECT -37.580 1866.380 -34.580 1866.390 ;
        RECT 58.020 1866.380 61.020 1866.390 ;
        RECT 238.020 1866.380 241.020 1866.390 ;
        RECT 418.020 1866.380 421.020 1866.390 ;
        RECT 598.020 1866.380 601.020 1866.390 ;
        RECT 778.020 1866.380 781.020 1866.390 ;
        RECT 958.020 1866.380 961.020 1866.390 ;
        RECT 1138.020 1866.380 1141.020 1866.390 ;
        RECT 1318.020 1866.380 1321.020 1866.390 ;
        RECT 1498.020 1866.380 1501.020 1866.390 ;
        RECT 1678.020 1866.380 1681.020 1866.390 ;
        RECT 1858.020 1866.380 1861.020 1866.390 ;
        RECT 2038.020 1866.380 2041.020 1866.390 ;
        RECT 2218.020 1866.380 2221.020 1866.390 ;
        RECT 2398.020 1866.380 2401.020 1866.390 ;
        RECT 2578.020 1866.380 2581.020 1866.390 ;
        RECT 2758.020 1866.380 2761.020 1866.390 ;
        RECT 2954.200 1866.380 2957.200 1866.390 ;
        RECT -42.180 1863.380 2961.800 1866.380 ;
        RECT -37.580 1863.370 -34.580 1863.380 ;
        RECT 58.020 1863.370 61.020 1863.380 ;
        RECT 238.020 1863.370 241.020 1863.380 ;
        RECT 418.020 1863.370 421.020 1863.380 ;
        RECT 598.020 1863.370 601.020 1863.380 ;
        RECT 778.020 1863.370 781.020 1863.380 ;
        RECT 958.020 1863.370 961.020 1863.380 ;
        RECT 1138.020 1863.370 1141.020 1863.380 ;
        RECT 1318.020 1863.370 1321.020 1863.380 ;
        RECT 1498.020 1863.370 1501.020 1863.380 ;
        RECT 1678.020 1863.370 1681.020 1863.380 ;
        RECT 1858.020 1863.370 1861.020 1863.380 ;
        RECT 2038.020 1863.370 2041.020 1863.380 ;
        RECT 2218.020 1863.370 2221.020 1863.380 ;
        RECT 2398.020 1863.370 2401.020 1863.380 ;
        RECT 2578.020 1863.370 2581.020 1863.380 ;
        RECT 2758.020 1863.370 2761.020 1863.380 ;
        RECT 2954.200 1863.370 2957.200 1863.380 ;
        RECT -37.580 1686.380 -34.580 1686.390 ;
        RECT 58.020 1686.380 61.020 1686.390 ;
        RECT 238.020 1686.380 241.020 1686.390 ;
        RECT 418.020 1686.380 421.020 1686.390 ;
        RECT 598.020 1686.380 601.020 1686.390 ;
        RECT 778.020 1686.380 781.020 1686.390 ;
        RECT 958.020 1686.380 961.020 1686.390 ;
        RECT 1138.020 1686.380 1141.020 1686.390 ;
        RECT 1318.020 1686.380 1321.020 1686.390 ;
        RECT 1498.020 1686.380 1501.020 1686.390 ;
        RECT 1678.020 1686.380 1681.020 1686.390 ;
        RECT 1858.020 1686.380 1861.020 1686.390 ;
        RECT 2038.020 1686.380 2041.020 1686.390 ;
        RECT 2218.020 1686.380 2221.020 1686.390 ;
        RECT 2398.020 1686.380 2401.020 1686.390 ;
        RECT 2578.020 1686.380 2581.020 1686.390 ;
        RECT 2758.020 1686.380 2761.020 1686.390 ;
        RECT 2954.200 1686.380 2957.200 1686.390 ;
        RECT -42.180 1683.380 2961.800 1686.380 ;
        RECT -37.580 1683.370 -34.580 1683.380 ;
        RECT 58.020 1683.370 61.020 1683.380 ;
        RECT 238.020 1683.370 241.020 1683.380 ;
        RECT 418.020 1683.370 421.020 1683.380 ;
        RECT 598.020 1683.370 601.020 1683.380 ;
        RECT 778.020 1683.370 781.020 1683.380 ;
        RECT 958.020 1683.370 961.020 1683.380 ;
        RECT 1138.020 1683.370 1141.020 1683.380 ;
        RECT 1318.020 1683.370 1321.020 1683.380 ;
        RECT 1498.020 1683.370 1501.020 1683.380 ;
        RECT 1678.020 1683.370 1681.020 1683.380 ;
        RECT 1858.020 1683.370 1861.020 1683.380 ;
        RECT 2038.020 1683.370 2041.020 1683.380 ;
        RECT 2218.020 1683.370 2221.020 1683.380 ;
        RECT 2398.020 1683.370 2401.020 1683.380 ;
        RECT 2578.020 1683.370 2581.020 1683.380 ;
        RECT 2758.020 1683.370 2761.020 1683.380 ;
        RECT 2954.200 1683.370 2957.200 1683.380 ;
        RECT -37.580 1506.380 -34.580 1506.390 ;
        RECT 58.020 1506.380 61.020 1506.390 ;
        RECT 238.020 1506.380 241.020 1506.390 ;
        RECT 418.020 1506.380 421.020 1506.390 ;
        RECT 598.020 1506.380 601.020 1506.390 ;
        RECT 778.020 1506.380 781.020 1506.390 ;
        RECT 958.020 1506.380 961.020 1506.390 ;
        RECT 1138.020 1506.380 1141.020 1506.390 ;
        RECT 1318.020 1506.380 1321.020 1506.390 ;
        RECT 1498.020 1506.380 1501.020 1506.390 ;
        RECT 1678.020 1506.380 1681.020 1506.390 ;
        RECT 1858.020 1506.380 1861.020 1506.390 ;
        RECT 2038.020 1506.380 2041.020 1506.390 ;
        RECT 2218.020 1506.380 2221.020 1506.390 ;
        RECT 2398.020 1506.380 2401.020 1506.390 ;
        RECT 2578.020 1506.380 2581.020 1506.390 ;
        RECT 2758.020 1506.380 2761.020 1506.390 ;
        RECT 2954.200 1506.380 2957.200 1506.390 ;
        RECT -42.180 1503.380 2961.800 1506.380 ;
        RECT -37.580 1503.370 -34.580 1503.380 ;
        RECT 58.020 1503.370 61.020 1503.380 ;
        RECT 238.020 1503.370 241.020 1503.380 ;
        RECT 418.020 1503.370 421.020 1503.380 ;
        RECT 598.020 1503.370 601.020 1503.380 ;
        RECT 778.020 1503.370 781.020 1503.380 ;
        RECT 958.020 1503.370 961.020 1503.380 ;
        RECT 1138.020 1503.370 1141.020 1503.380 ;
        RECT 1318.020 1503.370 1321.020 1503.380 ;
        RECT 1498.020 1503.370 1501.020 1503.380 ;
        RECT 1678.020 1503.370 1681.020 1503.380 ;
        RECT 1858.020 1503.370 1861.020 1503.380 ;
        RECT 2038.020 1503.370 2041.020 1503.380 ;
        RECT 2218.020 1503.370 2221.020 1503.380 ;
        RECT 2398.020 1503.370 2401.020 1503.380 ;
        RECT 2578.020 1503.370 2581.020 1503.380 ;
        RECT 2758.020 1503.370 2761.020 1503.380 ;
        RECT 2954.200 1503.370 2957.200 1503.380 ;
        RECT -37.580 1326.380 -34.580 1326.390 ;
        RECT 58.020 1326.380 61.020 1326.390 ;
        RECT 238.020 1326.380 241.020 1326.390 ;
        RECT 418.020 1326.380 421.020 1326.390 ;
        RECT 598.020 1326.380 601.020 1326.390 ;
        RECT 778.020 1326.380 781.020 1326.390 ;
        RECT 958.020 1326.380 961.020 1326.390 ;
        RECT 1138.020 1326.380 1141.020 1326.390 ;
        RECT 1318.020 1326.380 1321.020 1326.390 ;
        RECT 1498.020 1326.380 1501.020 1326.390 ;
        RECT 1678.020 1326.380 1681.020 1326.390 ;
        RECT 1858.020 1326.380 1861.020 1326.390 ;
        RECT 2038.020 1326.380 2041.020 1326.390 ;
        RECT 2218.020 1326.380 2221.020 1326.390 ;
        RECT 2398.020 1326.380 2401.020 1326.390 ;
        RECT 2578.020 1326.380 2581.020 1326.390 ;
        RECT 2758.020 1326.380 2761.020 1326.390 ;
        RECT 2954.200 1326.380 2957.200 1326.390 ;
        RECT -42.180 1323.380 2961.800 1326.380 ;
        RECT -37.580 1323.370 -34.580 1323.380 ;
        RECT 58.020 1323.370 61.020 1323.380 ;
        RECT 238.020 1323.370 241.020 1323.380 ;
        RECT 418.020 1323.370 421.020 1323.380 ;
        RECT 598.020 1323.370 601.020 1323.380 ;
        RECT 778.020 1323.370 781.020 1323.380 ;
        RECT 958.020 1323.370 961.020 1323.380 ;
        RECT 1138.020 1323.370 1141.020 1323.380 ;
        RECT 1318.020 1323.370 1321.020 1323.380 ;
        RECT 1498.020 1323.370 1501.020 1323.380 ;
        RECT 1678.020 1323.370 1681.020 1323.380 ;
        RECT 1858.020 1323.370 1861.020 1323.380 ;
        RECT 2038.020 1323.370 2041.020 1323.380 ;
        RECT 2218.020 1323.370 2221.020 1323.380 ;
        RECT 2398.020 1323.370 2401.020 1323.380 ;
        RECT 2578.020 1323.370 2581.020 1323.380 ;
        RECT 2758.020 1323.370 2761.020 1323.380 ;
        RECT 2954.200 1323.370 2957.200 1323.380 ;
        RECT -37.580 1146.380 -34.580 1146.390 ;
        RECT 58.020 1146.380 61.020 1146.390 ;
        RECT 238.020 1146.380 241.020 1146.390 ;
        RECT 418.020 1146.380 421.020 1146.390 ;
        RECT 598.020 1146.380 601.020 1146.390 ;
        RECT 778.020 1146.380 781.020 1146.390 ;
        RECT 958.020 1146.380 961.020 1146.390 ;
        RECT 1138.020 1146.380 1141.020 1146.390 ;
        RECT 1318.020 1146.380 1321.020 1146.390 ;
        RECT 1498.020 1146.380 1501.020 1146.390 ;
        RECT 1678.020 1146.380 1681.020 1146.390 ;
        RECT 1858.020 1146.380 1861.020 1146.390 ;
        RECT 2038.020 1146.380 2041.020 1146.390 ;
        RECT 2218.020 1146.380 2221.020 1146.390 ;
        RECT 2398.020 1146.380 2401.020 1146.390 ;
        RECT 2578.020 1146.380 2581.020 1146.390 ;
        RECT 2758.020 1146.380 2761.020 1146.390 ;
        RECT 2954.200 1146.380 2957.200 1146.390 ;
        RECT -42.180 1143.380 2961.800 1146.380 ;
        RECT -37.580 1143.370 -34.580 1143.380 ;
        RECT 58.020 1143.370 61.020 1143.380 ;
        RECT 238.020 1143.370 241.020 1143.380 ;
        RECT 418.020 1143.370 421.020 1143.380 ;
        RECT 598.020 1143.370 601.020 1143.380 ;
        RECT 778.020 1143.370 781.020 1143.380 ;
        RECT 958.020 1143.370 961.020 1143.380 ;
        RECT 1138.020 1143.370 1141.020 1143.380 ;
        RECT 1318.020 1143.370 1321.020 1143.380 ;
        RECT 1498.020 1143.370 1501.020 1143.380 ;
        RECT 1678.020 1143.370 1681.020 1143.380 ;
        RECT 1858.020 1143.370 1861.020 1143.380 ;
        RECT 2038.020 1143.370 2041.020 1143.380 ;
        RECT 2218.020 1143.370 2221.020 1143.380 ;
        RECT 2398.020 1143.370 2401.020 1143.380 ;
        RECT 2578.020 1143.370 2581.020 1143.380 ;
        RECT 2758.020 1143.370 2761.020 1143.380 ;
        RECT 2954.200 1143.370 2957.200 1143.380 ;
        RECT -37.580 966.380 -34.580 966.390 ;
        RECT 58.020 966.380 61.020 966.390 ;
        RECT 238.020 966.380 241.020 966.390 ;
        RECT 418.020 966.380 421.020 966.390 ;
        RECT 598.020 966.380 601.020 966.390 ;
        RECT 778.020 966.380 781.020 966.390 ;
        RECT 958.020 966.380 961.020 966.390 ;
        RECT 1138.020 966.380 1141.020 966.390 ;
        RECT 1318.020 966.380 1321.020 966.390 ;
        RECT 1498.020 966.380 1501.020 966.390 ;
        RECT 1678.020 966.380 1681.020 966.390 ;
        RECT 1858.020 966.380 1861.020 966.390 ;
        RECT 2038.020 966.380 2041.020 966.390 ;
        RECT 2218.020 966.380 2221.020 966.390 ;
        RECT 2398.020 966.380 2401.020 966.390 ;
        RECT 2578.020 966.380 2581.020 966.390 ;
        RECT 2758.020 966.380 2761.020 966.390 ;
        RECT 2954.200 966.380 2957.200 966.390 ;
        RECT -42.180 963.380 2961.800 966.380 ;
        RECT -37.580 963.370 -34.580 963.380 ;
        RECT 58.020 963.370 61.020 963.380 ;
        RECT 238.020 963.370 241.020 963.380 ;
        RECT 418.020 963.370 421.020 963.380 ;
        RECT 598.020 963.370 601.020 963.380 ;
        RECT 778.020 963.370 781.020 963.380 ;
        RECT 958.020 963.370 961.020 963.380 ;
        RECT 1138.020 963.370 1141.020 963.380 ;
        RECT 1318.020 963.370 1321.020 963.380 ;
        RECT 1498.020 963.370 1501.020 963.380 ;
        RECT 1678.020 963.370 1681.020 963.380 ;
        RECT 1858.020 963.370 1861.020 963.380 ;
        RECT 2038.020 963.370 2041.020 963.380 ;
        RECT 2218.020 963.370 2221.020 963.380 ;
        RECT 2398.020 963.370 2401.020 963.380 ;
        RECT 2578.020 963.370 2581.020 963.380 ;
        RECT 2758.020 963.370 2761.020 963.380 ;
        RECT 2954.200 963.370 2957.200 963.380 ;
        RECT -37.580 786.380 -34.580 786.390 ;
        RECT 58.020 786.380 61.020 786.390 ;
        RECT 238.020 786.380 241.020 786.390 ;
        RECT 418.020 786.380 421.020 786.390 ;
        RECT 598.020 786.380 601.020 786.390 ;
        RECT 778.020 786.380 781.020 786.390 ;
        RECT 958.020 786.380 961.020 786.390 ;
        RECT 1138.020 786.380 1141.020 786.390 ;
        RECT 1318.020 786.380 1321.020 786.390 ;
        RECT 1498.020 786.380 1501.020 786.390 ;
        RECT 1678.020 786.380 1681.020 786.390 ;
        RECT 1858.020 786.380 1861.020 786.390 ;
        RECT 2038.020 786.380 2041.020 786.390 ;
        RECT 2218.020 786.380 2221.020 786.390 ;
        RECT 2398.020 786.380 2401.020 786.390 ;
        RECT 2578.020 786.380 2581.020 786.390 ;
        RECT 2758.020 786.380 2761.020 786.390 ;
        RECT 2954.200 786.380 2957.200 786.390 ;
        RECT -42.180 783.380 2961.800 786.380 ;
        RECT -37.580 783.370 -34.580 783.380 ;
        RECT 58.020 783.370 61.020 783.380 ;
        RECT 238.020 783.370 241.020 783.380 ;
        RECT 418.020 783.370 421.020 783.380 ;
        RECT 598.020 783.370 601.020 783.380 ;
        RECT 778.020 783.370 781.020 783.380 ;
        RECT 958.020 783.370 961.020 783.380 ;
        RECT 1138.020 783.370 1141.020 783.380 ;
        RECT 1318.020 783.370 1321.020 783.380 ;
        RECT 1498.020 783.370 1501.020 783.380 ;
        RECT 1678.020 783.370 1681.020 783.380 ;
        RECT 1858.020 783.370 1861.020 783.380 ;
        RECT 2038.020 783.370 2041.020 783.380 ;
        RECT 2218.020 783.370 2221.020 783.380 ;
        RECT 2398.020 783.370 2401.020 783.380 ;
        RECT 2578.020 783.370 2581.020 783.380 ;
        RECT 2758.020 783.370 2761.020 783.380 ;
        RECT 2954.200 783.370 2957.200 783.380 ;
        RECT -37.580 606.380 -34.580 606.390 ;
        RECT 58.020 606.380 61.020 606.390 ;
        RECT 238.020 606.380 241.020 606.390 ;
        RECT 418.020 606.380 421.020 606.390 ;
        RECT 598.020 606.380 601.020 606.390 ;
        RECT 778.020 606.380 781.020 606.390 ;
        RECT 958.020 606.380 961.020 606.390 ;
        RECT 1138.020 606.380 1141.020 606.390 ;
        RECT 1318.020 606.380 1321.020 606.390 ;
        RECT 1498.020 606.380 1501.020 606.390 ;
        RECT 1678.020 606.380 1681.020 606.390 ;
        RECT 1858.020 606.380 1861.020 606.390 ;
        RECT 2038.020 606.380 2041.020 606.390 ;
        RECT 2218.020 606.380 2221.020 606.390 ;
        RECT 2398.020 606.380 2401.020 606.390 ;
        RECT 2578.020 606.380 2581.020 606.390 ;
        RECT 2758.020 606.380 2761.020 606.390 ;
        RECT 2954.200 606.380 2957.200 606.390 ;
        RECT -42.180 603.380 2961.800 606.380 ;
        RECT -37.580 603.370 -34.580 603.380 ;
        RECT 58.020 603.370 61.020 603.380 ;
        RECT 238.020 603.370 241.020 603.380 ;
        RECT 418.020 603.370 421.020 603.380 ;
        RECT 598.020 603.370 601.020 603.380 ;
        RECT 778.020 603.370 781.020 603.380 ;
        RECT 958.020 603.370 961.020 603.380 ;
        RECT 1138.020 603.370 1141.020 603.380 ;
        RECT 1318.020 603.370 1321.020 603.380 ;
        RECT 1498.020 603.370 1501.020 603.380 ;
        RECT 1678.020 603.370 1681.020 603.380 ;
        RECT 1858.020 603.370 1861.020 603.380 ;
        RECT 2038.020 603.370 2041.020 603.380 ;
        RECT 2218.020 603.370 2221.020 603.380 ;
        RECT 2398.020 603.370 2401.020 603.380 ;
        RECT 2578.020 603.370 2581.020 603.380 ;
        RECT 2758.020 603.370 2761.020 603.380 ;
        RECT 2954.200 603.370 2957.200 603.380 ;
        RECT -37.580 426.380 -34.580 426.390 ;
        RECT 58.020 426.380 61.020 426.390 ;
        RECT 238.020 426.380 241.020 426.390 ;
        RECT 418.020 426.380 421.020 426.390 ;
        RECT 598.020 426.380 601.020 426.390 ;
        RECT 778.020 426.380 781.020 426.390 ;
        RECT 958.020 426.380 961.020 426.390 ;
        RECT 1138.020 426.380 1141.020 426.390 ;
        RECT 1318.020 426.380 1321.020 426.390 ;
        RECT 1498.020 426.380 1501.020 426.390 ;
        RECT 1678.020 426.380 1681.020 426.390 ;
        RECT 1858.020 426.380 1861.020 426.390 ;
        RECT 2038.020 426.380 2041.020 426.390 ;
        RECT 2218.020 426.380 2221.020 426.390 ;
        RECT 2398.020 426.380 2401.020 426.390 ;
        RECT 2578.020 426.380 2581.020 426.390 ;
        RECT 2758.020 426.380 2761.020 426.390 ;
        RECT 2954.200 426.380 2957.200 426.390 ;
        RECT -42.180 423.380 2961.800 426.380 ;
        RECT -37.580 423.370 -34.580 423.380 ;
        RECT 58.020 423.370 61.020 423.380 ;
        RECT 238.020 423.370 241.020 423.380 ;
        RECT 418.020 423.370 421.020 423.380 ;
        RECT 598.020 423.370 601.020 423.380 ;
        RECT 778.020 423.370 781.020 423.380 ;
        RECT 958.020 423.370 961.020 423.380 ;
        RECT 1138.020 423.370 1141.020 423.380 ;
        RECT 1318.020 423.370 1321.020 423.380 ;
        RECT 1498.020 423.370 1501.020 423.380 ;
        RECT 1678.020 423.370 1681.020 423.380 ;
        RECT 1858.020 423.370 1861.020 423.380 ;
        RECT 2038.020 423.370 2041.020 423.380 ;
        RECT 2218.020 423.370 2221.020 423.380 ;
        RECT 2398.020 423.370 2401.020 423.380 ;
        RECT 2578.020 423.370 2581.020 423.380 ;
        RECT 2758.020 423.370 2761.020 423.380 ;
        RECT 2954.200 423.370 2957.200 423.380 ;
        RECT -37.580 246.380 -34.580 246.390 ;
        RECT 58.020 246.380 61.020 246.390 ;
        RECT 238.020 246.380 241.020 246.390 ;
        RECT 418.020 246.380 421.020 246.390 ;
        RECT 598.020 246.380 601.020 246.390 ;
        RECT 778.020 246.380 781.020 246.390 ;
        RECT 958.020 246.380 961.020 246.390 ;
        RECT 1138.020 246.380 1141.020 246.390 ;
        RECT 1318.020 246.380 1321.020 246.390 ;
        RECT 1498.020 246.380 1501.020 246.390 ;
        RECT 1678.020 246.380 1681.020 246.390 ;
        RECT 1858.020 246.380 1861.020 246.390 ;
        RECT 2038.020 246.380 2041.020 246.390 ;
        RECT 2218.020 246.380 2221.020 246.390 ;
        RECT 2398.020 246.380 2401.020 246.390 ;
        RECT 2578.020 246.380 2581.020 246.390 ;
        RECT 2758.020 246.380 2761.020 246.390 ;
        RECT 2954.200 246.380 2957.200 246.390 ;
        RECT -42.180 243.380 2961.800 246.380 ;
        RECT -37.580 243.370 -34.580 243.380 ;
        RECT 58.020 243.370 61.020 243.380 ;
        RECT 238.020 243.370 241.020 243.380 ;
        RECT 418.020 243.370 421.020 243.380 ;
        RECT 598.020 243.370 601.020 243.380 ;
        RECT 778.020 243.370 781.020 243.380 ;
        RECT 958.020 243.370 961.020 243.380 ;
        RECT 1138.020 243.370 1141.020 243.380 ;
        RECT 1318.020 243.370 1321.020 243.380 ;
        RECT 1498.020 243.370 1501.020 243.380 ;
        RECT 1678.020 243.370 1681.020 243.380 ;
        RECT 1858.020 243.370 1861.020 243.380 ;
        RECT 2038.020 243.370 2041.020 243.380 ;
        RECT 2218.020 243.370 2221.020 243.380 ;
        RECT 2398.020 243.370 2401.020 243.380 ;
        RECT 2578.020 243.370 2581.020 243.380 ;
        RECT 2758.020 243.370 2761.020 243.380 ;
        RECT 2954.200 243.370 2957.200 243.380 ;
        RECT -37.580 66.380 -34.580 66.390 ;
        RECT 58.020 66.380 61.020 66.390 ;
        RECT 238.020 66.380 241.020 66.390 ;
        RECT 418.020 66.380 421.020 66.390 ;
        RECT 598.020 66.380 601.020 66.390 ;
        RECT 778.020 66.380 781.020 66.390 ;
        RECT 958.020 66.380 961.020 66.390 ;
        RECT 1138.020 66.380 1141.020 66.390 ;
        RECT 1318.020 66.380 1321.020 66.390 ;
        RECT 1498.020 66.380 1501.020 66.390 ;
        RECT 1678.020 66.380 1681.020 66.390 ;
        RECT 1858.020 66.380 1861.020 66.390 ;
        RECT 2038.020 66.380 2041.020 66.390 ;
        RECT 2218.020 66.380 2221.020 66.390 ;
        RECT 2398.020 66.380 2401.020 66.390 ;
        RECT 2578.020 66.380 2581.020 66.390 ;
        RECT 2758.020 66.380 2761.020 66.390 ;
        RECT 2954.200 66.380 2957.200 66.390 ;
        RECT -42.180 63.380 2961.800 66.380 ;
        RECT -37.580 63.370 -34.580 63.380 ;
        RECT 58.020 63.370 61.020 63.380 ;
        RECT 238.020 63.370 241.020 63.380 ;
        RECT 418.020 63.370 421.020 63.380 ;
        RECT 598.020 63.370 601.020 63.380 ;
        RECT 778.020 63.370 781.020 63.380 ;
        RECT 958.020 63.370 961.020 63.380 ;
        RECT 1138.020 63.370 1141.020 63.380 ;
        RECT 1318.020 63.370 1321.020 63.380 ;
        RECT 1498.020 63.370 1501.020 63.380 ;
        RECT 1678.020 63.370 1681.020 63.380 ;
        RECT 1858.020 63.370 1861.020 63.380 ;
        RECT 2038.020 63.370 2041.020 63.380 ;
        RECT 2218.020 63.370 2221.020 63.380 ;
        RECT 2398.020 63.370 2401.020 63.380 ;
        RECT 2578.020 63.370 2581.020 63.380 ;
        RECT 2758.020 63.370 2761.020 63.380 ;
        RECT 2954.200 63.370 2957.200 63.380 ;
        RECT -37.580 -29.220 -34.580 -29.210 ;
        RECT 58.020 -29.220 61.020 -29.210 ;
        RECT 238.020 -29.220 241.020 -29.210 ;
        RECT 418.020 -29.220 421.020 -29.210 ;
        RECT 598.020 -29.220 601.020 -29.210 ;
        RECT 778.020 -29.220 781.020 -29.210 ;
        RECT 958.020 -29.220 961.020 -29.210 ;
        RECT 1138.020 -29.220 1141.020 -29.210 ;
        RECT 1318.020 -29.220 1321.020 -29.210 ;
        RECT 1498.020 -29.220 1501.020 -29.210 ;
        RECT 1678.020 -29.220 1681.020 -29.210 ;
        RECT 1858.020 -29.220 1861.020 -29.210 ;
        RECT 2038.020 -29.220 2041.020 -29.210 ;
        RECT 2218.020 -29.220 2221.020 -29.210 ;
        RECT 2398.020 -29.220 2401.020 -29.210 ;
        RECT 2578.020 -29.220 2581.020 -29.210 ;
        RECT 2758.020 -29.220 2761.020 -29.210 ;
        RECT 2954.200 -29.220 2957.200 -29.210 ;
        RECT -37.580 -32.220 2957.200 -29.220 ;
        RECT -37.580 -32.230 -34.580 -32.220 ;
        RECT 58.020 -32.230 61.020 -32.220 ;
        RECT 238.020 -32.230 241.020 -32.220 ;
        RECT 418.020 -32.230 421.020 -32.220 ;
        RECT 598.020 -32.230 601.020 -32.220 ;
        RECT 778.020 -32.230 781.020 -32.220 ;
        RECT 958.020 -32.230 961.020 -32.220 ;
        RECT 1138.020 -32.230 1141.020 -32.220 ;
        RECT 1318.020 -32.230 1321.020 -32.220 ;
        RECT 1498.020 -32.230 1501.020 -32.220 ;
        RECT 1678.020 -32.230 1681.020 -32.220 ;
        RECT 1858.020 -32.230 1861.020 -32.220 ;
        RECT 2038.020 -32.230 2041.020 -32.220 ;
        RECT 2218.020 -32.230 2221.020 -32.220 ;
        RECT 2398.020 -32.230 2401.020 -32.220 ;
        RECT 2578.020 -32.230 2581.020 -32.220 ;
        RECT 2758.020 -32.230 2761.020 -32.220 ;
        RECT 2954.200 -32.230 2957.200 -32.220 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -42.180 -36.820 -39.180 3556.500 ;
        RECT 148.020 -36.820 151.020 3556.500 ;
        RECT 328.020 -36.820 331.020 3556.500 ;
        RECT 508.020 -36.820 511.020 3556.500 ;
        RECT 688.020 -36.820 691.020 3556.500 ;
        RECT 868.020 -36.820 871.020 3556.500 ;
        RECT 1048.020 -36.820 1051.020 3556.500 ;
        RECT 1228.020 -36.820 1231.020 3556.500 ;
        RECT 1408.020 -36.820 1411.020 3556.500 ;
        RECT 1588.020 -36.820 1591.020 3556.500 ;
        RECT 1768.020 -36.820 1771.020 3556.500 ;
        RECT 1948.020 -36.820 1951.020 3556.500 ;
        RECT 2128.020 -36.820 2131.020 3556.500 ;
        RECT 2308.020 -36.820 2311.020 3556.500 ;
        RECT 2488.020 -36.820 2491.020 3556.500 ;
        RECT 2668.020 -36.820 2671.020 3556.500 ;
        RECT 2848.020 -36.820 2851.020 3556.500 ;
        RECT 2958.800 -36.820 2961.800 3556.500 ;
      LAYER via4 ;
        RECT -41.270 3555.210 -40.090 3556.390 ;
        RECT -41.270 3553.610 -40.090 3554.790 ;
        RECT -41.270 3395.090 -40.090 3396.270 ;
        RECT -41.270 3393.490 -40.090 3394.670 ;
        RECT -41.270 3215.090 -40.090 3216.270 ;
        RECT -41.270 3213.490 -40.090 3214.670 ;
        RECT -41.270 3035.090 -40.090 3036.270 ;
        RECT -41.270 3033.490 -40.090 3034.670 ;
        RECT -41.270 2855.090 -40.090 2856.270 ;
        RECT -41.270 2853.490 -40.090 2854.670 ;
        RECT -41.270 2675.090 -40.090 2676.270 ;
        RECT -41.270 2673.490 -40.090 2674.670 ;
        RECT -41.270 2495.090 -40.090 2496.270 ;
        RECT -41.270 2493.490 -40.090 2494.670 ;
        RECT -41.270 2315.090 -40.090 2316.270 ;
        RECT -41.270 2313.490 -40.090 2314.670 ;
        RECT -41.270 2135.090 -40.090 2136.270 ;
        RECT -41.270 2133.490 -40.090 2134.670 ;
        RECT -41.270 1955.090 -40.090 1956.270 ;
        RECT -41.270 1953.490 -40.090 1954.670 ;
        RECT -41.270 1775.090 -40.090 1776.270 ;
        RECT -41.270 1773.490 -40.090 1774.670 ;
        RECT -41.270 1595.090 -40.090 1596.270 ;
        RECT -41.270 1593.490 -40.090 1594.670 ;
        RECT -41.270 1415.090 -40.090 1416.270 ;
        RECT -41.270 1413.490 -40.090 1414.670 ;
        RECT -41.270 1235.090 -40.090 1236.270 ;
        RECT -41.270 1233.490 -40.090 1234.670 ;
        RECT -41.270 1055.090 -40.090 1056.270 ;
        RECT -41.270 1053.490 -40.090 1054.670 ;
        RECT -41.270 875.090 -40.090 876.270 ;
        RECT -41.270 873.490 -40.090 874.670 ;
        RECT -41.270 695.090 -40.090 696.270 ;
        RECT -41.270 693.490 -40.090 694.670 ;
        RECT -41.270 515.090 -40.090 516.270 ;
        RECT -41.270 513.490 -40.090 514.670 ;
        RECT -41.270 335.090 -40.090 336.270 ;
        RECT -41.270 333.490 -40.090 334.670 ;
        RECT -41.270 155.090 -40.090 156.270 ;
        RECT -41.270 153.490 -40.090 154.670 ;
        RECT -41.270 -35.110 -40.090 -33.930 ;
        RECT -41.270 -36.710 -40.090 -35.530 ;
        RECT 148.930 3555.210 150.110 3556.390 ;
        RECT 148.930 3553.610 150.110 3554.790 ;
        RECT 148.930 3395.090 150.110 3396.270 ;
        RECT 148.930 3393.490 150.110 3394.670 ;
        RECT 148.930 3215.090 150.110 3216.270 ;
        RECT 148.930 3213.490 150.110 3214.670 ;
        RECT 148.930 3035.090 150.110 3036.270 ;
        RECT 148.930 3033.490 150.110 3034.670 ;
        RECT 148.930 2855.090 150.110 2856.270 ;
        RECT 148.930 2853.490 150.110 2854.670 ;
        RECT 148.930 2675.090 150.110 2676.270 ;
        RECT 148.930 2673.490 150.110 2674.670 ;
        RECT 148.930 2495.090 150.110 2496.270 ;
        RECT 148.930 2493.490 150.110 2494.670 ;
        RECT 148.930 2315.090 150.110 2316.270 ;
        RECT 148.930 2313.490 150.110 2314.670 ;
        RECT 148.930 2135.090 150.110 2136.270 ;
        RECT 148.930 2133.490 150.110 2134.670 ;
        RECT 148.930 1955.090 150.110 1956.270 ;
        RECT 148.930 1953.490 150.110 1954.670 ;
        RECT 148.930 1775.090 150.110 1776.270 ;
        RECT 148.930 1773.490 150.110 1774.670 ;
        RECT 148.930 1595.090 150.110 1596.270 ;
        RECT 148.930 1593.490 150.110 1594.670 ;
        RECT 148.930 1415.090 150.110 1416.270 ;
        RECT 148.930 1413.490 150.110 1414.670 ;
        RECT 148.930 1235.090 150.110 1236.270 ;
        RECT 148.930 1233.490 150.110 1234.670 ;
        RECT 148.930 1055.090 150.110 1056.270 ;
        RECT 148.930 1053.490 150.110 1054.670 ;
        RECT 148.930 875.090 150.110 876.270 ;
        RECT 148.930 873.490 150.110 874.670 ;
        RECT 148.930 695.090 150.110 696.270 ;
        RECT 148.930 693.490 150.110 694.670 ;
        RECT 148.930 515.090 150.110 516.270 ;
        RECT 148.930 513.490 150.110 514.670 ;
        RECT 148.930 335.090 150.110 336.270 ;
        RECT 148.930 333.490 150.110 334.670 ;
        RECT 148.930 155.090 150.110 156.270 ;
        RECT 148.930 153.490 150.110 154.670 ;
        RECT 148.930 -35.110 150.110 -33.930 ;
        RECT 148.930 -36.710 150.110 -35.530 ;
        RECT 328.930 3555.210 330.110 3556.390 ;
        RECT 328.930 3553.610 330.110 3554.790 ;
        RECT 328.930 3395.090 330.110 3396.270 ;
        RECT 328.930 3393.490 330.110 3394.670 ;
        RECT 328.930 3215.090 330.110 3216.270 ;
        RECT 328.930 3213.490 330.110 3214.670 ;
        RECT 328.930 3035.090 330.110 3036.270 ;
        RECT 328.930 3033.490 330.110 3034.670 ;
        RECT 328.930 2855.090 330.110 2856.270 ;
        RECT 328.930 2853.490 330.110 2854.670 ;
        RECT 328.930 2675.090 330.110 2676.270 ;
        RECT 328.930 2673.490 330.110 2674.670 ;
        RECT 328.930 2495.090 330.110 2496.270 ;
        RECT 328.930 2493.490 330.110 2494.670 ;
        RECT 328.930 2315.090 330.110 2316.270 ;
        RECT 328.930 2313.490 330.110 2314.670 ;
        RECT 328.930 2135.090 330.110 2136.270 ;
        RECT 328.930 2133.490 330.110 2134.670 ;
        RECT 328.930 1955.090 330.110 1956.270 ;
        RECT 328.930 1953.490 330.110 1954.670 ;
        RECT 328.930 1775.090 330.110 1776.270 ;
        RECT 328.930 1773.490 330.110 1774.670 ;
        RECT 328.930 1595.090 330.110 1596.270 ;
        RECT 328.930 1593.490 330.110 1594.670 ;
        RECT 328.930 1415.090 330.110 1416.270 ;
        RECT 328.930 1413.490 330.110 1414.670 ;
        RECT 328.930 1235.090 330.110 1236.270 ;
        RECT 328.930 1233.490 330.110 1234.670 ;
        RECT 328.930 1055.090 330.110 1056.270 ;
        RECT 328.930 1053.490 330.110 1054.670 ;
        RECT 328.930 875.090 330.110 876.270 ;
        RECT 328.930 873.490 330.110 874.670 ;
        RECT 328.930 695.090 330.110 696.270 ;
        RECT 328.930 693.490 330.110 694.670 ;
        RECT 328.930 515.090 330.110 516.270 ;
        RECT 328.930 513.490 330.110 514.670 ;
        RECT 328.930 335.090 330.110 336.270 ;
        RECT 328.930 333.490 330.110 334.670 ;
        RECT 328.930 155.090 330.110 156.270 ;
        RECT 328.930 153.490 330.110 154.670 ;
        RECT 328.930 -35.110 330.110 -33.930 ;
        RECT 328.930 -36.710 330.110 -35.530 ;
        RECT 508.930 3555.210 510.110 3556.390 ;
        RECT 508.930 3553.610 510.110 3554.790 ;
        RECT 508.930 3395.090 510.110 3396.270 ;
        RECT 508.930 3393.490 510.110 3394.670 ;
        RECT 508.930 3215.090 510.110 3216.270 ;
        RECT 508.930 3213.490 510.110 3214.670 ;
        RECT 508.930 3035.090 510.110 3036.270 ;
        RECT 508.930 3033.490 510.110 3034.670 ;
        RECT 508.930 2855.090 510.110 2856.270 ;
        RECT 508.930 2853.490 510.110 2854.670 ;
        RECT 508.930 2675.090 510.110 2676.270 ;
        RECT 508.930 2673.490 510.110 2674.670 ;
        RECT 508.930 2495.090 510.110 2496.270 ;
        RECT 508.930 2493.490 510.110 2494.670 ;
        RECT 508.930 2315.090 510.110 2316.270 ;
        RECT 508.930 2313.490 510.110 2314.670 ;
        RECT 508.930 2135.090 510.110 2136.270 ;
        RECT 508.930 2133.490 510.110 2134.670 ;
        RECT 508.930 1955.090 510.110 1956.270 ;
        RECT 508.930 1953.490 510.110 1954.670 ;
        RECT 508.930 1775.090 510.110 1776.270 ;
        RECT 508.930 1773.490 510.110 1774.670 ;
        RECT 508.930 1595.090 510.110 1596.270 ;
        RECT 508.930 1593.490 510.110 1594.670 ;
        RECT 508.930 1415.090 510.110 1416.270 ;
        RECT 508.930 1413.490 510.110 1414.670 ;
        RECT 508.930 1235.090 510.110 1236.270 ;
        RECT 508.930 1233.490 510.110 1234.670 ;
        RECT 508.930 1055.090 510.110 1056.270 ;
        RECT 508.930 1053.490 510.110 1054.670 ;
        RECT 508.930 875.090 510.110 876.270 ;
        RECT 508.930 873.490 510.110 874.670 ;
        RECT 508.930 695.090 510.110 696.270 ;
        RECT 508.930 693.490 510.110 694.670 ;
        RECT 508.930 515.090 510.110 516.270 ;
        RECT 508.930 513.490 510.110 514.670 ;
        RECT 508.930 335.090 510.110 336.270 ;
        RECT 508.930 333.490 510.110 334.670 ;
        RECT 508.930 155.090 510.110 156.270 ;
        RECT 508.930 153.490 510.110 154.670 ;
        RECT 508.930 -35.110 510.110 -33.930 ;
        RECT 508.930 -36.710 510.110 -35.530 ;
        RECT 688.930 3555.210 690.110 3556.390 ;
        RECT 688.930 3553.610 690.110 3554.790 ;
        RECT 688.930 3395.090 690.110 3396.270 ;
        RECT 688.930 3393.490 690.110 3394.670 ;
        RECT 688.930 3215.090 690.110 3216.270 ;
        RECT 688.930 3213.490 690.110 3214.670 ;
        RECT 688.930 3035.090 690.110 3036.270 ;
        RECT 688.930 3033.490 690.110 3034.670 ;
        RECT 688.930 2855.090 690.110 2856.270 ;
        RECT 688.930 2853.490 690.110 2854.670 ;
        RECT 688.930 2675.090 690.110 2676.270 ;
        RECT 688.930 2673.490 690.110 2674.670 ;
        RECT 688.930 2495.090 690.110 2496.270 ;
        RECT 688.930 2493.490 690.110 2494.670 ;
        RECT 688.930 2315.090 690.110 2316.270 ;
        RECT 688.930 2313.490 690.110 2314.670 ;
        RECT 688.930 2135.090 690.110 2136.270 ;
        RECT 688.930 2133.490 690.110 2134.670 ;
        RECT 688.930 1955.090 690.110 1956.270 ;
        RECT 688.930 1953.490 690.110 1954.670 ;
        RECT 688.930 1775.090 690.110 1776.270 ;
        RECT 688.930 1773.490 690.110 1774.670 ;
        RECT 688.930 1595.090 690.110 1596.270 ;
        RECT 688.930 1593.490 690.110 1594.670 ;
        RECT 688.930 1415.090 690.110 1416.270 ;
        RECT 688.930 1413.490 690.110 1414.670 ;
        RECT 688.930 1235.090 690.110 1236.270 ;
        RECT 688.930 1233.490 690.110 1234.670 ;
        RECT 688.930 1055.090 690.110 1056.270 ;
        RECT 688.930 1053.490 690.110 1054.670 ;
        RECT 688.930 875.090 690.110 876.270 ;
        RECT 688.930 873.490 690.110 874.670 ;
        RECT 688.930 695.090 690.110 696.270 ;
        RECT 688.930 693.490 690.110 694.670 ;
        RECT 688.930 515.090 690.110 516.270 ;
        RECT 688.930 513.490 690.110 514.670 ;
        RECT 688.930 335.090 690.110 336.270 ;
        RECT 688.930 333.490 690.110 334.670 ;
        RECT 688.930 155.090 690.110 156.270 ;
        RECT 688.930 153.490 690.110 154.670 ;
        RECT 688.930 -35.110 690.110 -33.930 ;
        RECT 688.930 -36.710 690.110 -35.530 ;
        RECT 868.930 3555.210 870.110 3556.390 ;
        RECT 868.930 3553.610 870.110 3554.790 ;
        RECT 868.930 3395.090 870.110 3396.270 ;
        RECT 868.930 3393.490 870.110 3394.670 ;
        RECT 868.930 3215.090 870.110 3216.270 ;
        RECT 868.930 3213.490 870.110 3214.670 ;
        RECT 868.930 3035.090 870.110 3036.270 ;
        RECT 868.930 3033.490 870.110 3034.670 ;
        RECT 868.930 2855.090 870.110 2856.270 ;
        RECT 868.930 2853.490 870.110 2854.670 ;
        RECT 868.930 2675.090 870.110 2676.270 ;
        RECT 868.930 2673.490 870.110 2674.670 ;
        RECT 868.930 2495.090 870.110 2496.270 ;
        RECT 868.930 2493.490 870.110 2494.670 ;
        RECT 868.930 2315.090 870.110 2316.270 ;
        RECT 868.930 2313.490 870.110 2314.670 ;
        RECT 868.930 2135.090 870.110 2136.270 ;
        RECT 868.930 2133.490 870.110 2134.670 ;
        RECT 868.930 1955.090 870.110 1956.270 ;
        RECT 868.930 1953.490 870.110 1954.670 ;
        RECT 868.930 1775.090 870.110 1776.270 ;
        RECT 868.930 1773.490 870.110 1774.670 ;
        RECT 868.930 1595.090 870.110 1596.270 ;
        RECT 868.930 1593.490 870.110 1594.670 ;
        RECT 868.930 1415.090 870.110 1416.270 ;
        RECT 868.930 1413.490 870.110 1414.670 ;
        RECT 868.930 1235.090 870.110 1236.270 ;
        RECT 868.930 1233.490 870.110 1234.670 ;
        RECT 868.930 1055.090 870.110 1056.270 ;
        RECT 868.930 1053.490 870.110 1054.670 ;
        RECT 868.930 875.090 870.110 876.270 ;
        RECT 868.930 873.490 870.110 874.670 ;
        RECT 868.930 695.090 870.110 696.270 ;
        RECT 868.930 693.490 870.110 694.670 ;
        RECT 868.930 515.090 870.110 516.270 ;
        RECT 868.930 513.490 870.110 514.670 ;
        RECT 868.930 335.090 870.110 336.270 ;
        RECT 868.930 333.490 870.110 334.670 ;
        RECT 868.930 155.090 870.110 156.270 ;
        RECT 868.930 153.490 870.110 154.670 ;
        RECT 868.930 -35.110 870.110 -33.930 ;
        RECT 868.930 -36.710 870.110 -35.530 ;
        RECT 1048.930 3555.210 1050.110 3556.390 ;
        RECT 1048.930 3553.610 1050.110 3554.790 ;
        RECT 1048.930 3395.090 1050.110 3396.270 ;
        RECT 1048.930 3393.490 1050.110 3394.670 ;
        RECT 1048.930 3215.090 1050.110 3216.270 ;
        RECT 1048.930 3213.490 1050.110 3214.670 ;
        RECT 1048.930 3035.090 1050.110 3036.270 ;
        RECT 1048.930 3033.490 1050.110 3034.670 ;
        RECT 1048.930 2855.090 1050.110 2856.270 ;
        RECT 1048.930 2853.490 1050.110 2854.670 ;
        RECT 1048.930 2675.090 1050.110 2676.270 ;
        RECT 1048.930 2673.490 1050.110 2674.670 ;
        RECT 1048.930 2495.090 1050.110 2496.270 ;
        RECT 1048.930 2493.490 1050.110 2494.670 ;
        RECT 1048.930 2315.090 1050.110 2316.270 ;
        RECT 1048.930 2313.490 1050.110 2314.670 ;
        RECT 1048.930 2135.090 1050.110 2136.270 ;
        RECT 1048.930 2133.490 1050.110 2134.670 ;
        RECT 1048.930 1955.090 1050.110 1956.270 ;
        RECT 1048.930 1953.490 1050.110 1954.670 ;
        RECT 1048.930 1775.090 1050.110 1776.270 ;
        RECT 1048.930 1773.490 1050.110 1774.670 ;
        RECT 1048.930 1595.090 1050.110 1596.270 ;
        RECT 1048.930 1593.490 1050.110 1594.670 ;
        RECT 1048.930 1415.090 1050.110 1416.270 ;
        RECT 1048.930 1413.490 1050.110 1414.670 ;
        RECT 1048.930 1235.090 1050.110 1236.270 ;
        RECT 1048.930 1233.490 1050.110 1234.670 ;
        RECT 1048.930 1055.090 1050.110 1056.270 ;
        RECT 1048.930 1053.490 1050.110 1054.670 ;
        RECT 1048.930 875.090 1050.110 876.270 ;
        RECT 1048.930 873.490 1050.110 874.670 ;
        RECT 1048.930 695.090 1050.110 696.270 ;
        RECT 1048.930 693.490 1050.110 694.670 ;
        RECT 1048.930 515.090 1050.110 516.270 ;
        RECT 1048.930 513.490 1050.110 514.670 ;
        RECT 1048.930 335.090 1050.110 336.270 ;
        RECT 1048.930 333.490 1050.110 334.670 ;
        RECT 1048.930 155.090 1050.110 156.270 ;
        RECT 1048.930 153.490 1050.110 154.670 ;
        RECT 1048.930 -35.110 1050.110 -33.930 ;
        RECT 1048.930 -36.710 1050.110 -35.530 ;
        RECT 1228.930 3555.210 1230.110 3556.390 ;
        RECT 1228.930 3553.610 1230.110 3554.790 ;
        RECT 1228.930 3395.090 1230.110 3396.270 ;
        RECT 1228.930 3393.490 1230.110 3394.670 ;
        RECT 1228.930 3215.090 1230.110 3216.270 ;
        RECT 1228.930 3213.490 1230.110 3214.670 ;
        RECT 1228.930 3035.090 1230.110 3036.270 ;
        RECT 1228.930 3033.490 1230.110 3034.670 ;
        RECT 1228.930 2855.090 1230.110 2856.270 ;
        RECT 1228.930 2853.490 1230.110 2854.670 ;
        RECT 1228.930 2675.090 1230.110 2676.270 ;
        RECT 1228.930 2673.490 1230.110 2674.670 ;
        RECT 1228.930 2495.090 1230.110 2496.270 ;
        RECT 1228.930 2493.490 1230.110 2494.670 ;
        RECT 1228.930 2315.090 1230.110 2316.270 ;
        RECT 1228.930 2313.490 1230.110 2314.670 ;
        RECT 1228.930 2135.090 1230.110 2136.270 ;
        RECT 1228.930 2133.490 1230.110 2134.670 ;
        RECT 1228.930 1955.090 1230.110 1956.270 ;
        RECT 1228.930 1953.490 1230.110 1954.670 ;
        RECT 1228.930 1775.090 1230.110 1776.270 ;
        RECT 1228.930 1773.490 1230.110 1774.670 ;
        RECT 1228.930 1595.090 1230.110 1596.270 ;
        RECT 1228.930 1593.490 1230.110 1594.670 ;
        RECT 1228.930 1415.090 1230.110 1416.270 ;
        RECT 1228.930 1413.490 1230.110 1414.670 ;
        RECT 1228.930 1235.090 1230.110 1236.270 ;
        RECT 1228.930 1233.490 1230.110 1234.670 ;
        RECT 1228.930 1055.090 1230.110 1056.270 ;
        RECT 1228.930 1053.490 1230.110 1054.670 ;
        RECT 1228.930 875.090 1230.110 876.270 ;
        RECT 1228.930 873.490 1230.110 874.670 ;
        RECT 1228.930 695.090 1230.110 696.270 ;
        RECT 1228.930 693.490 1230.110 694.670 ;
        RECT 1228.930 515.090 1230.110 516.270 ;
        RECT 1228.930 513.490 1230.110 514.670 ;
        RECT 1228.930 335.090 1230.110 336.270 ;
        RECT 1228.930 333.490 1230.110 334.670 ;
        RECT 1228.930 155.090 1230.110 156.270 ;
        RECT 1228.930 153.490 1230.110 154.670 ;
        RECT 1228.930 -35.110 1230.110 -33.930 ;
        RECT 1228.930 -36.710 1230.110 -35.530 ;
        RECT 1408.930 3555.210 1410.110 3556.390 ;
        RECT 1408.930 3553.610 1410.110 3554.790 ;
        RECT 1408.930 3395.090 1410.110 3396.270 ;
        RECT 1408.930 3393.490 1410.110 3394.670 ;
        RECT 1408.930 3215.090 1410.110 3216.270 ;
        RECT 1408.930 3213.490 1410.110 3214.670 ;
        RECT 1408.930 3035.090 1410.110 3036.270 ;
        RECT 1408.930 3033.490 1410.110 3034.670 ;
        RECT 1408.930 2855.090 1410.110 2856.270 ;
        RECT 1408.930 2853.490 1410.110 2854.670 ;
        RECT 1408.930 2675.090 1410.110 2676.270 ;
        RECT 1408.930 2673.490 1410.110 2674.670 ;
        RECT 1408.930 2495.090 1410.110 2496.270 ;
        RECT 1408.930 2493.490 1410.110 2494.670 ;
        RECT 1408.930 2315.090 1410.110 2316.270 ;
        RECT 1408.930 2313.490 1410.110 2314.670 ;
        RECT 1408.930 2135.090 1410.110 2136.270 ;
        RECT 1408.930 2133.490 1410.110 2134.670 ;
        RECT 1408.930 1955.090 1410.110 1956.270 ;
        RECT 1408.930 1953.490 1410.110 1954.670 ;
        RECT 1408.930 1775.090 1410.110 1776.270 ;
        RECT 1408.930 1773.490 1410.110 1774.670 ;
        RECT 1408.930 1595.090 1410.110 1596.270 ;
        RECT 1408.930 1593.490 1410.110 1594.670 ;
        RECT 1408.930 1415.090 1410.110 1416.270 ;
        RECT 1408.930 1413.490 1410.110 1414.670 ;
        RECT 1408.930 1235.090 1410.110 1236.270 ;
        RECT 1408.930 1233.490 1410.110 1234.670 ;
        RECT 1408.930 1055.090 1410.110 1056.270 ;
        RECT 1408.930 1053.490 1410.110 1054.670 ;
        RECT 1408.930 875.090 1410.110 876.270 ;
        RECT 1408.930 873.490 1410.110 874.670 ;
        RECT 1408.930 695.090 1410.110 696.270 ;
        RECT 1408.930 693.490 1410.110 694.670 ;
        RECT 1408.930 515.090 1410.110 516.270 ;
        RECT 1408.930 513.490 1410.110 514.670 ;
        RECT 1408.930 335.090 1410.110 336.270 ;
        RECT 1408.930 333.490 1410.110 334.670 ;
        RECT 1408.930 155.090 1410.110 156.270 ;
        RECT 1408.930 153.490 1410.110 154.670 ;
        RECT 1408.930 -35.110 1410.110 -33.930 ;
        RECT 1408.930 -36.710 1410.110 -35.530 ;
        RECT 1588.930 3555.210 1590.110 3556.390 ;
        RECT 1588.930 3553.610 1590.110 3554.790 ;
        RECT 1588.930 3395.090 1590.110 3396.270 ;
        RECT 1588.930 3393.490 1590.110 3394.670 ;
        RECT 1588.930 3215.090 1590.110 3216.270 ;
        RECT 1588.930 3213.490 1590.110 3214.670 ;
        RECT 1588.930 3035.090 1590.110 3036.270 ;
        RECT 1588.930 3033.490 1590.110 3034.670 ;
        RECT 1588.930 2855.090 1590.110 2856.270 ;
        RECT 1588.930 2853.490 1590.110 2854.670 ;
        RECT 1588.930 2675.090 1590.110 2676.270 ;
        RECT 1588.930 2673.490 1590.110 2674.670 ;
        RECT 1588.930 2495.090 1590.110 2496.270 ;
        RECT 1588.930 2493.490 1590.110 2494.670 ;
        RECT 1588.930 2315.090 1590.110 2316.270 ;
        RECT 1588.930 2313.490 1590.110 2314.670 ;
        RECT 1588.930 2135.090 1590.110 2136.270 ;
        RECT 1588.930 2133.490 1590.110 2134.670 ;
        RECT 1588.930 1955.090 1590.110 1956.270 ;
        RECT 1588.930 1953.490 1590.110 1954.670 ;
        RECT 1588.930 1775.090 1590.110 1776.270 ;
        RECT 1588.930 1773.490 1590.110 1774.670 ;
        RECT 1588.930 1595.090 1590.110 1596.270 ;
        RECT 1588.930 1593.490 1590.110 1594.670 ;
        RECT 1588.930 1415.090 1590.110 1416.270 ;
        RECT 1588.930 1413.490 1590.110 1414.670 ;
        RECT 1588.930 1235.090 1590.110 1236.270 ;
        RECT 1588.930 1233.490 1590.110 1234.670 ;
        RECT 1588.930 1055.090 1590.110 1056.270 ;
        RECT 1588.930 1053.490 1590.110 1054.670 ;
        RECT 1588.930 875.090 1590.110 876.270 ;
        RECT 1588.930 873.490 1590.110 874.670 ;
        RECT 1588.930 695.090 1590.110 696.270 ;
        RECT 1588.930 693.490 1590.110 694.670 ;
        RECT 1588.930 515.090 1590.110 516.270 ;
        RECT 1588.930 513.490 1590.110 514.670 ;
        RECT 1588.930 335.090 1590.110 336.270 ;
        RECT 1588.930 333.490 1590.110 334.670 ;
        RECT 1588.930 155.090 1590.110 156.270 ;
        RECT 1588.930 153.490 1590.110 154.670 ;
        RECT 1588.930 -35.110 1590.110 -33.930 ;
        RECT 1588.930 -36.710 1590.110 -35.530 ;
        RECT 1768.930 3555.210 1770.110 3556.390 ;
        RECT 1768.930 3553.610 1770.110 3554.790 ;
        RECT 1768.930 3395.090 1770.110 3396.270 ;
        RECT 1768.930 3393.490 1770.110 3394.670 ;
        RECT 1768.930 3215.090 1770.110 3216.270 ;
        RECT 1768.930 3213.490 1770.110 3214.670 ;
        RECT 1768.930 3035.090 1770.110 3036.270 ;
        RECT 1768.930 3033.490 1770.110 3034.670 ;
        RECT 1768.930 2855.090 1770.110 2856.270 ;
        RECT 1768.930 2853.490 1770.110 2854.670 ;
        RECT 1768.930 2675.090 1770.110 2676.270 ;
        RECT 1768.930 2673.490 1770.110 2674.670 ;
        RECT 1768.930 2495.090 1770.110 2496.270 ;
        RECT 1768.930 2493.490 1770.110 2494.670 ;
        RECT 1768.930 2315.090 1770.110 2316.270 ;
        RECT 1768.930 2313.490 1770.110 2314.670 ;
        RECT 1768.930 2135.090 1770.110 2136.270 ;
        RECT 1768.930 2133.490 1770.110 2134.670 ;
        RECT 1768.930 1955.090 1770.110 1956.270 ;
        RECT 1768.930 1953.490 1770.110 1954.670 ;
        RECT 1768.930 1775.090 1770.110 1776.270 ;
        RECT 1768.930 1773.490 1770.110 1774.670 ;
        RECT 1768.930 1595.090 1770.110 1596.270 ;
        RECT 1768.930 1593.490 1770.110 1594.670 ;
        RECT 1768.930 1415.090 1770.110 1416.270 ;
        RECT 1768.930 1413.490 1770.110 1414.670 ;
        RECT 1768.930 1235.090 1770.110 1236.270 ;
        RECT 1768.930 1233.490 1770.110 1234.670 ;
        RECT 1768.930 1055.090 1770.110 1056.270 ;
        RECT 1768.930 1053.490 1770.110 1054.670 ;
        RECT 1768.930 875.090 1770.110 876.270 ;
        RECT 1768.930 873.490 1770.110 874.670 ;
        RECT 1768.930 695.090 1770.110 696.270 ;
        RECT 1768.930 693.490 1770.110 694.670 ;
        RECT 1768.930 515.090 1770.110 516.270 ;
        RECT 1768.930 513.490 1770.110 514.670 ;
        RECT 1768.930 335.090 1770.110 336.270 ;
        RECT 1768.930 333.490 1770.110 334.670 ;
        RECT 1768.930 155.090 1770.110 156.270 ;
        RECT 1768.930 153.490 1770.110 154.670 ;
        RECT 1768.930 -35.110 1770.110 -33.930 ;
        RECT 1768.930 -36.710 1770.110 -35.530 ;
        RECT 1948.930 3555.210 1950.110 3556.390 ;
        RECT 1948.930 3553.610 1950.110 3554.790 ;
        RECT 1948.930 3395.090 1950.110 3396.270 ;
        RECT 1948.930 3393.490 1950.110 3394.670 ;
        RECT 1948.930 3215.090 1950.110 3216.270 ;
        RECT 1948.930 3213.490 1950.110 3214.670 ;
        RECT 1948.930 3035.090 1950.110 3036.270 ;
        RECT 1948.930 3033.490 1950.110 3034.670 ;
        RECT 1948.930 2855.090 1950.110 2856.270 ;
        RECT 1948.930 2853.490 1950.110 2854.670 ;
        RECT 1948.930 2675.090 1950.110 2676.270 ;
        RECT 1948.930 2673.490 1950.110 2674.670 ;
        RECT 1948.930 2495.090 1950.110 2496.270 ;
        RECT 1948.930 2493.490 1950.110 2494.670 ;
        RECT 1948.930 2315.090 1950.110 2316.270 ;
        RECT 1948.930 2313.490 1950.110 2314.670 ;
        RECT 1948.930 2135.090 1950.110 2136.270 ;
        RECT 1948.930 2133.490 1950.110 2134.670 ;
        RECT 1948.930 1955.090 1950.110 1956.270 ;
        RECT 1948.930 1953.490 1950.110 1954.670 ;
        RECT 1948.930 1775.090 1950.110 1776.270 ;
        RECT 1948.930 1773.490 1950.110 1774.670 ;
        RECT 1948.930 1595.090 1950.110 1596.270 ;
        RECT 1948.930 1593.490 1950.110 1594.670 ;
        RECT 1948.930 1415.090 1950.110 1416.270 ;
        RECT 1948.930 1413.490 1950.110 1414.670 ;
        RECT 1948.930 1235.090 1950.110 1236.270 ;
        RECT 1948.930 1233.490 1950.110 1234.670 ;
        RECT 1948.930 1055.090 1950.110 1056.270 ;
        RECT 1948.930 1053.490 1950.110 1054.670 ;
        RECT 1948.930 875.090 1950.110 876.270 ;
        RECT 1948.930 873.490 1950.110 874.670 ;
        RECT 1948.930 695.090 1950.110 696.270 ;
        RECT 1948.930 693.490 1950.110 694.670 ;
        RECT 1948.930 515.090 1950.110 516.270 ;
        RECT 1948.930 513.490 1950.110 514.670 ;
        RECT 1948.930 335.090 1950.110 336.270 ;
        RECT 1948.930 333.490 1950.110 334.670 ;
        RECT 1948.930 155.090 1950.110 156.270 ;
        RECT 1948.930 153.490 1950.110 154.670 ;
        RECT 1948.930 -35.110 1950.110 -33.930 ;
        RECT 1948.930 -36.710 1950.110 -35.530 ;
        RECT 2128.930 3555.210 2130.110 3556.390 ;
        RECT 2128.930 3553.610 2130.110 3554.790 ;
        RECT 2128.930 3395.090 2130.110 3396.270 ;
        RECT 2128.930 3393.490 2130.110 3394.670 ;
        RECT 2128.930 3215.090 2130.110 3216.270 ;
        RECT 2128.930 3213.490 2130.110 3214.670 ;
        RECT 2128.930 3035.090 2130.110 3036.270 ;
        RECT 2128.930 3033.490 2130.110 3034.670 ;
        RECT 2128.930 2855.090 2130.110 2856.270 ;
        RECT 2128.930 2853.490 2130.110 2854.670 ;
        RECT 2128.930 2675.090 2130.110 2676.270 ;
        RECT 2128.930 2673.490 2130.110 2674.670 ;
        RECT 2128.930 2495.090 2130.110 2496.270 ;
        RECT 2128.930 2493.490 2130.110 2494.670 ;
        RECT 2128.930 2315.090 2130.110 2316.270 ;
        RECT 2128.930 2313.490 2130.110 2314.670 ;
        RECT 2128.930 2135.090 2130.110 2136.270 ;
        RECT 2128.930 2133.490 2130.110 2134.670 ;
        RECT 2128.930 1955.090 2130.110 1956.270 ;
        RECT 2128.930 1953.490 2130.110 1954.670 ;
        RECT 2128.930 1775.090 2130.110 1776.270 ;
        RECT 2128.930 1773.490 2130.110 1774.670 ;
        RECT 2128.930 1595.090 2130.110 1596.270 ;
        RECT 2128.930 1593.490 2130.110 1594.670 ;
        RECT 2128.930 1415.090 2130.110 1416.270 ;
        RECT 2128.930 1413.490 2130.110 1414.670 ;
        RECT 2128.930 1235.090 2130.110 1236.270 ;
        RECT 2128.930 1233.490 2130.110 1234.670 ;
        RECT 2128.930 1055.090 2130.110 1056.270 ;
        RECT 2128.930 1053.490 2130.110 1054.670 ;
        RECT 2128.930 875.090 2130.110 876.270 ;
        RECT 2128.930 873.490 2130.110 874.670 ;
        RECT 2128.930 695.090 2130.110 696.270 ;
        RECT 2128.930 693.490 2130.110 694.670 ;
        RECT 2128.930 515.090 2130.110 516.270 ;
        RECT 2128.930 513.490 2130.110 514.670 ;
        RECT 2128.930 335.090 2130.110 336.270 ;
        RECT 2128.930 333.490 2130.110 334.670 ;
        RECT 2128.930 155.090 2130.110 156.270 ;
        RECT 2128.930 153.490 2130.110 154.670 ;
        RECT 2128.930 -35.110 2130.110 -33.930 ;
        RECT 2128.930 -36.710 2130.110 -35.530 ;
        RECT 2308.930 3555.210 2310.110 3556.390 ;
        RECT 2308.930 3553.610 2310.110 3554.790 ;
        RECT 2308.930 3395.090 2310.110 3396.270 ;
        RECT 2308.930 3393.490 2310.110 3394.670 ;
        RECT 2308.930 3215.090 2310.110 3216.270 ;
        RECT 2308.930 3213.490 2310.110 3214.670 ;
        RECT 2308.930 3035.090 2310.110 3036.270 ;
        RECT 2308.930 3033.490 2310.110 3034.670 ;
        RECT 2308.930 2855.090 2310.110 2856.270 ;
        RECT 2308.930 2853.490 2310.110 2854.670 ;
        RECT 2308.930 2675.090 2310.110 2676.270 ;
        RECT 2308.930 2673.490 2310.110 2674.670 ;
        RECT 2308.930 2495.090 2310.110 2496.270 ;
        RECT 2308.930 2493.490 2310.110 2494.670 ;
        RECT 2308.930 2315.090 2310.110 2316.270 ;
        RECT 2308.930 2313.490 2310.110 2314.670 ;
        RECT 2308.930 2135.090 2310.110 2136.270 ;
        RECT 2308.930 2133.490 2310.110 2134.670 ;
        RECT 2308.930 1955.090 2310.110 1956.270 ;
        RECT 2308.930 1953.490 2310.110 1954.670 ;
        RECT 2308.930 1775.090 2310.110 1776.270 ;
        RECT 2308.930 1773.490 2310.110 1774.670 ;
        RECT 2308.930 1595.090 2310.110 1596.270 ;
        RECT 2308.930 1593.490 2310.110 1594.670 ;
        RECT 2308.930 1415.090 2310.110 1416.270 ;
        RECT 2308.930 1413.490 2310.110 1414.670 ;
        RECT 2308.930 1235.090 2310.110 1236.270 ;
        RECT 2308.930 1233.490 2310.110 1234.670 ;
        RECT 2308.930 1055.090 2310.110 1056.270 ;
        RECT 2308.930 1053.490 2310.110 1054.670 ;
        RECT 2308.930 875.090 2310.110 876.270 ;
        RECT 2308.930 873.490 2310.110 874.670 ;
        RECT 2308.930 695.090 2310.110 696.270 ;
        RECT 2308.930 693.490 2310.110 694.670 ;
        RECT 2308.930 515.090 2310.110 516.270 ;
        RECT 2308.930 513.490 2310.110 514.670 ;
        RECT 2308.930 335.090 2310.110 336.270 ;
        RECT 2308.930 333.490 2310.110 334.670 ;
        RECT 2308.930 155.090 2310.110 156.270 ;
        RECT 2308.930 153.490 2310.110 154.670 ;
        RECT 2308.930 -35.110 2310.110 -33.930 ;
        RECT 2308.930 -36.710 2310.110 -35.530 ;
        RECT 2488.930 3555.210 2490.110 3556.390 ;
        RECT 2488.930 3553.610 2490.110 3554.790 ;
        RECT 2488.930 3395.090 2490.110 3396.270 ;
        RECT 2488.930 3393.490 2490.110 3394.670 ;
        RECT 2488.930 3215.090 2490.110 3216.270 ;
        RECT 2488.930 3213.490 2490.110 3214.670 ;
        RECT 2488.930 3035.090 2490.110 3036.270 ;
        RECT 2488.930 3033.490 2490.110 3034.670 ;
        RECT 2488.930 2855.090 2490.110 2856.270 ;
        RECT 2488.930 2853.490 2490.110 2854.670 ;
        RECT 2488.930 2675.090 2490.110 2676.270 ;
        RECT 2488.930 2673.490 2490.110 2674.670 ;
        RECT 2488.930 2495.090 2490.110 2496.270 ;
        RECT 2488.930 2493.490 2490.110 2494.670 ;
        RECT 2488.930 2315.090 2490.110 2316.270 ;
        RECT 2488.930 2313.490 2490.110 2314.670 ;
        RECT 2488.930 2135.090 2490.110 2136.270 ;
        RECT 2488.930 2133.490 2490.110 2134.670 ;
        RECT 2488.930 1955.090 2490.110 1956.270 ;
        RECT 2488.930 1953.490 2490.110 1954.670 ;
        RECT 2488.930 1775.090 2490.110 1776.270 ;
        RECT 2488.930 1773.490 2490.110 1774.670 ;
        RECT 2488.930 1595.090 2490.110 1596.270 ;
        RECT 2488.930 1593.490 2490.110 1594.670 ;
        RECT 2488.930 1415.090 2490.110 1416.270 ;
        RECT 2488.930 1413.490 2490.110 1414.670 ;
        RECT 2488.930 1235.090 2490.110 1236.270 ;
        RECT 2488.930 1233.490 2490.110 1234.670 ;
        RECT 2488.930 1055.090 2490.110 1056.270 ;
        RECT 2488.930 1053.490 2490.110 1054.670 ;
        RECT 2488.930 875.090 2490.110 876.270 ;
        RECT 2488.930 873.490 2490.110 874.670 ;
        RECT 2488.930 695.090 2490.110 696.270 ;
        RECT 2488.930 693.490 2490.110 694.670 ;
        RECT 2488.930 515.090 2490.110 516.270 ;
        RECT 2488.930 513.490 2490.110 514.670 ;
        RECT 2488.930 335.090 2490.110 336.270 ;
        RECT 2488.930 333.490 2490.110 334.670 ;
        RECT 2488.930 155.090 2490.110 156.270 ;
        RECT 2488.930 153.490 2490.110 154.670 ;
        RECT 2488.930 -35.110 2490.110 -33.930 ;
        RECT 2488.930 -36.710 2490.110 -35.530 ;
        RECT 2668.930 3555.210 2670.110 3556.390 ;
        RECT 2668.930 3553.610 2670.110 3554.790 ;
        RECT 2668.930 3395.090 2670.110 3396.270 ;
        RECT 2668.930 3393.490 2670.110 3394.670 ;
        RECT 2668.930 3215.090 2670.110 3216.270 ;
        RECT 2668.930 3213.490 2670.110 3214.670 ;
        RECT 2668.930 3035.090 2670.110 3036.270 ;
        RECT 2668.930 3033.490 2670.110 3034.670 ;
        RECT 2668.930 2855.090 2670.110 2856.270 ;
        RECT 2668.930 2853.490 2670.110 2854.670 ;
        RECT 2668.930 2675.090 2670.110 2676.270 ;
        RECT 2668.930 2673.490 2670.110 2674.670 ;
        RECT 2668.930 2495.090 2670.110 2496.270 ;
        RECT 2668.930 2493.490 2670.110 2494.670 ;
        RECT 2668.930 2315.090 2670.110 2316.270 ;
        RECT 2668.930 2313.490 2670.110 2314.670 ;
        RECT 2668.930 2135.090 2670.110 2136.270 ;
        RECT 2668.930 2133.490 2670.110 2134.670 ;
        RECT 2668.930 1955.090 2670.110 1956.270 ;
        RECT 2668.930 1953.490 2670.110 1954.670 ;
        RECT 2668.930 1775.090 2670.110 1776.270 ;
        RECT 2668.930 1773.490 2670.110 1774.670 ;
        RECT 2668.930 1595.090 2670.110 1596.270 ;
        RECT 2668.930 1593.490 2670.110 1594.670 ;
        RECT 2668.930 1415.090 2670.110 1416.270 ;
        RECT 2668.930 1413.490 2670.110 1414.670 ;
        RECT 2668.930 1235.090 2670.110 1236.270 ;
        RECT 2668.930 1233.490 2670.110 1234.670 ;
        RECT 2668.930 1055.090 2670.110 1056.270 ;
        RECT 2668.930 1053.490 2670.110 1054.670 ;
        RECT 2668.930 875.090 2670.110 876.270 ;
        RECT 2668.930 873.490 2670.110 874.670 ;
        RECT 2668.930 695.090 2670.110 696.270 ;
        RECT 2668.930 693.490 2670.110 694.670 ;
        RECT 2668.930 515.090 2670.110 516.270 ;
        RECT 2668.930 513.490 2670.110 514.670 ;
        RECT 2668.930 335.090 2670.110 336.270 ;
        RECT 2668.930 333.490 2670.110 334.670 ;
        RECT 2668.930 155.090 2670.110 156.270 ;
        RECT 2668.930 153.490 2670.110 154.670 ;
        RECT 2668.930 -35.110 2670.110 -33.930 ;
        RECT 2668.930 -36.710 2670.110 -35.530 ;
        RECT 2848.930 3555.210 2850.110 3556.390 ;
        RECT 2848.930 3553.610 2850.110 3554.790 ;
        RECT 2848.930 3395.090 2850.110 3396.270 ;
        RECT 2848.930 3393.490 2850.110 3394.670 ;
        RECT 2848.930 3215.090 2850.110 3216.270 ;
        RECT 2848.930 3213.490 2850.110 3214.670 ;
        RECT 2848.930 3035.090 2850.110 3036.270 ;
        RECT 2848.930 3033.490 2850.110 3034.670 ;
        RECT 2848.930 2855.090 2850.110 2856.270 ;
        RECT 2848.930 2853.490 2850.110 2854.670 ;
        RECT 2848.930 2675.090 2850.110 2676.270 ;
        RECT 2848.930 2673.490 2850.110 2674.670 ;
        RECT 2848.930 2495.090 2850.110 2496.270 ;
        RECT 2848.930 2493.490 2850.110 2494.670 ;
        RECT 2848.930 2315.090 2850.110 2316.270 ;
        RECT 2848.930 2313.490 2850.110 2314.670 ;
        RECT 2848.930 2135.090 2850.110 2136.270 ;
        RECT 2848.930 2133.490 2850.110 2134.670 ;
        RECT 2848.930 1955.090 2850.110 1956.270 ;
        RECT 2848.930 1953.490 2850.110 1954.670 ;
        RECT 2848.930 1775.090 2850.110 1776.270 ;
        RECT 2848.930 1773.490 2850.110 1774.670 ;
        RECT 2848.930 1595.090 2850.110 1596.270 ;
        RECT 2848.930 1593.490 2850.110 1594.670 ;
        RECT 2848.930 1415.090 2850.110 1416.270 ;
        RECT 2848.930 1413.490 2850.110 1414.670 ;
        RECT 2848.930 1235.090 2850.110 1236.270 ;
        RECT 2848.930 1233.490 2850.110 1234.670 ;
        RECT 2848.930 1055.090 2850.110 1056.270 ;
        RECT 2848.930 1053.490 2850.110 1054.670 ;
        RECT 2848.930 875.090 2850.110 876.270 ;
        RECT 2848.930 873.490 2850.110 874.670 ;
        RECT 2848.930 695.090 2850.110 696.270 ;
        RECT 2848.930 693.490 2850.110 694.670 ;
        RECT 2848.930 515.090 2850.110 516.270 ;
        RECT 2848.930 513.490 2850.110 514.670 ;
        RECT 2848.930 335.090 2850.110 336.270 ;
        RECT 2848.930 333.490 2850.110 334.670 ;
        RECT 2848.930 155.090 2850.110 156.270 ;
        RECT 2848.930 153.490 2850.110 154.670 ;
        RECT 2848.930 -35.110 2850.110 -33.930 ;
        RECT 2848.930 -36.710 2850.110 -35.530 ;
        RECT 2959.710 3555.210 2960.890 3556.390 ;
        RECT 2959.710 3553.610 2960.890 3554.790 ;
        RECT 2959.710 3395.090 2960.890 3396.270 ;
        RECT 2959.710 3393.490 2960.890 3394.670 ;
        RECT 2959.710 3215.090 2960.890 3216.270 ;
        RECT 2959.710 3213.490 2960.890 3214.670 ;
        RECT 2959.710 3035.090 2960.890 3036.270 ;
        RECT 2959.710 3033.490 2960.890 3034.670 ;
        RECT 2959.710 2855.090 2960.890 2856.270 ;
        RECT 2959.710 2853.490 2960.890 2854.670 ;
        RECT 2959.710 2675.090 2960.890 2676.270 ;
        RECT 2959.710 2673.490 2960.890 2674.670 ;
        RECT 2959.710 2495.090 2960.890 2496.270 ;
        RECT 2959.710 2493.490 2960.890 2494.670 ;
        RECT 2959.710 2315.090 2960.890 2316.270 ;
        RECT 2959.710 2313.490 2960.890 2314.670 ;
        RECT 2959.710 2135.090 2960.890 2136.270 ;
        RECT 2959.710 2133.490 2960.890 2134.670 ;
        RECT 2959.710 1955.090 2960.890 1956.270 ;
        RECT 2959.710 1953.490 2960.890 1954.670 ;
        RECT 2959.710 1775.090 2960.890 1776.270 ;
        RECT 2959.710 1773.490 2960.890 1774.670 ;
        RECT 2959.710 1595.090 2960.890 1596.270 ;
        RECT 2959.710 1593.490 2960.890 1594.670 ;
        RECT 2959.710 1415.090 2960.890 1416.270 ;
        RECT 2959.710 1413.490 2960.890 1414.670 ;
        RECT 2959.710 1235.090 2960.890 1236.270 ;
        RECT 2959.710 1233.490 2960.890 1234.670 ;
        RECT 2959.710 1055.090 2960.890 1056.270 ;
        RECT 2959.710 1053.490 2960.890 1054.670 ;
        RECT 2959.710 875.090 2960.890 876.270 ;
        RECT 2959.710 873.490 2960.890 874.670 ;
        RECT 2959.710 695.090 2960.890 696.270 ;
        RECT 2959.710 693.490 2960.890 694.670 ;
        RECT 2959.710 515.090 2960.890 516.270 ;
        RECT 2959.710 513.490 2960.890 514.670 ;
        RECT 2959.710 335.090 2960.890 336.270 ;
        RECT 2959.710 333.490 2960.890 334.670 ;
        RECT 2959.710 155.090 2960.890 156.270 ;
        RECT 2959.710 153.490 2960.890 154.670 ;
        RECT 2959.710 -35.110 2960.890 -33.930 ;
        RECT 2959.710 -36.710 2960.890 -35.530 ;
      LAYER met5 ;
        RECT -42.180 3556.500 -39.180 3556.510 ;
        RECT 148.020 3556.500 151.020 3556.510 ;
        RECT 328.020 3556.500 331.020 3556.510 ;
        RECT 508.020 3556.500 511.020 3556.510 ;
        RECT 688.020 3556.500 691.020 3556.510 ;
        RECT 868.020 3556.500 871.020 3556.510 ;
        RECT 1048.020 3556.500 1051.020 3556.510 ;
        RECT 1228.020 3556.500 1231.020 3556.510 ;
        RECT 1408.020 3556.500 1411.020 3556.510 ;
        RECT 1588.020 3556.500 1591.020 3556.510 ;
        RECT 1768.020 3556.500 1771.020 3556.510 ;
        RECT 1948.020 3556.500 1951.020 3556.510 ;
        RECT 2128.020 3556.500 2131.020 3556.510 ;
        RECT 2308.020 3556.500 2311.020 3556.510 ;
        RECT 2488.020 3556.500 2491.020 3556.510 ;
        RECT 2668.020 3556.500 2671.020 3556.510 ;
        RECT 2848.020 3556.500 2851.020 3556.510 ;
        RECT 2958.800 3556.500 2961.800 3556.510 ;
        RECT -42.180 3553.500 2961.800 3556.500 ;
        RECT -42.180 3553.490 -39.180 3553.500 ;
        RECT 148.020 3553.490 151.020 3553.500 ;
        RECT 328.020 3553.490 331.020 3553.500 ;
        RECT 508.020 3553.490 511.020 3553.500 ;
        RECT 688.020 3553.490 691.020 3553.500 ;
        RECT 868.020 3553.490 871.020 3553.500 ;
        RECT 1048.020 3553.490 1051.020 3553.500 ;
        RECT 1228.020 3553.490 1231.020 3553.500 ;
        RECT 1408.020 3553.490 1411.020 3553.500 ;
        RECT 1588.020 3553.490 1591.020 3553.500 ;
        RECT 1768.020 3553.490 1771.020 3553.500 ;
        RECT 1948.020 3553.490 1951.020 3553.500 ;
        RECT 2128.020 3553.490 2131.020 3553.500 ;
        RECT 2308.020 3553.490 2311.020 3553.500 ;
        RECT 2488.020 3553.490 2491.020 3553.500 ;
        RECT 2668.020 3553.490 2671.020 3553.500 ;
        RECT 2848.020 3553.490 2851.020 3553.500 ;
        RECT 2958.800 3553.490 2961.800 3553.500 ;
        RECT -42.180 3396.380 -39.180 3396.390 ;
        RECT 148.020 3396.380 151.020 3396.390 ;
        RECT 328.020 3396.380 331.020 3396.390 ;
        RECT 508.020 3396.380 511.020 3396.390 ;
        RECT 688.020 3396.380 691.020 3396.390 ;
        RECT 868.020 3396.380 871.020 3396.390 ;
        RECT 1048.020 3396.380 1051.020 3396.390 ;
        RECT 1228.020 3396.380 1231.020 3396.390 ;
        RECT 1408.020 3396.380 1411.020 3396.390 ;
        RECT 1588.020 3396.380 1591.020 3396.390 ;
        RECT 1768.020 3396.380 1771.020 3396.390 ;
        RECT 1948.020 3396.380 1951.020 3396.390 ;
        RECT 2128.020 3396.380 2131.020 3396.390 ;
        RECT 2308.020 3396.380 2311.020 3396.390 ;
        RECT 2488.020 3396.380 2491.020 3396.390 ;
        RECT 2668.020 3396.380 2671.020 3396.390 ;
        RECT 2848.020 3396.380 2851.020 3396.390 ;
        RECT 2958.800 3396.380 2961.800 3396.390 ;
        RECT -42.180 3393.380 2961.800 3396.380 ;
        RECT -42.180 3393.370 -39.180 3393.380 ;
        RECT 148.020 3393.370 151.020 3393.380 ;
        RECT 328.020 3393.370 331.020 3393.380 ;
        RECT 508.020 3393.370 511.020 3393.380 ;
        RECT 688.020 3393.370 691.020 3393.380 ;
        RECT 868.020 3393.370 871.020 3393.380 ;
        RECT 1048.020 3393.370 1051.020 3393.380 ;
        RECT 1228.020 3393.370 1231.020 3393.380 ;
        RECT 1408.020 3393.370 1411.020 3393.380 ;
        RECT 1588.020 3393.370 1591.020 3393.380 ;
        RECT 1768.020 3393.370 1771.020 3393.380 ;
        RECT 1948.020 3393.370 1951.020 3393.380 ;
        RECT 2128.020 3393.370 2131.020 3393.380 ;
        RECT 2308.020 3393.370 2311.020 3393.380 ;
        RECT 2488.020 3393.370 2491.020 3393.380 ;
        RECT 2668.020 3393.370 2671.020 3393.380 ;
        RECT 2848.020 3393.370 2851.020 3393.380 ;
        RECT 2958.800 3393.370 2961.800 3393.380 ;
        RECT -42.180 3216.380 -39.180 3216.390 ;
        RECT 148.020 3216.380 151.020 3216.390 ;
        RECT 328.020 3216.380 331.020 3216.390 ;
        RECT 508.020 3216.380 511.020 3216.390 ;
        RECT 688.020 3216.380 691.020 3216.390 ;
        RECT 868.020 3216.380 871.020 3216.390 ;
        RECT 1048.020 3216.380 1051.020 3216.390 ;
        RECT 1228.020 3216.380 1231.020 3216.390 ;
        RECT 1408.020 3216.380 1411.020 3216.390 ;
        RECT 1588.020 3216.380 1591.020 3216.390 ;
        RECT 1768.020 3216.380 1771.020 3216.390 ;
        RECT 1948.020 3216.380 1951.020 3216.390 ;
        RECT 2128.020 3216.380 2131.020 3216.390 ;
        RECT 2308.020 3216.380 2311.020 3216.390 ;
        RECT 2488.020 3216.380 2491.020 3216.390 ;
        RECT 2668.020 3216.380 2671.020 3216.390 ;
        RECT 2848.020 3216.380 2851.020 3216.390 ;
        RECT 2958.800 3216.380 2961.800 3216.390 ;
        RECT -42.180 3213.380 2961.800 3216.380 ;
        RECT -42.180 3213.370 -39.180 3213.380 ;
        RECT 148.020 3213.370 151.020 3213.380 ;
        RECT 328.020 3213.370 331.020 3213.380 ;
        RECT 508.020 3213.370 511.020 3213.380 ;
        RECT 688.020 3213.370 691.020 3213.380 ;
        RECT 868.020 3213.370 871.020 3213.380 ;
        RECT 1048.020 3213.370 1051.020 3213.380 ;
        RECT 1228.020 3213.370 1231.020 3213.380 ;
        RECT 1408.020 3213.370 1411.020 3213.380 ;
        RECT 1588.020 3213.370 1591.020 3213.380 ;
        RECT 1768.020 3213.370 1771.020 3213.380 ;
        RECT 1948.020 3213.370 1951.020 3213.380 ;
        RECT 2128.020 3213.370 2131.020 3213.380 ;
        RECT 2308.020 3213.370 2311.020 3213.380 ;
        RECT 2488.020 3213.370 2491.020 3213.380 ;
        RECT 2668.020 3213.370 2671.020 3213.380 ;
        RECT 2848.020 3213.370 2851.020 3213.380 ;
        RECT 2958.800 3213.370 2961.800 3213.380 ;
        RECT -42.180 3036.380 -39.180 3036.390 ;
        RECT 148.020 3036.380 151.020 3036.390 ;
        RECT 328.020 3036.380 331.020 3036.390 ;
        RECT 508.020 3036.380 511.020 3036.390 ;
        RECT 688.020 3036.380 691.020 3036.390 ;
        RECT 868.020 3036.380 871.020 3036.390 ;
        RECT 1048.020 3036.380 1051.020 3036.390 ;
        RECT 1228.020 3036.380 1231.020 3036.390 ;
        RECT 1408.020 3036.380 1411.020 3036.390 ;
        RECT 1588.020 3036.380 1591.020 3036.390 ;
        RECT 1768.020 3036.380 1771.020 3036.390 ;
        RECT 1948.020 3036.380 1951.020 3036.390 ;
        RECT 2128.020 3036.380 2131.020 3036.390 ;
        RECT 2308.020 3036.380 2311.020 3036.390 ;
        RECT 2488.020 3036.380 2491.020 3036.390 ;
        RECT 2668.020 3036.380 2671.020 3036.390 ;
        RECT 2848.020 3036.380 2851.020 3036.390 ;
        RECT 2958.800 3036.380 2961.800 3036.390 ;
        RECT -42.180 3033.380 2961.800 3036.380 ;
        RECT -42.180 3033.370 -39.180 3033.380 ;
        RECT 148.020 3033.370 151.020 3033.380 ;
        RECT 328.020 3033.370 331.020 3033.380 ;
        RECT 508.020 3033.370 511.020 3033.380 ;
        RECT 688.020 3033.370 691.020 3033.380 ;
        RECT 868.020 3033.370 871.020 3033.380 ;
        RECT 1048.020 3033.370 1051.020 3033.380 ;
        RECT 1228.020 3033.370 1231.020 3033.380 ;
        RECT 1408.020 3033.370 1411.020 3033.380 ;
        RECT 1588.020 3033.370 1591.020 3033.380 ;
        RECT 1768.020 3033.370 1771.020 3033.380 ;
        RECT 1948.020 3033.370 1951.020 3033.380 ;
        RECT 2128.020 3033.370 2131.020 3033.380 ;
        RECT 2308.020 3033.370 2311.020 3033.380 ;
        RECT 2488.020 3033.370 2491.020 3033.380 ;
        RECT 2668.020 3033.370 2671.020 3033.380 ;
        RECT 2848.020 3033.370 2851.020 3033.380 ;
        RECT 2958.800 3033.370 2961.800 3033.380 ;
        RECT -42.180 2856.380 -39.180 2856.390 ;
        RECT 148.020 2856.380 151.020 2856.390 ;
        RECT 328.020 2856.380 331.020 2856.390 ;
        RECT 508.020 2856.380 511.020 2856.390 ;
        RECT 688.020 2856.380 691.020 2856.390 ;
        RECT 868.020 2856.380 871.020 2856.390 ;
        RECT 1048.020 2856.380 1051.020 2856.390 ;
        RECT 1228.020 2856.380 1231.020 2856.390 ;
        RECT 1408.020 2856.380 1411.020 2856.390 ;
        RECT 1588.020 2856.380 1591.020 2856.390 ;
        RECT 1768.020 2856.380 1771.020 2856.390 ;
        RECT 1948.020 2856.380 1951.020 2856.390 ;
        RECT 2128.020 2856.380 2131.020 2856.390 ;
        RECT 2308.020 2856.380 2311.020 2856.390 ;
        RECT 2488.020 2856.380 2491.020 2856.390 ;
        RECT 2668.020 2856.380 2671.020 2856.390 ;
        RECT 2848.020 2856.380 2851.020 2856.390 ;
        RECT 2958.800 2856.380 2961.800 2856.390 ;
        RECT -42.180 2853.380 2961.800 2856.380 ;
        RECT -42.180 2853.370 -39.180 2853.380 ;
        RECT 148.020 2853.370 151.020 2853.380 ;
        RECT 328.020 2853.370 331.020 2853.380 ;
        RECT 508.020 2853.370 511.020 2853.380 ;
        RECT 688.020 2853.370 691.020 2853.380 ;
        RECT 868.020 2853.370 871.020 2853.380 ;
        RECT 1048.020 2853.370 1051.020 2853.380 ;
        RECT 1228.020 2853.370 1231.020 2853.380 ;
        RECT 1408.020 2853.370 1411.020 2853.380 ;
        RECT 1588.020 2853.370 1591.020 2853.380 ;
        RECT 1768.020 2853.370 1771.020 2853.380 ;
        RECT 1948.020 2853.370 1951.020 2853.380 ;
        RECT 2128.020 2853.370 2131.020 2853.380 ;
        RECT 2308.020 2853.370 2311.020 2853.380 ;
        RECT 2488.020 2853.370 2491.020 2853.380 ;
        RECT 2668.020 2853.370 2671.020 2853.380 ;
        RECT 2848.020 2853.370 2851.020 2853.380 ;
        RECT 2958.800 2853.370 2961.800 2853.380 ;
        RECT -42.180 2676.380 -39.180 2676.390 ;
        RECT 148.020 2676.380 151.020 2676.390 ;
        RECT 328.020 2676.380 331.020 2676.390 ;
        RECT 508.020 2676.380 511.020 2676.390 ;
        RECT 688.020 2676.380 691.020 2676.390 ;
        RECT 868.020 2676.380 871.020 2676.390 ;
        RECT 1048.020 2676.380 1051.020 2676.390 ;
        RECT 1228.020 2676.380 1231.020 2676.390 ;
        RECT 1408.020 2676.380 1411.020 2676.390 ;
        RECT 1588.020 2676.380 1591.020 2676.390 ;
        RECT 1768.020 2676.380 1771.020 2676.390 ;
        RECT 1948.020 2676.380 1951.020 2676.390 ;
        RECT 2128.020 2676.380 2131.020 2676.390 ;
        RECT 2308.020 2676.380 2311.020 2676.390 ;
        RECT 2488.020 2676.380 2491.020 2676.390 ;
        RECT 2668.020 2676.380 2671.020 2676.390 ;
        RECT 2848.020 2676.380 2851.020 2676.390 ;
        RECT 2958.800 2676.380 2961.800 2676.390 ;
        RECT -42.180 2673.380 2961.800 2676.380 ;
        RECT -42.180 2673.370 -39.180 2673.380 ;
        RECT 148.020 2673.370 151.020 2673.380 ;
        RECT 328.020 2673.370 331.020 2673.380 ;
        RECT 508.020 2673.370 511.020 2673.380 ;
        RECT 688.020 2673.370 691.020 2673.380 ;
        RECT 868.020 2673.370 871.020 2673.380 ;
        RECT 1048.020 2673.370 1051.020 2673.380 ;
        RECT 1228.020 2673.370 1231.020 2673.380 ;
        RECT 1408.020 2673.370 1411.020 2673.380 ;
        RECT 1588.020 2673.370 1591.020 2673.380 ;
        RECT 1768.020 2673.370 1771.020 2673.380 ;
        RECT 1948.020 2673.370 1951.020 2673.380 ;
        RECT 2128.020 2673.370 2131.020 2673.380 ;
        RECT 2308.020 2673.370 2311.020 2673.380 ;
        RECT 2488.020 2673.370 2491.020 2673.380 ;
        RECT 2668.020 2673.370 2671.020 2673.380 ;
        RECT 2848.020 2673.370 2851.020 2673.380 ;
        RECT 2958.800 2673.370 2961.800 2673.380 ;
        RECT -42.180 2496.380 -39.180 2496.390 ;
        RECT 148.020 2496.380 151.020 2496.390 ;
        RECT 328.020 2496.380 331.020 2496.390 ;
        RECT 508.020 2496.380 511.020 2496.390 ;
        RECT 688.020 2496.380 691.020 2496.390 ;
        RECT 868.020 2496.380 871.020 2496.390 ;
        RECT 1048.020 2496.380 1051.020 2496.390 ;
        RECT 1228.020 2496.380 1231.020 2496.390 ;
        RECT 1408.020 2496.380 1411.020 2496.390 ;
        RECT 1588.020 2496.380 1591.020 2496.390 ;
        RECT 1768.020 2496.380 1771.020 2496.390 ;
        RECT 1948.020 2496.380 1951.020 2496.390 ;
        RECT 2128.020 2496.380 2131.020 2496.390 ;
        RECT 2308.020 2496.380 2311.020 2496.390 ;
        RECT 2488.020 2496.380 2491.020 2496.390 ;
        RECT 2668.020 2496.380 2671.020 2496.390 ;
        RECT 2848.020 2496.380 2851.020 2496.390 ;
        RECT 2958.800 2496.380 2961.800 2496.390 ;
        RECT -42.180 2493.380 2961.800 2496.380 ;
        RECT -42.180 2493.370 -39.180 2493.380 ;
        RECT 148.020 2493.370 151.020 2493.380 ;
        RECT 328.020 2493.370 331.020 2493.380 ;
        RECT 508.020 2493.370 511.020 2493.380 ;
        RECT 688.020 2493.370 691.020 2493.380 ;
        RECT 868.020 2493.370 871.020 2493.380 ;
        RECT 1048.020 2493.370 1051.020 2493.380 ;
        RECT 1228.020 2493.370 1231.020 2493.380 ;
        RECT 1408.020 2493.370 1411.020 2493.380 ;
        RECT 1588.020 2493.370 1591.020 2493.380 ;
        RECT 1768.020 2493.370 1771.020 2493.380 ;
        RECT 1948.020 2493.370 1951.020 2493.380 ;
        RECT 2128.020 2493.370 2131.020 2493.380 ;
        RECT 2308.020 2493.370 2311.020 2493.380 ;
        RECT 2488.020 2493.370 2491.020 2493.380 ;
        RECT 2668.020 2493.370 2671.020 2493.380 ;
        RECT 2848.020 2493.370 2851.020 2493.380 ;
        RECT 2958.800 2493.370 2961.800 2493.380 ;
        RECT -42.180 2316.380 -39.180 2316.390 ;
        RECT 148.020 2316.380 151.020 2316.390 ;
        RECT 328.020 2316.380 331.020 2316.390 ;
        RECT 508.020 2316.380 511.020 2316.390 ;
        RECT 688.020 2316.380 691.020 2316.390 ;
        RECT 868.020 2316.380 871.020 2316.390 ;
        RECT 1048.020 2316.380 1051.020 2316.390 ;
        RECT 1228.020 2316.380 1231.020 2316.390 ;
        RECT 1408.020 2316.380 1411.020 2316.390 ;
        RECT 1588.020 2316.380 1591.020 2316.390 ;
        RECT 1768.020 2316.380 1771.020 2316.390 ;
        RECT 1948.020 2316.380 1951.020 2316.390 ;
        RECT 2128.020 2316.380 2131.020 2316.390 ;
        RECT 2308.020 2316.380 2311.020 2316.390 ;
        RECT 2488.020 2316.380 2491.020 2316.390 ;
        RECT 2668.020 2316.380 2671.020 2316.390 ;
        RECT 2848.020 2316.380 2851.020 2316.390 ;
        RECT 2958.800 2316.380 2961.800 2316.390 ;
        RECT -42.180 2313.380 2961.800 2316.380 ;
        RECT -42.180 2313.370 -39.180 2313.380 ;
        RECT 148.020 2313.370 151.020 2313.380 ;
        RECT 328.020 2313.370 331.020 2313.380 ;
        RECT 508.020 2313.370 511.020 2313.380 ;
        RECT 688.020 2313.370 691.020 2313.380 ;
        RECT 868.020 2313.370 871.020 2313.380 ;
        RECT 1048.020 2313.370 1051.020 2313.380 ;
        RECT 1228.020 2313.370 1231.020 2313.380 ;
        RECT 1408.020 2313.370 1411.020 2313.380 ;
        RECT 1588.020 2313.370 1591.020 2313.380 ;
        RECT 1768.020 2313.370 1771.020 2313.380 ;
        RECT 1948.020 2313.370 1951.020 2313.380 ;
        RECT 2128.020 2313.370 2131.020 2313.380 ;
        RECT 2308.020 2313.370 2311.020 2313.380 ;
        RECT 2488.020 2313.370 2491.020 2313.380 ;
        RECT 2668.020 2313.370 2671.020 2313.380 ;
        RECT 2848.020 2313.370 2851.020 2313.380 ;
        RECT 2958.800 2313.370 2961.800 2313.380 ;
        RECT -42.180 2136.380 -39.180 2136.390 ;
        RECT 148.020 2136.380 151.020 2136.390 ;
        RECT 328.020 2136.380 331.020 2136.390 ;
        RECT 508.020 2136.380 511.020 2136.390 ;
        RECT 688.020 2136.380 691.020 2136.390 ;
        RECT 868.020 2136.380 871.020 2136.390 ;
        RECT 1048.020 2136.380 1051.020 2136.390 ;
        RECT 1228.020 2136.380 1231.020 2136.390 ;
        RECT 1408.020 2136.380 1411.020 2136.390 ;
        RECT 1588.020 2136.380 1591.020 2136.390 ;
        RECT 1768.020 2136.380 1771.020 2136.390 ;
        RECT 1948.020 2136.380 1951.020 2136.390 ;
        RECT 2128.020 2136.380 2131.020 2136.390 ;
        RECT 2308.020 2136.380 2311.020 2136.390 ;
        RECT 2488.020 2136.380 2491.020 2136.390 ;
        RECT 2668.020 2136.380 2671.020 2136.390 ;
        RECT 2848.020 2136.380 2851.020 2136.390 ;
        RECT 2958.800 2136.380 2961.800 2136.390 ;
        RECT -42.180 2133.380 2961.800 2136.380 ;
        RECT -42.180 2133.370 -39.180 2133.380 ;
        RECT 148.020 2133.370 151.020 2133.380 ;
        RECT 328.020 2133.370 331.020 2133.380 ;
        RECT 508.020 2133.370 511.020 2133.380 ;
        RECT 688.020 2133.370 691.020 2133.380 ;
        RECT 868.020 2133.370 871.020 2133.380 ;
        RECT 1048.020 2133.370 1051.020 2133.380 ;
        RECT 1228.020 2133.370 1231.020 2133.380 ;
        RECT 1408.020 2133.370 1411.020 2133.380 ;
        RECT 1588.020 2133.370 1591.020 2133.380 ;
        RECT 1768.020 2133.370 1771.020 2133.380 ;
        RECT 1948.020 2133.370 1951.020 2133.380 ;
        RECT 2128.020 2133.370 2131.020 2133.380 ;
        RECT 2308.020 2133.370 2311.020 2133.380 ;
        RECT 2488.020 2133.370 2491.020 2133.380 ;
        RECT 2668.020 2133.370 2671.020 2133.380 ;
        RECT 2848.020 2133.370 2851.020 2133.380 ;
        RECT 2958.800 2133.370 2961.800 2133.380 ;
        RECT -42.180 1956.380 -39.180 1956.390 ;
        RECT 148.020 1956.380 151.020 1956.390 ;
        RECT 328.020 1956.380 331.020 1956.390 ;
        RECT 508.020 1956.380 511.020 1956.390 ;
        RECT 688.020 1956.380 691.020 1956.390 ;
        RECT 868.020 1956.380 871.020 1956.390 ;
        RECT 1048.020 1956.380 1051.020 1956.390 ;
        RECT 1228.020 1956.380 1231.020 1956.390 ;
        RECT 1408.020 1956.380 1411.020 1956.390 ;
        RECT 1588.020 1956.380 1591.020 1956.390 ;
        RECT 1768.020 1956.380 1771.020 1956.390 ;
        RECT 1948.020 1956.380 1951.020 1956.390 ;
        RECT 2128.020 1956.380 2131.020 1956.390 ;
        RECT 2308.020 1956.380 2311.020 1956.390 ;
        RECT 2488.020 1956.380 2491.020 1956.390 ;
        RECT 2668.020 1956.380 2671.020 1956.390 ;
        RECT 2848.020 1956.380 2851.020 1956.390 ;
        RECT 2958.800 1956.380 2961.800 1956.390 ;
        RECT -42.180 1953.380 2961.800 1956.380 ;
        RECT -42.180 1953.370 -39.180 1953.380 ;
        RECT 148.020 1953.370 151.020 1953.380 ;
        RECT 328.020 1953.370 331.020 1953.380 ;
        RECT 508.020 1953.370 511.020 1953.380 ;
        RECT 688.020 1953.370 691.020 1953.380 ;
        RECT 868.020 1953.370 871.020 1953.380 ;
        RECT 1048.020 1953.370 1051.020 1953.380 ;
        RECT 1228.020 1953.370 1231.020 1953.380 ;
        RECT 1408.020 1953.370 1411.020 1953.380 ;
        RECT 1588.020 1953.370 1591.020 1953.380 ;
        RECT 1768.020 1953.370 1771.020 1953.380 ;
        RECT 1948.020 1953.370 1951.020 1953.380 ;
        RECT 2128.020 1953.370 2131.020 1953.380 ;
        RECT 2308.020 1953.370 2311.020 1953.380 ;
        RECT 2488.020 1953.370 2491.020 1953.380 ;
        RECT 2668.020 1953.370 2671.020 1953.380 ;
        RECT 2848.020 1953.370 2851.020 1953.380 ;
        RECT 2958.800 1953.370 2961.800 1953.380 ;
        RECT -42.180 1776.380 -39.180 1776.390 ;
        RECT 148.020 1776.380 151.020 1776.390 ;
        RECT 328.020 1776.380 331.020 1776.390 ;
        RECT 508.020 1776.380 511.020 1776.390 ;
        RECT 688.020 1776.380 691.020 1776.390 ;
        RECT 868.020 1776.380 871.020 1776.390 ;
        RECT 1048.020 1776.380 1051.020 1776.390 ;
        RECT 1228.020 1776.380 1231.020 1776.390 ;
        RECT 1408.020 1776.380 1411.020 1776.390 ;
        RECT 1588.020 1776.380 1591.020 1776.390 ;
        RECT 1768.020 1776.380 1771.020 1776.390 ;
        RECT 1948.020 1776.380 1951.020 1776.390 ;
        RECT 2128.020 1776.380 2131.020 1776.390 ;
        RECT 2308.020 1776.380 2311.020 1776.390 ;
        RECT 2488.020 1776.380 2491.020 1776.390 ;
        RECT 2668.020 1776.380 2671.020 1776.390 ;
        RECT 2848.020 1776.380 2851.020 1776.390 ;
        RECT 2958.800 1776.380 2961.800 1776.390 ;
        RECT -42.180 1773.380 2961.800 1776.380 ;
        RECT -42.180 1773.370 -39.180 1773.380 ;
        RECT 148.020 1773.370 151.020 1773.380 ;
        RECT 328.020 1773.370 331.020 1773.380 ;
        RECT 508.020 1773.370 511.020 1773.380 ;
        RECT 688.020 1773.370 691.020 1773.380 ;
        RECT 868.020 1773.370 871.020 1773.380 ;
        RECT 1048.020 1773.370 1051.020 1773.380 ;
        RECT 1228.020 1773.370 1231.020 1773.380 ;
        RECT 1408.020 1773.370 1411.020 1773.380 ;
        RECT 1588.020 1773.370 1591.020 1773.380 ;
        RECT 1768.020 1773.370 1771.020 1773.380 ;
        RECT 1948.020 1773.370 1951.020 1773.380 ;
        RECT 2128.020 1773.370 2131.020 1773.380 ;
        RECT 2308.020 1773.370 2311.020 1773.380 ;
        RECT 2488.020 1773.370 2491.020 1773.380 ;
        RECT 2668.020 1773.370 2671.020 1773.380 ;
        RECT 2848.020 1773.370 2851.020 1773.380 ;
        RECT 2958.800 1773.370 2961.800 1773.380 ;
        RECT -42.180 1596.380 -39.180 1596.390 ;
        RECT 148.020 1596.380 151.020 1596.390 ;
        RECT 328.020 1596.380 331.020 1596.390 ;
        RECT 508.020 1596.380 511.020 1596.390 ;
        RECT 688.020 1596.380 691.020 1596.390 ;
        RECT 868.020 1596.380 871.020 1596.390 ;
        RECT 1048.020 1596.380 1051.020 1596.390 ;
        RECT 1228.020 1596.380 1231.020 1596.390 ;
        RECT 1408.020 1596.380 1411.020 1596.390 ;
        RECT 1588.020 1596.380 1591.020 1596.390 ;
        RECT 1768.020 1596.380 1771.020 1596.390 ;
        RECT 1948.020 1596.380 1951.020 1596.390 ;
        RECT 2128.020 1596.380 2131.020 1596.390 ;
        RECT 2308.020 1596.380 2311.020 1596.390 ;
        RECT 2488.020 1596.380 2491.020 1596.390 ;
        RECT 2668.020 1596.380 2671.020 1596.390 ;
        RECT 2848.020 1596.380 2851.020 1596.390 ;
        RECT 2958.800 1596.380 2961.800 1596.390 ;
        RECT -42.180 1593.380 2961.800 1596.380 ;
        RECT -42.180 1593.370 -39.180 1593.380 ;
        RECT 148.020 1593.370 151.020 1593.380 ;
        RECT 328.020 1593.370 331.020 1593.380 ;
        RECT 508.020 1593.370 511.020 1593.380 ;
        RECT 688.020 1593.370 691.020 1593.380 ;
        RECT 868.020 1593.370 871.020 1593.380 ;
        RECT 1048.020 1593.370 1051.020 1593.380 ;
        RECT 1228.020 1593.370 1231.020 1593.380 ;
        RECT 1408.020 1593.370 1411.020 1593.380 ;
        RECT 1588.020 1593.370 1591.020 1593.380 ;
        RECT 1768.020 1593.370 1771.020 1593.380 ;
        RECT 1948.020 1593.370 1951.020 1593.380 ;
        RECT 2128.020 1593.370 2131.020 1593.380 ;
        RECT 2308.020 1593.370 2311.020 1593.380 ;
        RECT 2488.020 1593.370 2491.020 1593.380 ;
        RECT 2668.020 1593.370 2671.020 1593.380 ;
        RECT 2848.020 1593.370 2851.020 1593.380 ;
        RECT 2958.800 1593.370 2961.800 1593.380 ;
        RECT -42.180 1416.380 -39.180 1416.390 ;
        RECT 148.020 1416.380 151.020 1416.390 ;
        RECT 328.020 1416.380 331.020 1416.390 ;
        RECT 508.020 1416.380 511.020 1416.390 ;
        RECT 688.020 1416.380 691.020 1416.390 ;
        RECT 868.020 1416.380 871.020 1416.390 ;
        RECT 1048.020 1416.380 1051.020 1416.390 ;
        RECT 1228.020 1416.380 1231.020 1416.390 ;
        RECT 1408.020 1416.380 1411.020 1416.390 ;
        RECT 1588.020 1416.380 1591.020 1416.390 ;
        RECT 1768.020 1416.380 1771.020 1416.390 ;
        RECT 1948.020 1416.380 1951.020 1416.390 ;
        RECT 2128.020 1416.380 2131.020 1416.390 ;
        RECT 2308.020 1416.380 2311.020 1416.390 ;
        RECT 2488.020 1416.380 2491.020 1416.390 ;
        RECT 2668.020 1416.380 2671.020 1416.390 ;
        RECT 2848.020 1416.380 2851.020 1416.390 ;
        RECT 2958.800 1416.380 2961.800 1416.390 ;
        RECT -42.180 1413.380 2961.800 1416.380 ;
        RECT -42.180 1413.370 -39.180 1413.380 ;
        RECT 148.020 1413.370 151.020 1413.380 ;
        RECT 328.020 1413.370 331.020 1413.380 ;
        RECT 508.020 1413.370 511.020 1413.380 ;
        RECT 688.020 1413.370 691.020 1413.380 ;
        RECT 868.020 1413.370 871.020 1413.380 ;
        RECT 1048.020 1413.370 1051.020 1413.380 ;
        RECT 1228.020 1413.370 1231.020 1413.380 ;
        RECT 1408.020 1413.370 1411.020 1413.380 ;
        RECT 1588.020 1413.370 1591.020 1413.380 ;
        RECT 1768.020 1413.370 1771.020 1413.380 ;
        RECT 1948.020 1413.370 1951.020 1413.380 ;
        RECT 2128.020 1413.370 2131.020 1413.380 ;
        RECT 2308.020 1413.370 2311.020 1413.380 ;
        RECT 2488.020 1413.370 2491.020 1413.380 ;
        RECT 2668.020 1413.370 2671.020 1413.380 ;
        RECT 2848.020 1413.370 2851.020 1413.380 ;
        RECT 2958.800 1413.370 2961.800 1413.380 ;
        RECT -42.180 1236.380 -39.180 1236.390 ;
        RECT 148.020 1236.380 151.020 1236.390 ;
        RECT 328.020 1236.380 331.020 1236.390 ;
        RECT 508.020 1236.380 511.020 1236.390 ;
        RECT 688.020 1236.380 691.020 1236.390 ;
        RECT 868.020 1236.380 871.020 1236.390 ;
        RECT 1048.020 1236.380 1051.020 1236.390 ;
        RECT 1228.020 1236.380 1231.020 1236.390 ;
        RECT 1408.020 1236.380 1411.020 1236.390 ;
        RECT 1588.020 1236.380 1591.020 1236.390 ;
        RECT 1768.020 1236.380 1771.020 1236.390 ;
        RECT 1948.020 1236.380 1951.020 1236.390 ;
        RECT 2128.020 1236.380 2131.020 1236.390 ;
        RECT 2308.020 1236.380 2311.020 1236.390 ;
        RECT 2488.020 1236.380 2491.020 1236.390 ;
        RECT 2668.020 1236.380 2671.020 1236.390 ;
        RECT 2848.020 1236.380 2851.020 1236.390 ;
        RECT 2958.800 1236.380 2961.800 1236.390 ;
        RECT -42.180 1233.380 2961.800 1236.380 ;
        RECT -42.180 1233.370 -39.180 1233.380 ;
        RECT 148.020 1233.370 151.020 1233.380 ;
        RECT 328.020 1233.370 331.020 1233.380 ;
        RECT 508.020 1233.370 511.020 1233.380 ;
        RECT 688.020 1233.370 691.020 1233.380 ;
        RECT 868.020 1233.370 871.020 1233.380 ;
        RECT 1048.020 1233.370 1051.020 1233.380 ;
        RECT 1228.020 1233.370 1231.020 1233.380 ;
        RECT 1408.020 1233.370 1411.020 1233.380 ;
        RECT 1588.020 1233.370 1591.020 1233.380 ;
        RECT 1768.020 1233.370 1771.020 1233.380 ;
        RECT 1948.020 1233.370 1951.020 1233.380 ;
        RECT 2128.020 1233.370 2131.020 1233.380 ;
        RECT 2308.020 1233.370 2311.020 1233.380 ;
        RECT 2488.020 1233.370 2491.020 1233.380 ;
        RECT 2668.020 1233.370 2671.020 1233.380 ;
        RECT 2848.020 1233.370 2851.020 1233.380 ;
        RECT 2958.800 1233.370 2961.800 1233.380 ;
        RECT -42.180 1056.380 -39.180 1056.390 ;
        RECT 148.020 1056.380 151.020 1056.390 ;
        RECT 328.020 1056.380 331.020 1056.390 ;
        RECT 508.020 1056.380 511.020 1056.390 ;
        RECT 688.020 1056.380 691.020 1056.390 ;
        RECT 868.020 1056.380 871.020 1056.390 ;
        RECT 1048.020 1056.380 1051.020 1056.390 ;
        RECT 1228.020 1056.380 1231.020 1056.390 ;
        RECT 1408.020 1056.380 1411.020 1056.390 ;
        RECT 1588.020 1056.380 1591.020 1056.390 ;
        RECT 1768.020 1056.380 1771.020 1056.390 ;
        RECT 1948.020 1056.380 1951.020 1056.390 ;
        RECT 2128.020 1056.380 2131.020 1056.390 ;
        RECT 2308.020 1056.380 2311.020 1056.390 ;
        RECT 2488.020 1056.380 2491.020 1056.390 ;
        RECT 2668.020 1056.380 2671.020 1056.390 ;
        RECT 2848.020 1056.380 2851.020 1056.390 ;
        RECT 2958.800 1056.380 2961.800 1056.390 ;
        RECT -42.180 1053.380 2961.800 1056.380 ;
        RECT -42.180 1053.370 -39.180 1053.380 ;
        RECT 148.020 1053.370 151.020 1053.380 ;
        RECT 328.020 1053.370 331.020 1053.380 ;
        RECT 508.020 1053.370 511.020 1053.380 ;
        RECT 688.020 1053.370 691.020 1053.380 ;
        RECT 868.020 1053.370 871.020 1053.380 ;
        RECT 1048.020 1053.370 1051.020 1053.380 ;
        RECT 1228.020 1053.370 1231.020 1053.380 ;
        RECT 1408.020 1053.370 1411.020 1053.380 ;
        RECT 1588.020 1053.370 1591.020 1053.380 ;
        RECT 1768.020 1053.370 1771.020 1053.380 ;
        RECT 1948.020 1053.370 1951.020 1053.380 ;
        RECT 2128.020 1053.370 2131.020 1053.380 ;
        RECT 2308.020 1053.370 2311.020 1053.380 ;
        RECT 2488.020 1053.370 2491.020 1053.380 ;
        RECT 2668.020 1053.370 2671.020 1053.380 ;
        RECT 2848.020 1053.370 2851.020 1053.380 ;
        RECT 2958.800 1053.370 2961.800 1053.380 ;
        RECT -42.180 876.380 -39.180 876.390 ;
        RECT 148.020 876.380 151.020 876.390 ;
        RECT 328.020 876.380 331.020 876.390 ;
        RECT 508.020 876.380 511.020 876.390 ;
        RECT 688.020 876.380 691.020 876.390 ;
        RECT 868.020 876.380 871.020 876.390 ;
        RECT 1048.020 876.380 1051.020 876.390 ;
        RECT 1228.020 876.380 1231.020 876.390 ;
        RECT 1408.020 876.380 1411.020 876.390 ;
        RECT 1588.020 876.380 1591.020 876.390 ;
        RECT 1768.020 876.380 1771.020 876.390 ;
        RECT 1948.020 876.380 1951.020 876.390 ;
        RECT 2128.020 876.380 2131.020 876.390 ;
        RECT 2308.020 876.380 2311.020 876.390 ;
        RECT 2488.020 876.380 2491.020 876.390 ;
        RECT 2668.020 876.380 2671.020 876.390 ;
        RECT 2848.020 876.380 2851.020 876.390 ;
        RECT 2958.800 876.380 2961.800 876.390 ;
        RECT -42.180 873.380 2961.800 876.380 ;
        RECT -42.180 873.370 -39.180 873.380 ;
        RECT 148.020 873.370 151.020 873.380 ;
        RECT 328.020 873.370 331.020 873.380 ;
        RECT 508.020 873.370 511.020 873.380 ;
        RECT 688.020 873.370 691.020 873.380 ;
        RECT 868.020 873.370 871.020 873.380 ;
        RECT 1048.020 873.370 1051.020 873.380 ;
        RECT 1228.020 873.370 1231.020 873.380 ;
        RECT 1408.020 873.370 1411.020 873.380 ;
        RECT 1588.020 873.370 1591.020 873.380 ;
        RECT 1768.020 873.370 1771.020 873.380 ;
        RECT 1948.020 873.370 1951.020 873.380 ;
        RECT 2128.020 873.370 2131.020 873.380 ;
        RECT 2308.020 873.370 2311.020 873.380 ;
        RECT 2488.020 873.370 2491.020 873.380 ;
        RECT 2668.020 873.370 2671.020 873.380 ;
        RECT 2848.020 873.370 2851.020 873.380 ;
        RECT 2958.800 873.370 2961.800 873.380 ;
        RECT -42.180 696.380 -39.180 696.390 ;
        RECT 148.020 696.380 151.020 696.390 ;
        RECT 328.020 696.380 331.020 696.390 ;
        RECT 508.020 696.380 511.020 696.390 ;
        RECT 688.020 696.380 691.020 696.390 ;
        RECT 868.020 696.380 871.020 696.390 ;
        RECT 1048.020 696.380 1051.020 696.390 ;
        RECT 1228.020 696.380 1231.020 696.390 ;
        RECT 1408.020 696.380 1411.020 696.390 ;
        RECT 1588.020 696.380 1591.020 696.390 ;
        RECT 1768.020 696.380 1771.020 696.390 ;
        RECT 1948.020 696.380 1951.020 696.390 ;
        RECT 2128.020 696.380 2131.020 696.390 ;
        RECT 2308.020 696.380 2311.020 696.390 ;
        RECT 2488.020 696.380 2491.020 696.390 ;
        RECT 2668.020 696.380 2671.020 696.390 ;
        RECT 2848.020 696.380 2851.020 696.390 ;
        RECT 2958.800 696.380 2961.800 696.390 ;
        RECT -42.180 693.380 2961.800 696.380 ;
        RECT -42.180 693.370 -39.180 693.380 ;
        RECT 148.020 693.370 151.020 693.380 ;
        RECT 328.020 693.370 331.020 693.380 ;
        RECT 508.020 693.370 511.020 693.380 ;
        RECT 688.020 693.370 691.020 693.380 ;
        RECT 868.020 693.370 871.020 693.380 ;
        RECT 1048.020 693.370 1051.020 693.380 ;
        RECT 1228.020 693.370 1231.020 693.380 ;
        RECT 1408.020 693.370 1411.020 693.380 ;
        RECT 1588.020 693.370 1591.020 693.380 ;
        RECT 1768.020 693.370 1771.020 693.380 ;
        RECT 1948.020 693.370 1951.020 693.380 ;
        RECT 2128.020 693.370 2131.020 693.380 ;
        RECT 2308.020 693.370 2311.020 693.380 ;
        RECT 2488.020 693.370 2491.020 693.380 ;
        RECT 2668.020 693.370 2671.020 693.380 ;
        RECT 2848.020 693.370 2851.020 693.380 ;
        RECT 2958.800 693.370 2961.800 693.380 ;
        RECT -42.180 516.380 -39.180 516.390 ;
        RECT 148.020 516.380 151.020 516.390 ;
        RECT 328.020 516.380 331.020 516.390 ;
        RECT 508.020 516.380 511.020 516.390 ;
        RECT 688.020 516.380 691.020 516.390 ;
        RECT 868.020 516.380 871.020 516.390 ;
        RECT 1048.020 516.380 1051.020 516.390 ;
        RECT 1228.020 516.380 1231.020 516.390 ;
        RECT 1408.020 516.380 1411.020 516.390 ;
        RECT 1588.020 516.380 1591.020 516.390 ;
        RECT 1768.020 516.380 1771.020 516.390 ;
        RECT 1948.020 516.380 1951.020 516.390 ;
        RECT 2128.020 516.380 2131.020 516.390 ;
        RECT 2308.020 516.380 2311.020 516.390 ;
        RECT 2488.020 516.380 2491.020 516.390 ;
        RECT 2668.020 516.380 2671.020 516.390 ;
        RECT 2848.020 516.380 2851.020 516.390 ;
        RECT 2958.800 516.380 2961.800 516.390 ;
        RECT -42.180 513.380 2961.800 516.380 ;
        RECT -42.180 513.370 -39.180 513.380 ;
        RECT 148.020 513.370 151.020 513.380 ;
        RECT 328.020 513.370 331.020 513.380 ;
        RECT 508.020 513.370 511.020 513.380 ;
        RECT 688.020 513.370 691.020 513.380 ;
        RECT 868.020 513.370 871.020 513.380 ;
        RECT 1048.020 513.370 1051.020 513.380 ;
        RECT 1228.020 513.370 1231.020 513.380 ;
        RECT 1408.020 513.370 1411.020 513.380 ;
        RECT 1588.020 513.370 1591.020 513.380 ;
        RECT 1768.020 513.370 1771.020 513.380 ;
        RECT 1948.020 513.370 1951.020 513.380 ;
        RECT 2128.020 513.370 2131.020 513.380 ;
        RECT 2308.020 513.370 2311.020 513.380 ;
        RECT 2488.020 513.370 2491.020 513.380 ;
        RECT 2668.020 513.370 2671.020 513.380 ;
        RECT 2848.020 513.370 2851.020 513.380 ;
        RECT 2958.800 513.370 2961.800 513.380 ;
        RECT -42.180 336.380 -39.180 336.390 ;
        RECT 148.020 336.380 151.020 336.390 ;
        RECT 328.020 336.380 331.020 336.390 ;
        RECT 508.020 336.380 511.020 336.390 ;
        RECT 688.020 336.380 691.020 336.390 ;
        RECT 868.020 336.380 871.020 336.390 ;
        RECT 1048.020 336.380 1051.020 336.390 ;
        RECT 1228.020 336.380 1231.020 336.390 ;
        RECT 1408.020 336.380 1411.020 336.390 ;
        RECT 1588.020 336.380 1591.020 336.390 ;
        RECT 1768.020 336.380 1771.020 336.390 ;
        RECT 1948.020 336.380 1951.020 336.390 ;
        RECT 2128.020 336.380 2131.020 336.390 ;
        RECT 2308.020 336.380 2311.020 336.390 ;
        RECT 2488.020 336.380 2491.020 336.390 ;
        RECT 2668.020 336.380 2671.020 336.390 ;
        RECT 2848.020 336.380 2851.020 336.390 ;
        RECT 2958.800 336.380 2961.800 336.390 ;
        RECT -42.180 333.380 2961.800 336.380 ;
        RECT -42.180 333.370 -39.180 333.380 ;
        RECT 148.020 333.370 151.020 333.380 ;
        RECT 328.020 333.370 331.020 333.380 ;
        RECT 508.020 333.370 511.020 333.380 ;
        RECT 688.020 333.370 691.020 333.380 ;
        RECT 868.020 333.370 871.020 333.380 ;
        RECT 1048.020 333.370 1051.020 333.380 ;
        RECT 1228.020 333.370 1231.020 333.380 ;
        RECT 1408.020 333.370 1411.020 333.380 ;
        RECT 1588.020 333.370 1591.020 333.380 ;
        RECT 1768.020 333.370 1771.020 333.380 ;
        RECT 1948.020 333.370 1951.020 333.380 ;
        RECT 2128.020 333.370 2131.020 333.380 ;
        RECT 2308.020 333.370 2311.020 333.380 ;
        RECT 2488.020 333.370 2491.020 333.380 ;
        RECT 2668.020 333.370 2671.020 333.380 ;
        RECT 2848.020 333.370 2851.020 333.380 ;
        RECT 2958.800 333.370 2961.800 333.380 ;
        RECT -42.180 156.380 -39.180 156.390 ;
        RECT 148.020 156.380 151.020 156.390 ;
        RECT 328.020 156.380 331.020 156.390 ;
        RECT 508.020 156.380 511.020 156.390 ;
        RECT 688.020 156.380 691.020 156.390 ;
        RECT 868.020 156.380 871.020 156.390 ;
        RECT 1048.020 156.380 1051.020 156.390 ;
        RECT 1228.020 156.380 1231.020 156.390 ;
        RECT 1408.020 156.380 1411.020 156.390 ;
        RECT 1588.020 156.380 1591.020 156.390 ;
        RECT 1768.020 156.380 1771.020 156.390 ;
        RECT 1948.020 156.380 1951.020 156.390 ;
        RECT 2128.020 156.380 2131.020 156.390 ;
        RECT 2308.020 156.380 2311.020 156.390 ;
        RECT 2488.020 156.380 2491.020 156.390 ;
        RECT 2668.020 156.380 2671.020 156.390 ;
        RECT 2848.020 156.380 2851.020 156.390 ;
        RECT 2958.800 156.380 2961.800 156.390 ;
        RECT -42.180 153.380 2961.800 156.380 ;
        RECT -42.180 153.370 -39.180 153.380 ;
        RECT 148.020 153.370 151.020 153.380 ;
        RECT 328.020 153.370 331.020 153.380 ;
        RECT 508.020 153.370 511.020 153.380 ;
        RECT 688.020 153.370 691.020 153.380 ;
        RECT 868.020 153.370 871.020 153.380 ;
        RECT 1048.020 153.370 1051.020 153.380 ;
        RECT 1228.020 153.370 1231.020 153.380 ;
        RECT 1408.020 153.370 1411.020 153.380 ;
        RECT 1588.020 153.370 1591.020 153.380 ;
        RECT 1768.020 153.370 1771.020 153.380 ;
        RECT 1948.020 153.370 1951.020 153.380 ;
        RECT 2128.020 153.370 2131.020 153.380 ;
        RECT 2308.020 153.370 2311.020 153.380 ;
        RECT 2488.020 153.370 2491.020 153.380 ;
        RECT 2668.020 153.370 2671.020 153.380 ;
        RECT 2848.020 153.370 2851.020 153.380 ;
        RECT 2958.800 153.370 2961.800 153.380 ;
        RECT -42.180 -33.820 -39.180 -33.810 ;
        RECT 148.020 -33.820 151.020 -33.810 ;
        RECT 328.020 -33.820 331.020 -33.810 ;
        RECT 508.020 -33.820 511.020 -33.810 ;
        RECT 688.020 -33.820 691.020 -33.810 ;
        RECT 868.020 -33.820 871.020 -33.810 ;
        RECT 1048.020 -33.820 1051.020 -33.810 ;
        RECT 1228.020 -33.820 1231.020 -33.810 ;
        RECT 1408.020 -33.820 1411.020 -33.810 ;
        RECT 1588.020 -33.820 1591.020 -33.810 ;
        RECT 1768.020 -33.820 1771.020 -33.810 ;
        RECT 1948.020 -33.820 1951.020 -33.810 ;
        RECT 2128.020 -33.820 2131.020 -33.810 ;
        RECT 2308.020 -33.820 2311.020 -33.810 ;
        RECT 2488.020 -33.820 2491.020 -33.810 ;
        RECT 2668.020 -33.820 2671.020 -33.810 ;
        RECT 2848.020 -33.820 2851.020 -33.810 ;
        RECT 2958.800 -33.820 2961.800 -33.810 ;
        RECT -42.180 -36.820 2961.800 -33.820 ;
        RECT -42.180 -36.830 -39.180 -36.820 ;
        RECT 148.020 -36.830 151.020 -36.820 ;
        RECT 328.020 -36.830 331.020 -36.820 ;
        RECT 508.020 -36.830 511.020 -36.820 ;
        RECT 688.020 -36.830 691.020 -36.820 ;
        RECT 868.020 -36.830 871.020 -36.820 ;
        RECT 1048.020 -36.830 1051.020 -36.820 ;
        RECT 1228.020 -36.830 1231.020 -36.820 ;
        RECT 1408.020 -36.830 1411.020 -36.820 ;
        RECT 1588.020 -36.830 1591.020 -36.820 ;
        RECT 1768.020 -36.830 1771.020 -36.820 ;
        RECT 1948.020 -36.830 1951.020 -36.820 ;
        RECT 2128.020 -36.830 2131.020 -36.820 ;
        RECT 2308.020 -36.830 2311.020 -36.820 ;
        RECT 2488.020 -36.830 2491.020 -36.820 ;
        RECT 2668.020 -36.830 2671.020 -36.820 ;
        RECT 2848.020 -36.830 2851.020 -36.820 ;
        RECT 2958.800 -36.830 2961.800 -36.820 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 855.520 1110.795 1844.060 2587.925 ;
      LAYER met1 ;
        RECT 850.990 1108.880 1847.210 2588.080 ;
      LAYER met2 ;
        RECT 1828.510 2596.000 1828.790 2600.000 ;
        RECT 1836.790 2596.000 1837.070 2600.000 ;
        RECT 1845.530 2596.000 1845.810 2600.000 ;
      LAYER met2 ;
        RECT 851.020 2595.720 853.950 2596.000 ;
        RECT 854.790 2595.720 862.230 2596.000 ;
        RECT 863.070 2595.720 870.970 2596.000 ;
        RECT 871.810 2595.720 879.250 2596.000 ;
        RECT 880.090 2595.720 887.990 2596.000 ;
        RECT 888.830 2595.720 896.270 2596.000 ;
        RECT 897.110 2595.720 905.010 2596.000 ;
        RECT 905.850 2595.720 913.750 2596.000 ;
        RECT 914.590 2595.720 922.030 2596.000 ;
        RECT 922.870 2595.720 930.770 2596.000 ;
        RECT 931.610 2595.720 939.050 2596.000 ;
        RECT 939.890 2595.720 947.790 2596.000 ;
        RECT 948.630 2595.720 956.070 2596.000 ;
        RECT 956.910 2595.720 964.810 2596.000 ;
        RECT 965.650 2595.720 973.550 2596.000 ;
        RECT 974.390 2595.720 981.830 2596.000 ;
        RECT 982.670 2595.720 990.570 2596.000 ;
        RECT 991.410 2595.720 998.850 2596.000 ;
        RECT 999.690 2595.720 1007.590 2596.000 ;
        RECT 1008.430 2595.720 1016.330 2596.000 ;
        RECT 1017.170 2595.720 1024.610 2596.000 ;
        RECT 1025.450 2595.720 1033.350 2596.000 ;
        RECT 1034.190 2595.720 1041.630 2596.000 ;
        RECT 1042.470 2595.720 1050.370 2596.000 ;
        RECT 1051.210 2595.720 1058.650 2596.000 ;
        RECT 1059.490 2595.720 1067.390 2596.000 ;
        RECT 1068.230 2595.720 1076.130 2596.000 ;
        RECT 1076.970 2595.720 1084.410 2596.000 ;
        RECT 1085.250 2595.720 1093.150 2596.000 ;
        RECT 1093.990 2595.720 1101.430 2596.000 ;
        RECT 1102.270 2595.720 1110.170 2596.000 ;
        RECT 1111.010 2595.720 1118.910 2596.000 ;
        RECT 1119.750 2595.720 1127.190 2596.000 ;
        RECT 1128.030 2595.720 1135.930 2596.000 ;
        RECT 1136.770 2595.720 1144.210 2596.000 ;
        RECT 1145.050 2595.720 1152.950 2596.000 ;
        RECT 1153.790 2595.720 1161.230 2596.000 ;
        RECT 1162.070 2595.720 1169.970 2596.000 ;
        RECT 1170.810 2595.720 1178.710 2596.000 ;
        RECT 1179.550 2595.720 1186.990 2596.000 ;
        RECT 1187.830 2595.720 1195.730 2596.000 ;
        RECT 1196.570 2595.720 1204.010 2596.000 ;
        RECT 1204.850 2595.720 1212.750 2596.000 ;
        RECT 1213.590 2595.720 1221.030 2596.000 ;
        RECT 1221.870 2595.720 1229.770 2596.000 ;
        RECT 1230.610 2595.720 1238.510 2596.000 ;
        RECT 1239.350 2595.720 1246.790 2596.000 ;
        RECT 1247.630 2595.720 1255.530 2596.000 ;
        RECT 1256.370 2595.720 1263.810 2596.000 ;
        RECT 1264.650 2595.720 1272.550 2596.000 ;
        RECT 1273.390 2595.720 1281.290 2596.000 ;
        RECT 1282.130 2595.720 1289.570 2596.000 ;
        RECT 1290.410 2595.720 1298.310 2596.000 ;
        RECT 1299.150 2595.720 1306.590 2596.000 ;
        RECT 1307.430 2595.720 1315.330 2596.000 ;
        RECT 1316.170 2595.720 1323.610 2596.000 ;
        RECT 1324.450 2595.720 1332.350 2596.000 ;
        RECT 1333.190 2595.720 1341.090 2596.000 ;
        RECT 1341.930 2595.720 1349.370 2596.000 ;
        RECT 1350.210 2595.720 1358.110 2596.000 ;
        RECT 1358.950 2595.720 1366.390 2596.000 ;
        RECT 1367.230 2595.720 1375.130 2596.000 ;
        RECT 1375.970 2595.720 1383.870 2596.000 ;
        RECT 1384.710 2595.720 1392.150 2596.000 ;
        RECT 1392.990 2595.720 1400.890 2596.000 ;
        RECT 1401.730 2595.720 1409.170 2596.000 ;
        RECT 1410.010 2595.720 1417.910 2596.000 ;
        RECT 1418.750 2595.720 1426.190 2596.000 ;
        RECT 1427.030 2595.720 1434.930 2596.000 ;
        RECT 1435.770 2595.720 1443.670 2596.000 ;
        RECT 1444.510 2595.720 1451.950 2596.000 ;
        RECT 1452.790 2595.720 1460.690 2596.000 ;
        RECT 1461.530 2595.720 1468.970 2596.000 ;
        RECT 1469.810 2595.720 1477.710 2596.000 ;
        RECT 1478.550 2595.720 1486.450 2596.000 ;
        RECT 1487.290 2595.720 1494.730 2596.000 ;
        RECT 1495.570 2595.720 1503.470 2596.000 ;
        RECT 1504.310 2595.720 1511.750 2596.000 ;
        RECT 1512.590 2595.720 1520.490 2596.000 ;
        RECT 1521.330 2595.720 1528.770 2596.000 ;
        RECT 1529.610 2595.720 1537.510 2596.000 ;
        RECT 1538.350 2595.720 1546.250 2596.000 ;
        RECT 1547.090 2595.720 1554.530 2596.000 ;
        RECT 1555.370 2595.720 1563.270 2596.000 ;
        RECT 1564.110 2595.720 1571.550 2596.000 ;
        RECT 1572.390 2595.720 1580.290 2596.000 ;
        RECT 1581.130 2595.720 1588.570 2596.000 ;
        RECT 1589.410 2595.720 1597.310 2596.000 ;
        RECT 1598.150 2595.720 1606.050 2596.000 ;
        RECT 1606.890 2595.720 1614.330 2596.000 ;
        RECT 1615.170 2595.720 1623.070 2596.000 ;
        RECT 1623.910 2595.720 1631.350 2596.000 ;
        RECT 1632.190 2595.720 1640.090 2596.000 ;
        RECT 1640.930 2595.720 1648.830 2596.000 ;
        RECT 1649.670 2595.720 1657.110 2596.000 ;
        RECT 1657.950 2595.720 1665.850 2596.000 ;
        RECT 1666.690 2595.720 1674.130 2596.000 ;
        RECT 1674.970 2595.720 1682.870 2596.000 ;
        RECT 1683.710 2595.720 1691.150 2596.000 ;
        RECT 1691.990 2595.720 1699.890 2596.000 ;
        RECT 1700.730 2595.720 1708.630 2596.000 ;
        RECT 1709.470 2595.720 1716.910 2596.000 ;
        RECT 1717.750 2595.720 1725.650 2596.000 ;
        RECT 1726.490 2595.720 1733.930 2596.000 ;
        RECT 1734.770 2595.720 1742.670 2596.000 ;
        RECT 1743.510 2595.720 1751.410 2596.000 ;
        RECT 1752.250 2595.720 1759.690 2596.000 ;
        RECT 1760.530 2595.720 1768.430 2596.000 ;
        RECT 1769.270 2595.720 1776.710 2596.000 ;
        RECT 1777.550 2595.720 1785.450 2596.000 ;
        RECT 1786.290 2595.720 1793.730 2596.000 ;
        RECT 1794.570 2595.720 1802.470 2596.000 ;
        RECT 1803.310 2595.720 1811.210 2596.000 ;
        RECT 1812.050 2595.720 1819.490 2596.000 ;
        RECT 1820.330 2595.720 1828.230 2596.000 ;
        RECT 1829.070 2595.720 1836.510 2596.000 ;
        RECT 1837.350 2595.720 1845.250 2596.000 ;
        RECT 1846.090 2595.720 1847.180 2596.000 ;
        RECT 851.020 1104.280 1847.180 2595.720 ;
        RECT 851.570 1104.000 852.570 1104.280 ;
        RECT 853.410 1104.000 854.410 1104.280 ;
        RECT 855.250 1104.000 856.710 1104.280 ;
        RECT 857.550 1104.000 858.550 1104.280 ;
        RECT 859.390 1104.000 860.850 1104.280 ;
        RECT 861.690 1104.000 862.690 1104.280 ;
        RECT 863.530 1104.000 864.990 1104.280 ;
        RECT 865.830 1104.000 866.830 1104.280 ;
        RECT 867.670 1104.000 868.670 1104.280 ;
        RECT 869.510 1104.000 870.970 1104.280 ;
        RECT 871.810 1104.000 872.810 1104.280 ;
        RECT 873.650 1104.000 875.110 1104.280 ;
        RECT 875.950 1104.000 876.950 1104.280 ;
        RECT 877.790 1104.000 879.250 1104.280 ;
        RECT 880.090 1104.000 881.090 1104.280 ;
        RECT 881.930 1104.000 882.930 1104.280 ;
        RECT 883.770 1104.000 885.230 1104.280 ;
        RECT 886.070 1104.000 887.070 1104.280 ;
        RECT 887.910 1104.000 889.370 1104.280 ;
        RECT 890.210 1104.000 891.210 1104.280 ;
        RECT 892.050 1104.000 893.510 1104.280 ;
        RECT 894.350 1104.000 895.350 1104.280 ;
        RECT 896.190 1104.000 897.650 1104.280 ;
        RECT 898.490 1104.000 899.490 1104.280 ;
        RECT 900.330 1104.000 901.330 1104.280 ;
        RECT 902.170 1104.000 903.630 1104.280 ;
        RECT 904.470 1104.000 905.470 1104.280 ;
        RECT 906.310 1104.000 907.770 1104.280 ;
        RECT 908.610 1104.000 909.610 1104.280 ;
        RECT 910.450 1104.000 911.910 1104.280 ;
        RECT 912.750 1104.000 913.750 1104.280 ;
        RECT 914.590 1104.000 915.590 1104.280 ;
        RECT 916.430 1104.000 917.890 1104.280 ;
        RECT 918.730 1104.000 919.730 1104.280 ;
        RECT 920.570 1104.000 922.030 1104.280 ;
        RECT 922.870 1104.000 923.870 1104.280 ;
        RECT 924.710 1104.000 926.170 1104.280 ;
        RECT 927.010 1104.000 928.010 1104.280 ;
        RECT 928.850 1104.000 930.310 1104.280 ;
        RECT 931.150 1104.000 932.150 1104.280 ;
        RECT 932.990 1104.000 933.990 1104.280 ;
        RECT 934.830 1104.000 936.290 1104.280 ;
        RECT 937.130 1104.000 938.130 1104.280 ;
        RECT 938.970 1104.000 940.430 1104.280 ;
        RECT 941.270 1104.000 942.270 1104.280 ;
        RECT 943.110 1104.000 944.570 1104.280 ;
        RECT 945.410 1104.000 946.410 1104.280 ;
        RECT 947.250 1104.000 948.250 1104.280 ;
        RECT 949.090 1104.000 950.550 1104.280 ;
        RECT 951.390 1104.000 952.390 1104.280 ;
        RECT 953.230 1104.000 954.690 1104.280 ;
        RECT 955.530 1104.000 956.530 1104.280 ;
        RECT 957.370 1104.000 958.830 1104.280 ;
        RECT 959.670 1104.000 960.670 1104.280 ;
        RECT 961.510 1104.000 962.970 1104.280 ;
        RECT 963.810 1104.000 964.810 1104.280 ;
        RECT 965.650 1104.000 966.650 1104.280 ;
        RECT 967.490 1104.000 968.950 1104.280 ;
        RECT 969.790 1104.000 970.790 1104.280 ;
        RECT 971.630 1104.000 973.090 1104.280 ;
        RECT 973.930 1104.000 974.930 1104.280 ;
        RECT 975.770 1104.000 977.230 1104.280 ;
        RECT 978.070 1104.000 979.070 1104.280 ;
        RECT 979.910 1104.000 980.910 1104.280 ;
        RECT 981.750 1104.000 983.210 1104.280 ;
        RECT 984.050 1104.000 985.050 1104.280 ;
        RECT 985.890 1104.000 987.350 1104.280 ;
        RECT 988.190 1104.000 989.190 1104.280 ;
        RECT 990.030 1104.000 991.490 1104.280 ;
        RECT 992.330 1104.000 993.330 1104.280 ;
        RECT 994.170 1104.000 995.630 1104.280 ;
        RECT 996.470 1104.000 997.470 1104.280 ;
        RECT 998.310 1104.000 999.310 1104.280 ;
        RECT 1000.150 1104.000 1001.610 1104.280 ;
        RECT 1002.450 1104.000 1003.450 1104.280 ;
        RECT 1004.290 1104.000 1005.750 1104.280 ;
        RECT 1006.590 1104.000 1007.590 1104.280 ;
        RECT 1008.430 1104.000 1009.890 1104.280 ;
        RECT 1010.730 1104.000 1011.730 1104.280 ;
        RECT 1012.570 1104.000 1013.570 1104.280 ;
        RECT 1014.410 1104.000 1015.870 1104.280 ;
        RECT 1016.710 1104.000 1017.710 1104.280 ;
        RECT 1018.550 1104.000 1020.010 1104.280 ;
        RECT 1020.850 1104.000 1021.850 1104.280 ;
        RECT 1022.690 1104.000 1024.150 1104.280 ;
        RECT 1024.990 1104.000 1025.990 1104.280 ;
        RECT 1026.830 1104.000 1027.830 1104.280 ;
        RECT 1028.670 1104.000 1030.130 1104.280 ;
        RECT 1030.970 1104.000 1031.970 1104.280 ;
        RECT 1032.810 1104.000 1034.270 1104.280 ;
        RECT 1035.110 1104.000 1036.110 1104.280 ;
        RECT 1036.950 1104.000 1038.410 1104.280 ;
        RECT 1039.250 1104.000 1040.250 1104.280 ;
        RECT 1041.090 1104.000 1042.550 1104.280 ;
        RECT 1043.390 1104.000 1044.390 1104.280 ;
        RECT 1045.230 1104.000 1046.230 1104.280 ;
        RECT 1047.070 1104.000 1048.530 1104.280 ;
        RECT 1049.370 1104.000 1050.370 1104.280 ;
        RECT 1051.210 1104.000 1052.670 1104.280 ;
        RECT 1053.510 1104.000 1054.510 1104.280 ;
        RECT 1055.350 1104.000 1056.810 1104.280 ;
        RECT 1057.650 1104.000 1058.650 1104.280 ;
        RECT 1059.490 1104.000 1060.490 1104.280 ;
        RECT 1061.330 1104.000 1062.790 1104.280 ;
        RECT 1063.630 1104.000 1064.630 1104.280 ;
        RECT 1065.470 1104.000 1066.930 1104.280 ;
        RECT 1067.770 1104.000 1068.770 1104.280 ;
        RECT 1069.610 1104.000 1071.070 1104.280 ;
        RECT 1071.910 1104.000 1072.910 1104.280 ;
        RECT 1073.750 1104.000 1075.210 1104.280 ;
        RECT 1076.050 1104.000 1077.050 1104.280 ;
        RECT 1077.890 1104.000 1078.890 1104.280 ;
        RECT 1079.730 1104.000 1081.190 1104.280 ;
        RECT 1082.030 1104.000 1083.030 1104.280 ;
        RECT 1083.870 1104.000 1085.330 1104.280 ;
        RECT 1086.170 1104.000 1087.170 1104.280 ;
        RECT 1088.010 1104.000 1089.470 1104.280 ;
        RECT 1090.310 1104.000 1091.310 1104.280 ;
        RECT 1092.150 1104.000 1093.150 1104.280 ;
        RECT 1093.990 1104.000 1095.450 1104.280 ;
        RECT 1096.290 1104.000 1097.290 1104.280 ;
        RECT 1098.130 1104.000 1099.590 1104.280 ;
        RECT 1100.430 1104.000 1101.430 1104.280 ;
        RECT 1102.270 1104.000 1103.730 1104.280 ;
        RECT 1104.570 1104.000 1105.570 1104.280 ;
        RECT 1106.410 1104.000 1107.870 1104.280 ;
        RECT 1108.710 1104.000 1109.710 1104.280 ;
        RECT 1110.550 1104.000 1111.550 1104.280 ;
        RECT 1112.390 1104.000 1113.850 1104.280 ;
        RECT 1114.690 1104.000 1115.690 1104.280 ;
        RECT 1116.530 1104.000 1117.990 1104.280 ;
        RECT 1118.830 1104.000 1119.830 1104.280 ;
        RECT 1120.670 1104.000 1122.130 1104.280 ;
        RECT 1122.970 1104.000 1123.970 1104.280 ;
        RECT 1124.810 1104.000 1125.810 1104.280 ;
        RECT 1126.650 1104.000 1128.110 1104.280 ;
        RECT 1128.950 1104.000 1129.950 1104.280 ;
        RECT 1130.790 1104.000 1132.250 1104.280 ;
        RECT 1133.090 1104.000 1134.090 1104.280 ;
        RECT 1134.930 1104.000 1136.390 1104.280 ;
        RECT 1137.230 1104.000 1138.230 1104.280 ;
        RECT 1139.070 1104.000 1140.530 1104.280 ;
        RECT 1141.370 1104.000 1142.370 1104.280 ;
        RECT 1143.210 1104.000 1144.210 1104.280 ;
        RECT 1145.050 1104.000 1146.510 1104.280 ;
        RECT 1147.350 1104.000 1148.350 1104.280 ;
        RECT 1149.190 1104.000 1150.650 1104.280 ;
        RECT 1151.490 1104.000 1152.490 1104.280 ;
        RECT 1153.330 1104.000 1154.790 1104.280 ;
        RECT 1155.630 1104.000 1156.630 1104.280 ;
        RECT 1157.470 1104.000 1158.470 1104.280 ;
        RECT 1159.310 1104.000 1160.770 1104.280 ;
        RECT 1161.610 1104.000 1162.610 1104.280 ;
        RECT 1163.450 1104.000 1164.910 1104.280 ;
        RECT 1165.750 1104.000 1166.750 1104.280 ;
        RECT 1167.590 1104.000 1169.050 1104.280 ;
        RECT 1169.890 1104.000 1170.890 1104.280 ;
        RECT 1171.730 1104.000 1173.190 1104.280 ;
        RECT 1174.030 1104.000 1175.030 1104.280 ;
        RECT 1175.870 1104.000 1176.870 1104.280 ;
        RECT 1177.710 1104.000 1179.170 1104.280 ;
        RECT 1180.010 1104.000 1181.010 1104.280 ;
        RECT 1181.850 1104.000 1183.310 1104.280 ;
        RECT 1184.150 1104.000 1185.150 1104.280 ;
        RECT 1185.990 1104.000 1187.450 1104.280 ;
        RECT 1188.290 1104.000 1189.290 1104.280 ;
        RECT 1190.130 1104.000 1191.130 1104.280 ;
        RECT 1191.970 1104.000 1193.430 1104.280 ;
        RECT 1194.270 1104.000 1195.270 1104.280 ;
        RECT 1196.110 1104.000 1197.570 1104.280 ;
        RECT 1198.410 1104.000 1199.410 1104.280 ;
        RECT 1200.250 1104.000 1201.710 1104.280 ;
        RECT 1202.550 1104.000 1203.550 1104.280 ;
        RECT 1204.390 1104.000 1205.390 1104.280 ;
        RECT 1206.230 1104.000 1207.690 1104.280 ;
        RECT 1208.530 1104.000 1209.530 1104.280 ;
        RECT 1210.370 1104.000 1211.830 1104.280 ;
        RECT 1212.670 1104.000 1213.670 1104.280 ;
        RECT 1214.510 1104.000 1215.970 1104.280 ;
        RECT 1216.810 1104.000 1217.810 1104.280 ;
        RECT 1218.650 1104.000 1220.110 1104.280 ;
        RECT 1220.950 1104.000 1221.950 1104.280 ;
        RECT 1222.790 1104.000 1223.790 1104.280 ;
        RECT 1224.630 1104.000 1226.090 1104.280 ;
        RECT 1226.930 1104.000 1227.930 1104.280 ;
        RECT 1228.770 1104.000 1230.230 1104.280 ;
        RECT 1231.070 1104.000 1232.070 1104.280 ;
        RECT 1232.910 1104.000 1234.370 1104.280 ;
        RECT 1235.210 1104.000 1236.210 1104.280 ;
        RECT 1237.050 1104.000 1238.050 1104.280 ;
        RECT 1238.890 1104.000 1240.350 1104.280 ;
        RECT 1241.190 1104.000 1242.190 1104.280 ;
        RECT 1243.030 1104.000 1244.490 1104.280 ;
        RECT 1245.330 1104.000 1246.330 1104.280 ;
        RECT 1247.170 1104.000 1248.630 1104.280 ;
        RECT 1249.470 1104.000 1250.470 1104.280 ;
        RECT 1251.310 1104.000 1252.770 1104.280 ;
        RECT 1253.610 1104.000 1254.610 1104.280 ;
        RECT 1255.450 1104.000 1256.450 1104.280 ;
        RECT 1257.290 1104.000 1258.750 1104.280 ;
        RECT 1259.590 1104.000 1260.590 1104.280 ;
        RECT 1261.430 1104.000 1262.890 1104.280 ;
        RECT 1263.730 1104.000 1264.730 1104.280 ;
        RECT 1265.570 1104.000 1267.030 1104.280 ;
        RECT 1267.870 1104.000 1268.870 1104.280 ;
        RECT 1269.710 1104.000 1270.710 1104.280 ;
        RECT 1271.550 1104.000 1273.010 1104.280 ;
        RECT 1273.850 1104.000 1274.850 1104.280 ;
        RECT 1275.690 1104.000 1277.150 1104.280 ;
        RECT 1277.990 1104.000 1278.990 1104.280 ;
        RECT 1279.830 1104.000 1281.290 1104.280 ;
        RECT 1282.130 1104.000 1283.130 1104.280 ;
        RECT 1283.970 1104.000 1285.430 1104.280 ;
        RECT 1286.270 1104.000 1287.270 1104.280 ;
        RECT 1288.110 1104.000 1289.110 1104.280 ;
        RECT 1289.950 1104.000 1291.410 1104.280 ;
        RECT 1292.250 1104.000 1293.250 1104.280 ;
        RECT 1294.090 1104.000 1295.550 1104.280 ;
        RECT 1296.390 1104.000 1297.390 1104.280 ;
        RECT 1298.230 1104.000 1299.690 1104.280 ;
        RECT 1300.530 1104.000 1301.530 1104.280 ;
        RECT 1302.370 1104.000 1303.370 1104.280 ;
        RECT 1304.210 1104.000 1305.670 1104.280 ;
        RECT 1306.510 1104.000 1307.510 1104.280 ;
        RECT 1308.350 1104.000 1309.810 1104.280 ;
        RECT 1310.650 1104.000 1311.650 1104.280 ;
        RECT 1312.490 1104.000 1313.950 1104.280 ;
        RECT 1314.790 1104.000 1315.790 1104.280 ;
        RECT 1316.630 1104.000 1318.090 1104.280 ;
        RECT 1318.930 1104.000 1319.930 1104.280 ;
        RECT 1320.770 1104.000 1321.770 1104.280 ;
        RECT 1322.610 1104.000 1324.070 1104.280 ;
        RECT 1324.910 1104.000 1325.910 1104.280 ;
        RECT 1326.750 1104.000 1328.210 1104.280 ;
        RECT 1329.050 1104.000 1330.050 1104.280 ;
        RECT 1330.890 1104.000 1332.350 1104.280 ;
        RECT 1333.190 1104.000 1334.190 1104.280 ;
        RECT 1335.030 1104.000 1336.030 1104.280 ;
        RECT 1336.870 1104.000 1338.330 1104.280 ;
        RECT 1339.170 1104.000 1340.170 1104.280 ;
        RECT 1341.010 1104.000 1342.470 1104.280 ;
        RECT 1343.310 1104.000 1344.310 1104.280 ;
        RECT 1345.150 1104.000 1346.610 1104.280 ;
        RECT 1347.450 1104.000 1348.450 1104.280 ;
        RECT 1349.290 1104.000 1350.750 1104.280 ;
        RECT 1351.590 1104.000 1352.590 1104.280 ;
        RECT 1353.430 1104.000 1354.430 1104.280 ;
        RECT 1355.270 1104.000 1356.730 1104.280 ;
        RECT 1357.570 1104.000 1358.570 1104.280 ;
        RECT 1359.410 1104.000 1360.870 1104.280 ;
        RECT 1361.710 1104.000 1362.710 1104.280 ;
        RECT 1363.550 1104.000 1365.010 1104.280 ;
        RECT 1365.850 1104.000 1366.850 1104.280 ;
        RECT 1367.690 1104.000 1368.690 1104.280 ;
        RECT 1369.530 1104.000 1370.990 1104.280 ;
        RECT 1371.830 1104.000 1372.830 1104.280 ;
        RECT 1373.670 1104.000 1375.130 1104.280 ;
        RECT 1375.970 1104.000 1376.970 1104.280 ;
        RECT 1377.810 1104.000 1379.270 1104.280 ;
        RECT 1380.110 1104.000 1381.110 1104.280 ;
        RECT 1381.950 1104.000 1382.950 1104.280 ;
        RECT 1383.790 1104.000 1385.250 1104.280 ;
        RECT 1386.090 1104.000 1387.090 1104.280 ;
        RECT 1387.930 1104.000 1389.390 1104.280 ;
        RECT 1390.230 1104.000 1391.230 1104.280 ;
        RECT 1392.070 1104.000 1393.530 1104.280 ;
        RECT 1394.370 1104.000 1395.370 1104.280 ;
        RECT 1396.210 1104.000 1397.670 1104.280 ;
        RECT 1398.510 1104.000 1399.510 1104.280 ;
        RECT 1400.350 1104.000 1401.350 1104.280 ;
        RECT 1402.190 1104.000 1403.650 1104.280 ;
        RECT 1404.490 1104.000 1405.490 1104.280 ;
        RECT 1406.330 1104.000 1407.790 1104.280 ;
        RECT 1408.630 1104.000 1409.630 1104.280 ;
        RECT 1410.470 1104.000 1411.930 1104.280 ;
        RECT 1412.770 1104.000 1413.770 1104.280 ;
        RECT 1414.610 1104.000 1415.610 1104.280 ;
        RECT 1416.450 1104.000 1417.910 1104.280 ;
        RECT 1418.750 1104.000 1419.750 1104.280 ;
        RECT 1420.590 1104.000 1422.050 1104.280 ;
        RECT 1422.890 1104.000 1423.890 1104.280 ;
        RECT 1424.730 1104.000 1426.190 1104.280 ;
        RECT 1427.030 1104.000 1428.030 1104.280 ;
        RECT 1428.870 1104.000 1430.330 1104.280 ;
        RECT 1431.170 1104.000 1432.170 1104.280 ;
        RECT 1433.010 1104.000 1434.010 1104.280 ;
        RECT 1434.850 1104.000 1436.310 1104.280 ;
        RECT 1437.150 1104.000 1438.150 1104.280 ;
        RECT 1438.990 1104.000 1440.450 1104.280 ;
        RECT 1441.290 1104.000 1442.290 1104.280 ;
        RECT 1443.130 1104.000 1444.590 1104.280 ;
        RECT 1445.430 1104.000 1446.430 1104.280 ;
        RECT 1447.270 1104.000 1448.270 1104.280 ;
        RECT 1449.110 1104.000 1450.570 1104.280 ;
        RECT 1451.410 1104.000 1452.410 1104.280 ;
        RECT 1453.250 1104.000 1454.710 1104.280 ;
        RECT 1455.550 1104.000 1456.550 1104.280 ;
        RECT 1457.390 1104.000 1458.850 1104.280 ;
        RECT 1459.690 1104.000 1460.690 1104.280 ;
        RECT 1461.530 1104.000 1462.990 1104.280 ;
        RECT 1463.830 1104.000 1464.830 1104.280 ;
        RECT 1465.670 1104.000 1466.670 1104.280 ;
        RECT 1467.510 1104.000 1468.970 1104.280 ;
        RECT 1469.810 1104.000 1470.810 1104.280 ;
        RECT 1471.650 1104.000 1473.110 1104.280 ;
        RECT 1473.950 1104.000 1474.950 1104.280 ;
        RECT 1475.790 1104.000 1477.250 1104.280 ;
        RECT 1478.090 1104.000 1479.090 1104.280 ;
        RECT 1479.930 1104.000 1480.930 1104.280 ;
        RECT 1481.770 1104.000 1483.230 1104.280 ;
        RECT 1484.070 1104.000 1485.070 1104.280 ;
        RECT 1485.910 1104.000 1487.370 1104.280 ;
        RECT 1488.210 1104.000 1489.210 1104.280 ;
        RECT 1490.050 1104.000 1491.510 1104.280 ;
        RECT 1492.350 1104.000 1493.350 1104.280 ;
        RECT 1494.190 1104.000 1495.650 1104.280 ;
        RECT 1496.490 1104.000 1497.490 1104.280 ;
        RECT 1498.330 1104.000 1499.330 1104.280 ;
        RECT 1500.170 1104.000 1501.630 1104.280 ;
        RECT 1502.470 1104.000 1503.470 1104.280 ;
        RECT 1504.310 1104.000 1505.770 1104.280 ;
        RECT 1506.610 1104.000 1507.610 1104.280 ;
        RECT 1508.450 1104.000 1509.910 1104.280 ;
        RECT 1510.750 1104.000 1511.750 1104.280 ;
        RECT 1512.590 1104.000 1513.590 1104.280 ;
        RECT 1514.430 1104.000 1515.890 1104.280 ;
        RECT 1516.730 1104.000 1517.730 1104.280 ;
        RECT 1518.570 1104.000 1520.030 1104.280 ;
        RECT 1520.870 1104.000 1521.870 1104.280 ;
        RECT 1522.710 1104.000 1524.170 1104.280 ;
        RECT 1525.010 1104.000 1526.010 1104.280 ;
        RECT 1526.850 1104.000 1527.850 1104.280 ;
        RECT 1528.690 1104.000 1530.150 1104.280 ;
        RECT 1530.990 1104.000 1531.990 1104.280 ;
        RECT 1532.830 1104.000 1534.290 1104.280 ;
        RECT 1535.130 1104.000 1536.130 1104.280 ;
        RECT 1536.970 1104.000 1538.430 1104.280 ;
        RECT 1539.270 1104.000 1540.270 1104.280 ;
        RECT 1541.110 1104.000 1542.570 1104.280 ;
        RECT 1543.410 1104.000 1544.410 1104.280 ;
        RECT 1545.250 1104.000 1546.250 1104.280 ;
        RECT 1547.090 1104.000 1548.550 1104.280 ;
        RECT 1549.390 1104.000 1550.390 1104.280 ;
        RECT 1551.230 1104.000 1552.690 1104.280 ;
        RECT 1553.530 1104.000 1554.530 1104.280 ;
        RECT 1555.370 1104.000 1556.830 1104.280 ;
        RECT 1557.670 1104.000 1558.670 1104.280 ;
        RECT 1559.510 1104.000 1560.510 1104.280 ;
        RECT 1561.350 1104.000 1562.810 1104.280 ;
        RECT 1563.650 1104.000 1564.650 1104.280 ;
        RECT 1565.490 1104.000 1566.950 1104.280 ;
        RECT 1567.790 1104.000 1568.790 1104.280 ;
        RECT 1569.630 1104.000 1571.090 1104.280 ;
        RECT 1571.930 1104.000 1572.930 1104.280 ;
        RECT 1573.770 1104.000 1575.230 1104.280 ;
        RECT 1576.070 1104.000 1577.070 1104.280 ;
        RECT 1577.910 1104.000 1578.910 1104.280 ;
        RECT 1579.750 1104.000 1581.210 1104.280 ;
        RECT 1582.050 1104.000 1583.050 1104.280 ;
        RECT 1583.890 1104.000 1585.350 1104.280 ;
        RECT 1586.190 1104.000 1587.190 1104.280 ;
        RECT 1588.030 1104.000 1589.490 1104.280 ;
        RECT 1590.330 1104.000 1591.330 1104.280 ;
        RECT 1592.170 1104.000 1593.170 1104.280 ;
        RECT 1594.010 1104.000 1595.470 1104.280 ;
        RECT 1596.310 1104.000 1597.310 1104.280 ;
        RECT 1598.150 1104.000 1599.610 1104.280 ;
        RECT 1600.450 1104.000 1601.450 1104.280 ;
        RECT 1602.290 1104.000 1603.750 1104.280 ;
        RECT 1604.590 1104.000 1605.590 1104.280 ;
        RECT 1606.430 1104.000 1607.890 1104.280 ;
        RECT 1608.730 1104.000 1609.730 1104.280 ;
        RECT 1610.570 1104.000 1611.570 1104.280 ;
        RECT 1612.410 1104.000 1613.870 1104.280 ;
        RECT 1614.710 1104.000 1615.710 1104.280 ;
        RECT 1616.550 1104.000 1618.010 1104.280 ;
        RECT 1618.850 1104.000 1619.850 1104.280 ;
        RECT 1620.690 1104.000 1622.150 1104.280 ;
        RECT 1622.990 1104.000 1623.990 1104.280 ;
        RECT 1624.830 1104.000 1625.830 1104.280 ;
        RECT 1626.670 1104.000 1628.130 1104.280 ;
        RECT 1628.970 1104.000 1629.970 1104.280 ;
        RECT 1630.810 1104.000 1632.270 1104.280 ;
        RECT 1633.110 1104.000 1634.110 1104.280 ;
        RECT 1634.950 1104.000 1636.410 1104.280 ;
        RECT 1637.250 1104.000 1638.250 1104.280 ;
        RECT 1639.090 1104.000 1640.550 1104.280 ;
        RECT 1641.390 1104.000 1642.390 1104.280 ;
        RECT 1643.230 1104.000 1644.230 1104.280 ;
        RECT 1645.070 1104.000 1646.530 1104.280 ;
        RECT 1647.370 1104.000 1648.370 1104.280 ;
        RECT 1649.210 1104.000 1650.670 1104.280 ;
        RECT 1651.510 1104.000 1652.510 1104.280 ;
        RECT 1653.350 1104.000 1654.810 1104.280 ;
        RECT 1655.650 1104.000 1656.650 1104.280 ;
        RECT 1657.490 1104.000 1658.490 1104.280 ;
        RECT 1659.330 1104.000 1660.790 1104.280 ;
        RECT 1661.630 1104.000 1662.630 1104.280 ;
        RECT 1663.470 1104.000 1664.930 1104.280 ;
        RECT 1665.770 1104.000 1666.770 1104.280 ;
        RECT 1667.610 1104.000 1669.070 1104.280 ;
        RECT 1669.910 1104.000 1670.910 1104.280 ;
        RECT 1671.750 1104.000 1673.210 1104.280 ;
        RECT 1674.050 1104.000 1675.050 1104.280 ;
        RECT 1675.890 1104.000 1676.890 1104.280 ;
        RECT 1677.730 1104.000 1679.190 1104.280 ;
        RECT 1680.030 1104.000 1681.030 1104.280 ;
        RECT 1681.870 1104.000 1683.330 1104.280 ;
        RECT 1684.170 1104.000 1685.170 1104.280 ;
        RECT 1686.010 1104.000 1687.470 1104.280 ;
        RECT 1688.310 1104.000 1689.310 1104.280 ;
        RECT 1690.150 1104.000 1691.150 1104.280 ;
        RECT 1691.990 1104.000 1693.450 1104.280 ;
        RECT 1694.290 1104.000 1695.290 1104.280 ;
        RECT 1696.130 1104.000 1697.590 1104.280 ;
        RECT 1698.430 1104.000 1699.430 1104.280 ;
        RECT 1700.270 1104.000 1701.730 1104.280 ;
        RECT 1702.570 1104.000 1703.570 1104.280 ;
        RECT 1704.410 1104.000 1705.410 1104.280 ;
        RECT 1706.250 1104.000 1707.710 1104.280 ;
        RECT 1708.550 1104.000 1709.550 1104.280 ;
        RECT 1710.390 1104.000 1711.850 1104.280 ;
        RECT 1712.690 1104.000 1713.690 1104.280 ;
        RECT 1714.530 1104.000 1715.990 1104.280 ;
        RECT 1716.830 1104.000 1717.830 1104.280 ;
        RECT 1718.670 1104.000 1720.130 1104.280 ;
        RECT 1720.970 1104.000 1721.970 1104.280 ;
        RECT 1722.810 1104.000 1723.810 1104.280 ;
        RECT 1724.650 1104.000 1726.110 1104.280 ;
        RECT 1726.950 1104.000 1727.950 1104.280 ;
        RECT 1728.790 1104.000 1730.250 1104.280 ;
        RECT 1731.090 1104.000 1732.090 1104.280 ;
        RECT 1732.930 1104.000 1734.390 1104.280 ;
        RECT 1735.230 1104.000 1736.230 1104.280 ;
        RECT 1737.070 1104.000 1738.070 1104.280 ;
        RECT 1738.910 1104.000 1740.370 1104.280 ;
        RECT 1741.210 1104.000 1742.210 1104.280 ;
        RECT 1743.050 1104.000 1744.510 1104.280 ;
        RECT 1745.350 1104.000 1746.350 1104.280 ;
        RECT 1747.190 1104.000 1748.650 1104.280 ;
        RECT 1749.490 1104.000 1750.490 1104.280 ;
        RECT 1751.330 1104.000 1752.790 1104.280 ;
        RECT 1753.630 1104.000 1754.630 1104.280 ;
        RECT 1755.470 1104.000 1756.470 1104.280 ;
        RECT 1757.310 1104.000 1758.770 1104.280 ;
        RECT 1759.610 1104.000 1760.610 1104.280 ;
        RECT 1761.450 1104.000 1762.910 1104.280 ;
        RECT 1763.750 1104.000 1764.750 1104.280 ;
        RECT 1765.590 1104.000 1767.050 1104.280 ;
        RECT 1767.890 1104.000 1768.890 1104.280 ;
        RECT 1769.730 1104.000 1770.730 1104.280 ;
        RECT 1771.570 1104.000 1773.030 1104.280 ;
        RECT 1773.870 1104.000 1774.870 1104.280 ;
        RECT 1775.710 1104.000 1777.170 1104.280 ;
        RECT 1778.010 1104.000 1779.010 1104.280 ;
        RECT 1779.850 1104.000 1781.310 1104.280 ;
        RECT 1782.150 1104.000 1783.150 1104.280 ;
        RECT 1783.990 1104.000 1785.450 1104.280 ;
        RECT 1786.290 1104.000 1787.290 1104.280 ;
        RECT 1788.130 1104.000 1789.130 1104.280 ;
        RECT 1789.970 1104.000 1791.430 1104.280 ;
        RECT 1792.270 1104.000 1793.270 1104.280 ;
        RECT 1794.110 1104.000 1795.570 1104.280 ;
        RECT 1796.410 1104.000 1797.410 1104.280 ;
        RECT 1798.250 1104.000 1799.710 1104.280 ;
        RECT 1800.550 1104.000 1801.550 1104.280 ;
        RECT 1802.390 1104.000 1803.390 1104.280 ;
        RECT 1804.230 1104.000 1805.690 1104.280 ;
        RECT 1806.530 1104.000 1807.530 1104.280 ;
        RECT 1808.370 1104.000 1809.830 1104.280 ;
        RECT 1810.670 1104.000 1811.670 1104.280 ;
        RECT 1812.510 1104.000 1813.970 1104.280 ;
        RECT 1814.810 1104.000 1815.810 1104.280 ;
        RECT 1816.650 1104.000 1818.110 1104.280 ;
        RECT 1818.950 1104.000 1819.950 1104.280 ;
        RECT 1820.790 1104.000 1821.790 1104.280 ;
        RECT 1822.630 1104.000 1824.090 1104.280 ;
        RECT 1824.930 1104.000 1825.930 1104.280 ;
        RECT 1826.770 1104.000 1828.230 1104.280 ;
        RECT 1829.070 1104.000 1830.070 1104.280 ;
        RECT 1830.910 1104.000 1832.370 1104.280 ;
        RECT 1833.210 1104.000 1834.210 1104.280 ;
        RECT 1835.050 1104.000 1836.050 1104.280 ;
        RECT 1836.890 1104.000 1838.350 1104.280 ;
        RECT 1839.190 1104.000 1840.190 1104.280 ;
        RECT 1841.030 1104.000 1842.490 1104.280 ;
        RECT 1843.330 1104.000 1844.330 1104.280 ;
        RECT 1845.170 1104.000 1846.630 1104.280 ;
      LAYER met3 ;
        RECT 850.000 2411.760 854.000 2412.360 ;
        RECT 850.000 2037.080 854.000 2037.680 ;
        RECT 850.000 1661.720 854.000 1662.320 ;
        RECT 850.000 1287.040 854.000 1287.640 ;
      LAYER met3 ;
        RECT 863.405 1104.255 1794.240 2588.005 ;
      LAYER met3 ;
        RECT 1846.000 1850.080 1850.000 1850.680 ;
      LAYER met4 ;
        RECT 871.040 1110.640 872.640 2588.080 ;
      LAYER met4 ;
        RECT 873.040 1110.640 904.020 2588.080 ;
        RECT 907.020 1110.640 922.020 2588.080 ;
        RECT 925.020 1110.640 940.020 2588.080 ;
        RECT 943.020 1110.640 947.440 2588.080 ;
      LAYER met4 ;
        RECT 947.840 1110.640 949.440 2588.080 ;
      LAYER met4 ;
        RECT 949.840 1110.640 958.020 2588.080 ;
        RECT 961.020 1110.640 994.020 2588.080 ;
        RECT 997.020 1110.640 1012.020 2588.080 ;
        RECT 1015.020 1110.640 1030.020 2588.080 ;
        RECT 1033.020 1110.640 1048.020 2588.080 ;
        RECT 1051.020 1110.640 1084.020 2588.080 ;
        RECT 1087.020 1110.640 1102.020 2588.080 ;
        RECT 1105.020 1110.640 1120.020 2588.080 ;
        RECT 1123.020 1110.640 1138.020 2588.080 ;
        RECT 1141.020 1110.640 1174.020 2588.080 ;
        RECT 1177.020 1110.640 1192.020 2588.080 ;
        RECT 1195.020 1110.640 1210.020 2588.080 ;
        RECT 1213.020 1110.640 1228.020 2588.080 ;
        RECT 1231.020 1110.640 1264.020 2588.080 ;
        RECT 1267.020 1110.640 1282.020 2588.080 ;
        RECT 1285.020 1110.640 1300.020 2588.080 ;
        RECT 1303.020 1110.640 1318.020 2588.080 ;
        RECT 1321.020 1110.640 1354.020 2588.080 ;
        RECT 1357.020 1110.640 1372.020 2588.080 ;
        RECT 1375.020 1110.640 1390.020 2588.080 ;
        RECT 1393.020 1110.640 1408.020 2588.080 ;
        RECT 1411.020 1110.640 1444.020 2588.080 ;
        RECT 1447.020 1110.640 1462.020 2588.080 ;
        RECT 1465.020 1110.640 1480.020 2588.080 ;
        RECT 1483.020 1110.640 1498.020 2588.080 ;
        RECT 1501.020 1110.640 1534.020 2588.080 ;
        RECT 1537.020 1110.640 1552.020 2588.080 ;
        RECT 1555.020 1110.640 1570.020 2588.080 ;
        RECT 1573.020 1110.640 1588.020 2588.080 ;
        RECT 1591.020 1110.640 1624.020 2588.080 ;
        RECT 1627.020 1110.640 1642.020 2588.080 ;
        RECT 1645.020 1110.640 1660.020 2588.080 ;
        RECT 1663.020 1110.640 1678.020 2588.080 ;
        RECT 1681.020 1110.640 1714.020 2588.080 ;
        RECT 1717.020 1110.640 1732.020 2588.080 ;
        RECT 1735.020 1110.640 1750.020 2588.080 ;
        RECT 1753.020 1110.640 1768.020 2588.080 ;
        RECT 1771.020 1110.640 1794.240 2588.080 ;
  END
END user_project_wrapper
END LIBRARY

