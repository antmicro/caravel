magic
tech sky130A
magscale 1 2
timestamp 1611670034
<< obsli1 >>
rect 1104 2159 198812 297585
<< obsm1 >>
rect 198 1300 198812 297616
<< metal2 >>
rect 846 299200 902 300000
rect 2502 299200 2558 300000
rect 4250 299200 4306 300000
rect 5998 299200 6054 300000
rect 7654 299200 7710 300000
rect 9402 299200 9458 300000
rect 11150 299200 11206 300000
rect 12898 299200 12954 300000
rect 14554 299200 14610 300000
rect 16302 299200 16358 300000
rect 18050 299200 18106 300000
rect 19798 299200 19854 300000
rect 21454 299200 21510 300000
rect 23202 299200 23258 300000
rect 24950 299200 25006 300000
rect 26698 299200 26754 300000
rect 28354 299200 28410 300000
rect 30102 299200 30158 300000
rect 31850 299200 31906 300000
rect 33598 299200 33654 300000
rect 35254 299200 35310 300000
rect 37002 299200 37058 300000
rect 38750 299200 38806 300000
rect 40498 299200 40554 300000
rect 42154 299200 42210 300000
rect 43902 299200 43958 300000
rect 45650 299200 45706 300000
rect 47398 299200 47454 300000
rect 49054 299200 49110 300000
rect 50802 299200 50858 300000
rect 52550 299200 52606 300000
rect 54206 299200 54262 300000
rect 55954 299200 56010 300000
rect 57702 299200 57758 300000
rect 59450 299200 59506 300000
rect 61106 299200 61162 300000
rect 62854 299200 62910 300000
rect 64602 299200 64658 300000
rect 66350 299200 66406 300000
rect 68006 299200 68062 300000
rect 69754 299200 69810 300000
rect 71502 299200 71558 300000
rect 73250 299200 73306 300000
rect 74906 299200 74962 300000
rect 76654 299200 76710 300000
rect 78402 299200 78458 300000
rect 80150 299200 80206 300000
rect 81806 299200 81862 300000
rect 83554 299200 83610 300000
rect 85302 299200 85358 300000
rect 87050 299200 87106 300000
rect 88706 299200 88762 300000
rect 90454 299200 90510 300000
rect 92202 299200 92258 300000
rect 93950 299200 94006 300000
rect 95606 299200 95662 300000
rect 97354 299200 97410 300000
rect 99102 299200 99158 300000
rect 100850 299200 100906 300000
rect 102506 299200 102562 300000
rect 104254 299200 104310 300000
rect 106002 299200 106058 300000
rect 107658 299200 107714 300000
rect 109406 299200 109462 300000
rect 111154 299200 111210 300000
rect 112902 299200 112958 300000
rect 114558 299200 114614 300000
rect 116306 299200 116362 300000
rect 118054 299200 118110 300000
rect 119802 299200 119858 300000
rect 121458 299200 121514 300000
rect 123206 299200 123262 300000
rect 124954 299200 125010 300000
rect 126702 299200 126758 300000
rect 128358 299200 128414 300000
rect 130106 299200 130162 300000
rect 131854 299200 131910 300000
rect 133602 299200 133658 300000
rect 135258 299200 135314 300000
rect 137006 299200 137062 300000
rect 138754 299200 138810 300000
rect 140502 299200 140558 300000
rect 142158 299200 142214 300000
rect 143906 299200 143962 300000
rect 145654 299200 145710 300000
rect 147402 299200 147458 300000
rect 149058 299200 149114 300000
rect 150806 299200 150862 300000
rect 152554 299200 152610 300000
rect 154210 299200 154266 300000
rect 155958 299200 156014 300000
rect 157706 299200 157762 300000
rect 159454 299200 159510 300000
rect 161110 299200 161166 300000
rect 162858 299200 162914 300000
rect 164606 299200 164662 300000
rect 166354 299200 166410 300000
rect 168010 299200 168066 300000
rect 169758 299200 169814 300000
rect 171506 299200 171562 300000
rect 173254 299200 173310 300000
rect 174910 299200 174966 300000
rect 176658 299200 176714 300000
rect 178406 299200 178462 300000
rect 180154 299200 180210 300000
rect 181810 299200 181866 300000
rect 183558 299200 183614 300000
rect 185306 299200 185362 300000
rect 187054 299200 187110 300000
rect 188710 299200 188766 300000
rect 190458 299200 190514 300000
rect 192206 299200 192262 300000
rect 193954 299200 194010 300000
rect 195610 299200 195666 300000
rect 197358 299200 197414 300000
rect 199106 299200 199162 300000
rect 202 0 258 800
rect 570 0 626 800
rect 938 0 994 800
rect 1398 0 1454 800
rect 1766 0 1822 800
rect 2226 0 2282 800
rect 2594 0 2650 800
rect 2962 0 3018 800
rect 3422 0 3478 800
rect 3790 0 3846 800
rect 4250 0 4306 800
rect 4618 0 4674 800
rect 5078 0 5134 800
rect 5446 0 5502 800
rect 5814 0 5870 800
rect 6274 0 6330 800
rect 6642 0 6698 800
rect 7102 0 7158 800
rect 7470 0 7526 800
rect 7838 0 7894 800
rect 8298 0 8354 800
rect 8666 0 8722 800
rect 9126 0 9182 800
rect 9494 0 9550 800
rect 9954 0 10010 800
rect 10322 0 10378 800
rect 10690 0 10746 800
rect 11150 0 11206 800
rect 11518 0 11574 800
rect 11978 0 12034 800
rect 12346 0 12402 800
rect 12714 0 12770 800
rect 13174 0 13230 800
rect 13542 0 13598 800
rect 14002 0 14058 800
rect 14370 0 14426 800
rect 14830 0 14886 800
rect 15198 0 15254 800
rect 15566 0 15622 800
rect 16026 0 16082 800
rect 16394 0 16450 800
rect 16854 0 16910 800
rect 17222 0 17278 800
rect 17682 0 17738 800
rect 18050 0 18106 800
rect 18418 0 18474 800
rect 18878 0 18934 800
rect 19246 0 19302 800
rect 19706 0 19762 800
rect 20074 0 20130 800
rect 20442 0 20498 800
rect 20902 0 20958 800
rect 21270 0 21326 800
rect 21730 0 21786 800
rect 22098 0 22154 800
rect 22558 0 22614 800
rect 22926 0 22982 800
rect 23294 0 23350 800
rect 23754 0 23810 800
rect 24122 0 24178 800
rect 24582 0 24638 800
rect 24950 0 25006 800
rect 25318 0 25374 800
rect 25778 0 25834 800
rect 26146 0 26202 800
rect 26606 0 26662 800
rect 26974 0 27030 800
rect 27434 0 27490 800
rect 27802 0 27858 800
rect 28170 0 28226 800
rect 28630 0 28686 800
rect 28998 0 29054 800
rect 29458 0 29514 800
rect 29826 0 29882 800
rect 30194 0 30250 800
rect 30654 0 30710 800
rect 31022 0 31078 800
rect 31482 0 31538 800
rect 31850 0 31906 800
rect 32310 0 32366 800
rect 32678 0 32734 800
rect 33046 0 33102 800
rect 33506 0 33562 800
rect 33874 0 33930 800
rect 34334 0 34390 800
rect 34702 0 34758 800
rect 35162 0 35218 800
rect 35530 0 35586 800
rect 35898 0 35954 800
rect 36358 0 36414 800
rect 36726 0 36782 800
rect 37186 0 37242 800
rect 37554 0 37610 800
rect 37922 0 37978 800
rect 38382 0 38438 800
rect 38750 0 38806 800
rect 39210 0 39266 800
rect 39578 0 39634 800
rect 40038 0 40094 800
rect 40406 0 40462 800
rect 40774 0 40830 800
rect 41234 0 41290 800
rect 41602 0 41658 800
rect 42062 0 42118 800
rect 42430 0 42486 800
rect 42798 0 42854 800
rect 43258 0 43314 800
rect 43626 0 43682 800
rect 44086 0 44142 800
rect 44454 0 44510 800
rect 44914 0 44970 800
rect 45282 0 45338 800
rect 45650 0 45706 800
rect 46110 0 46166 800
rect 46478 0 46534 800
rect 46938 0 46994 800
rect 47306 0 47362 800
rect 47674 0 47730 800
rect 48134 0 48190 800
rect 48502 0 48558 800
rect 48962 0 49018 800
rect 49330 0 49386 800
rect 49790 0 49846 800
rect 50158 0 50214 800
rect 50526 0 50582 800
rect 50986 0 51042 800
rect 51354 0 51410 800
rect 51814 0 51870 800
rect 52182 0 52238 800
rect 52642 0 52698 800
rect 53010 0 53066 800
rect 53378 0 53434 800
rect 53838 0 53894 800
rect 54206 0 54262 800
rect 54666 0 54722 800
rect 55034 0 55090 800
rect 55402 0 55458 800
rect 55862 0 55918 800
rect 56230 0 56286 800
rect 56690 0 56746 800
rect 57058 0 57114 800
rect 57518 0 57574 800
rect 57886 0 57942 800
rect 58254 0 58310 800
rect 58714 0 58770 800
rect 59082 0 59138 800
rect 59542 0 59598 800
rect 59910 0 59966 800
rect 60278 0 60334 800
rect 60738 0 60794 800
rect 61106 0 61162 800
rect 61566 0 61622 800
rect 61934 0 61990 800
rect 62394 0 62450 800
rect 62762 0 62818 800
rect 63130 0 63186 800
rect 63590 0 63646 800
rect 63958 0 64014 800
rect 64418 0 64474 800
rect 64786 0 64842 800
rect 65154 0 65210 800
rect 65614 0 65670 800
rect 65982 0 66038 800
rect 66442 0 66498 800
rect 66810 0 66866 800
rect 67270 0 67326 800
rect 67638 0 67694 800
rect 68006 0 68062 800
rect 68466 0 68522 800
rect 68834 0 68890 800
rect 69294 0 69350 800
rect 69662 0 69718 800
rect 70122 0 70178 800
rect 70490 0 70546 800
rect 70858 0 70914 800
rect 71318 0 71374 800
rect 71686 0 71742 800
rect 72146 0 72202 800
rect 72514 0 72570 800
rect 72882 0 72938 800
rect 73342 0 73398 800
rect 73710 0 73766 800
rect 74170 0 74226 800
rect 74538 0 74594 800
rect 74998 0 75054 800
rect 75366 0 75422 800
rect 75734 0 75790 800
rect 76194 0 76250 800
rect 76562 0 76618 800
rect 77022 0 77078 800
rect 77390 0 77446 800
rect 77758 0 77814 800
rect 78218 0 78274 800
rect 78586 0 78642 800
rect 79046 0 79102 800
rect 79414 0 79470 800
rect 79874 0 79930 800
rect 80242 0 80298 800
rect 80610 0 80666 800
rect 81070 0 81126 800
rect 81438 0 81494 800
rect 81898 0 81954 800
rect 82266 0 82322 800
rect 82634 0 82690 800
rect 83094 0 83150 800
rect 83462 0 83518 800
rect 83922 0 83978 800
rect 84290 0 84346 800
rect 84750 0 84806 800
rect 85118 0 85174 800
rect 85486 0 85542 800
rect 85946 0 86002 800
rect 86314 0 86370 800
rect 86774 0 86830 800
rect 87142 0 87198 800
rect 87602 0 87658 800
rect 87970 0 88026 800
rect 88338 0 88394 800
rect 88798 0 88854 800
rect 89166 0 89222 800
rect 89626 0 89682 800
rect 89994 0 90050 800
rect 90362 0 90418 800
rect 90822 0 90878 800
rect 91190 0 91246 800
rect 91650 0 91706 800
rect 92018 0 92074 800
rect 92478 0 92534 800
rect 92846 0 92902 800
rect 93214 0 93270 800
rect 93674 0 93730 800
rect 94042 0 94098 800
rect 94502 0 94558 800
rect 94870 0 94926 800
rect 95238 0 95294 800
rect 95698 0 95754 800
rect 96066 0 96122 800
rect 96526 0 96582 800
rect 96894 0 96950 800
rect 97354 0 97410 800
rect 97722 0 97778 800
rect 98090 0 98146 800
rect 98550 0 98606 800
rect 98918 0 98974 800
rect 99378 0 99434 800
rect 99746 0 99802 800
rect 100206 0 100262 800
rect 100574 0 100630 800
rect 100942 0 100998 800
rect 101402 0 101458 800
rect 101770 0 101826 800
rect 102230 0 102286 800
rect 102598 0 102654 800
rect 102966 0 103022 800
rect 103426 0 103482 800
rect 103794 0 103850 800
rect 104254 0 104310 800
rect 104622 0 104678 800
rect 105082 0 105138 800
rect 105450 0 105506 800
rect 105818 0 105874 800
rect 106278 0 106334 800
rect 106646 0 106702 800
rect 107106 0 107162 800
rect 107474 0 107530 800
rect 107842 0 107898 800
rect 108302 0 108358 800
rect 108670 0 108726 800
rect 109130 0 109186 800
rect 109498 0 109554 800
rect 109958 0 110014 800
rect 110326 0 110382 800
rect 110694 0 110750 800
rect 111154 0 111210 800
rect 111522 0 111578 800
rect 111982 0 112038 800
rect 112350 0 112406 800
rect 112718 0 112774 800
rect 113178 0 113234 800
rect 113546 0 113602 800
rect 114006 0 114062 800
rect 114374 0 114430 800
rect 114834 0 114890 800
rect 115202 0 115258 800
rect 115570 0 115626 800
rect 116030 0 116086 800
rect 116398 0 116454 800
rect 116858 0 116914 800
rect 117226 0 117282 800
rect 117686 0 117742 800
rect 118054 0 118110 800
rect 118422 0 118478 800
rect 118882 0 118938 800
rect 119250 0 119306 800
rect 119710 0 119766 800
rect 120078 0 120134 800
rect 120446 0 120502 800
rect 120906 0 120962 800
rect 121274 0 121330 800
rect 121734 0 121790 800
rect 122102 0 122158 800
rect 122562 0 122618 800
rect 122930 0 122986 800
rect 123298 0 123354 800
rect 123758 0 123814 800
rect 124126 0 124182 800
rect 124586 0 124642 800
rect 124954 0 125010 800
rect 125322 0 125378 800
rect 125782 0 125838 800
rect 126150 0 126206 800
rect 126610 0 126666 800
rect 126978 0 127034 800
rect 127438 0 127494 800
rect 127806 0 127862 800
rect 128174 0 128230 800
rect 128634 0 128690 800
rect 129002 0 129058 800
rect 129462 0 129518 800
rect 129830 0 129886 800
rect 130198 0 130254 800
rect 130658 0 130714 800
rect 131026 0 131082 800
rect 131486 0 131542 800
rect 131854 0 131910 800
rect 132314 0 132370 800
rect 132682 0 132738 800
rect 133050 0 133106 800
rect 133510 0 133566 800
rect 133878 0 133934 800
rect 134338 0 134394 800
rect 134706 0 134762 800
rect 135166 0 135222 800
rect 135534 0 135590 800
rect 135902 0 135958 800
rect 136362 0 136418 800
rect 136730 0 136786 800
rect 137190 0 137246 800
rect 137558 0 137614 800
rect 137926 0 137982 800
rect 138386 0 138442 800
rect 138754 0 138810 800
rect 139214 0 139270 800
rect 139582 0 139638 800
rect 140042 0 140098 800
rect 140410 0 140466 800
rect 140778 0 140834 800
rect 141238 0 141294 800
rect 141606 0 141662 800
rect 142066 0 142122 800
rect 142434 0 142490 800
rect 142802 0 142858 800
rect 143262 0 143318 800
rect 143630 0 143686 800
rect 144090 0 144146 800
rect 144458 0 144514 800
rect 144918 0 144974 800
rect 145286 0 145342 800
rect 145654 0 145710 800
rect 146114 0 146170 800
rect 146482 0 146538 800
rect 146942 0 146998 800
rect 147310 0 147366 800
rect 147678 0 147734 800
rect 148138 0 148194 800
rect 148506 0 148562 800
rect 148966 0 149022 800
rect 149334 0 149390 800
rect 149794 0 149850 800
rect 150162 0 150218 800
rect 150530 0 150586 800
rect 150990 0 151046 800
rect 151358 0 151414 800
rect 151818 0 151874 800
rect 152186 0 152242 800
rect 152646 0 152702 800
rect 153014 0 153070 800
rect 153382 0 153438 800
rect 153842 0 153898 800
rect 154210 0 154266 800
rect 154670 0 154726 800
rect 155038 0 155094 800
rect 155406 0 155462 800
rect 155866 0 155922 800
rect 156234 0 156290 800
rect 156694 0 156750 800
rect 157062 0 157118 800
rect 157522 0 157578 800
rect 157890 0 157946 800
rect 158258 0 158314 800
rect 158718 0 158774 800
rect 159086 0 159142 800
rect 159546 0 159602 800
rect 159914 0 159970 800
rect 160282 0 160338 800
rect 160742 0 160798 800
rect 161110 0 161166 800
rect 161570 0 161626 800
rect 161938 0 161994 800
rect 162398 0 162454 800
rect 162766 0 162822 800
rect 163134 0 163190 800
rect 163594 0 163650 800
rect 163962 0 164018 800
rect 164422 0 164478 800
rect 164790 0 164846 800
rect 165158 0 165214 800
rect 165618 0 165674 800
rect 165986 0 166042 800
rect 166446 0 166502 800
rect 166814 0 166870 800
rect 167274 0 167330 800
rect 167642 0 167698 800
rect 168010 0 168066 800
rect 168470 0 168526 800
rect 168838 0 168894 800
rect 169298 0 169354 800
rect 169666 0 169722 800
rect 170126 0 170182 800
rect 170494 0 170550 800
rect 170862 0 170918 800
rect 171322 0 171378 800
rect 171690 0 171746 800
rect 172150 0 172206 800
rect 172518 0 172574 800
rect 172886 0 172942 800
rect 173346 0 173402 800
rect 173714 0 173770 800
rect 174174 0 174230 800
rect 174542 0 174598 800
rect 175002 0 175058 800
rect 175370 0 175426 800
rect 175738 0 175794 800
rect 176198 0 176254 800
rect 176566 0 176622 800
rect 177026 0 177082 800
rect 177394 0 177450 800
rect 177762 0 177818 800
rect 178222 0 178278 800
rect 178590 0 178646 800
rect 179050 0 179106 800
rect 179418 0 179474 800
rect 179878 0 179934 800
rect 180246 0 180302 800
rect 180614 0 180670 800
rect 181074 0 181130 800
rect 181442 0 181498 800
rect 181902 0 181958 800
rect 182270 0 182326 800
rect 182638 0 182694 800
rect 183098 0 183154 800
rect 183466 0 183522 800
rect 183926 0 183982 800
rect 184294 0 184350 800
rect 184754 0 184810 800
rect 185122 0 185178 800
rect 185490 0 185546 800
rect 185950 0 186006 800
rect 186318 0 186374 800
rect 186778 0 186834 800
rect 187146 0 187202 800
rect 187606 0 187662 800
rect 187974 0 188030 800
rect 188342 0 188398 800
rect 188802 0 188858 800
rect 189170 0 189226 800
rect 189630 0 189686 800
rect 189998 0 190054 800
rect 190366 0 190422 800
rect 190826 0 190882 800
rect 191194 0 191250 800
rect 191654 0 191710 800
rect 192022 0 192078 800
rect 192482 0 192538 800
rect 192850 0 192906 800
rect 193218 0 193274 800
rect 193678 0 193734 800
rect 194046 0 194102 800
rect 194506 0 194562 800
rect 194874 0 194930 800
rect 195242 0 195298 800
rect 195702 0 195758 800
rect 196070 0 196126 800
rect 196530 0 196586 800
rect 196898 0 196954 800
rect 197358 0 197414 800
rect 197726 0 197782 800
rect 198094 0 198150 800
rect 198554 0 198610 800
rect 198922 0 198978 800
rect 199382 0 199438 800
rect 199750 0 199806 800
<< obsm2 >>
rect 204 299144 790 299200
rect 958 299144 2446 299200
rect 2614 299144 4194 299200
rect 4362 299144 5942 299200
rect 6110 299144 7598 299200
rect 7766 299144 9346 299200
rect 9514 299144 11094 299200
rect 11262 299144 12842 299200
rect 13010 299144 14498 299200
rect 14666 299144 16246 299200
rect 16414 299144 17994 299200
rect 18162 299144 19742 299200
rect 19910 299144 21398 299200
rect 21566 299144 23146 299200
rect 23314 299144 24894 299200
rect 25062 299144 26642 299200
rect 26810 299144 28298 299200
rect 28466 299144 30046 299200
rect 30214 299144 31794 299200
rect 31962 299144 33542 299200
rect 33710 299144 35198 299200
rect 35366 299144 36946 299200
rect 37114 299144 38694 299200
rect 38862 299144 40442 299200
rect 40610 299144 42098 299200
rect 42266 299144 43846 299200
rect 44014 299144 45594 299200
rect 45762 299144 47342 299200
rect 47510 299144 48998 299200
rect 49166 299144 50746 299200
rect 50914 299144 52494 299200
rect 52662 299144 54150 299200
rect 54318 299144 55898 299200
rect 56066 299144 57646 299200
rect 57814 299144 59394 299200
rect 59562 299144 61050 299200
rect 61218 299144 62798 299200
rect 62966 299144 64546 299200
rect 64714 299144 66294 299200
rect 66462 299144 67950 299200
rect 68118 299144 69698 299200
rect 69866 299144 71446 299200
rect 71614 299144 73194 299200
rect 73362 299144 74850 299200
rect 75018 299144 76598 299200
rect 76766 299144 78346 299200
rect 78514 299144 80094 299200
rect 80262 299144 81750 299200
rect 81918 299144 83498 299200
rect 83666 299144 85246 299200
rect 85414 299144 86994 299200
rect 87162 299144 88650 299200
rect 88818 299144 90398 299200
rect 90566 299144 92146 299200
rect 92314 299144 93894 299200
rect 94062 299144 95550 299200
rect 95718 299144 97298 299200
rect 97466 299144 99046 299200
rect 99214 299144 100794 299200
rect 100962 299144 102450 299200
rect 102618 299144 104198 299200
rect 104366 299144 105946 299200
rect 106114 299144 107602 299200
rect 107770 299144 109350 299200
rect 109518 299144 111098 299200
rect 111266 299144 112846 299200
rect 113014 299144 114502 299200
rect 114670 299144 116250 299200
rect 116418 299144 117998 299200
rect 118166 299144 119746 299200
rect 119914 299144 121402 299200
rect 121570 299144 123150 299200
rect 123318 299144 124898 299200
rect 125066 299144 126646 299200
rect 126814 299144 128302 299200
rect 128470 299144 130050 299200
rect 130218 299144 131798 299200
rect 131966 299144 133546 299200
rect 133714 299144 135202 299200
rect 135370 299144 136950 299200
rect 137118 299144 138698 299200
rect 138866 299144 140446 299200
rect 140614 299144 142102 299200
rect 142270 299144 143850 299200
rect 144018 299144 145598 299200
rect 145766 299144 147346 299200
rect 147514 299144 149002 299200
rect 149170 299144 150750 299200
rect 150918 299144 152498 299200
rect 152666 299144 154154 299200
rect 154322 299144 155902 299200
rect 156070 299144 157650 299200
rect 157818 299144 159398 299200
rect 159566 299144 161054 299200
rect 161222 299144 162802 299200
rect 162970 299144 164550 299200
rect 164718 299144 166298 299200
rect 166466 299144 167954 299200
rect 168122 299144 169702 299200
rect 169870 299144 171450 299200
rect 171618 299144 173198 299200
rect 173366 299144 174854 299200
rect 175022 299144 176602 299200
rect 176770 299144 178350 299200
rect 178518 299144 180098 299200
rect 180266 299144 181754 299200
rect 181922 299144 183502 299200
rect 183670 299144 185250 299200
rect 185418 299144 186998 299200
rect 187166 299144 188654 299200
rect 188822 299144 190402 299200
rect 190570 299144 192150 299200
rect 192318 299144 193898 299200
rect 194066 299144 195554 299200
rect 195722 299144 197302 299200
rect 197470 299144 198608 299200
rect 204 856 198608 299144
rect 314 800 514 856
rect 682 800 882 856
rect 1050 800 1342 856
rect 1510 800 1710 856
rect 1878 800 2170 856
rect 2338 800 2538 856
rect 2706 800 2906 856
rect 3074 800 3366 856
rect 3534 800 3734 856
rect 3902 800 4194 856
rect 4362 800 4562 856
rect 4730 800 5022 856
rect 5190 800 5390 856
rect 5558 800 5758 856
rect 5926 800 6218 856
rect 6386 800 6586 856
rect 6754 800 7046 856
rect 7214 800 7414 856
rect 7582 800 7782 856
rect 7950 800 8242 856
rect 8410 800 8610 856
rect 8778 800 9070 856
rect 9238 800 9438 856
rect 9606 800 9898 856
rect 10066 800 10266 856
rect 10434 800 10634 856
rect 10802 800 11094 856
rect 11262 800 11462 856
rect 11630 800 11922 856
rect 12090 800 12290 856
rect 12458 800 12658 856
rect 12826 800 13118 856
rect 13286 800 13486 856
rect 13654 800 13946 856
rect 14114 800 14314 856
rect 14482 800 14774 856
rect 14942 800 15142 856
rect 15310 800 15510 856
rect 15678 800 15970 856
rect 16138 800 16338 856
rect 16506 800 16798 856
rect 16966 800 17166 856
rect 17334 800 17626 856
rect 17794 800 17994 856
rect 18162 800 18362 856
rect 18530 800 18822 856
rect 18990 800 19190 856
rect 19358 800 19650 856
rect 19818 800 20018 856
rect 20186 800 20386 856
rect 20554 800 20846 856
rect 21014 800 21214 856
rect 21382 800 21674 856
rect 21842 800 22042 856
rect 22210 800 22502 856
rect 22670 800 22870 856
rect 23038 800 23238 856
rect 23406 800 23698 856
rect 23866 800 24066 856
rect 24234 800 24526 856
rect 24694 800 24894 856
rect 25062 800 25262 856
rect 25430 800 25722 856
rect 25890 800 26090 856
rect 26258 800 26550 856
rect 26718 800 26918 856
rect 27086 800 27378 856
rect 27546 800 27746 856
rect 27914 800 28114 856
rect 28282 800 28574 856
rect 28742 800 28942 856
rect 29110 800 29402 856
rect 29570 800 29770 856
rect 29938 800 30138 856
rect 30306 800 30598 856
rect 30766 800 30966 856
rect 31134 800 31426 856
rect 31594 800 31794 856
rect 31962 800 32254 856
rect 32422 800 32622 856
rect 32790 800 32990 856
rect 33158 800 33450 856
rect 33618 800 33818 856
rect 33986 800 34278 856
rect 34446 800 34646 856
rect 34814 800 35106 856
rect 35274 800 35474 856
rect 35642 800 35842 856
rect 36010 800 36302 856
rect 36470 800 36670 856
rect 36838 800 37130 856
rect 37298 800 37498 856
rect 37666 800 37866 856
rect 38034 800 38326 856
rect 38494 800 38694 856
rect 38862 800 39154 856
rect 39322 800 39522 856
rect 39690 800 39982 856
rect 40150 800 40350 856
rect 40518 800 40718 856
rect 40886 800 41178 856
rect 41346 800 41546 856
rect 41714 800 42006 856
rect 42174 800 42374 856
rect 42542 800 42742 856
rect 42910 800 43202 856
rect 43370 800 43570 856
rect 43738 800 44030 856
rect 44198 800 44398 856
rect 44566 800 44858 856
rect 45026 800 45226 856
rect 45394 800 45594 856
rect 45762 800 46054 856
rect 46222 800 46422 856
rect 46590 800 46882 856
rect 47050 800 47250 856
rect 47418 800 47618 856
rect 47786 800 48078 856
rect 48246 800 48446 856
rect 48614 800 48906 856
rect 49074 800 49274 856
rect 49442 800 49734 856
rect 49902 800 50102 856
rect 50270 800 50470 856
rect 50638 800 50930 856
rect 51098 800 51298 856
rect 51466 800 51758 856
rect 51926 800 52126 856
rect 52294 800 52586 856
rect 52754 800 52954 856
rect 53122 800 53322 856
rect 53490 800 53782 856
rect 53950 800 54150 856
rect 54318 800 54610 856
rect 54778 800 54978 856
rect 55146 800 55346 856
rect 55514 800 55806 856
rect 55974 800 56174 856
rect 56342 800 56634 856
rect 56802 800 57002 856
rect 57170 800 57462 856
rect 57630 800 57830 856
rect 57998 800 58198 856
rect 58366 800 58658 856
rect 58826 800 59026 856
rect 59194 800 59486 856
rect 59654 800 59854 856
rect 60022 800 60222 856
rect 60390 800 60682 856
rect 60850 800 61050 856
rect 61218 800 61510 856
rect 61678 800 61878 856
rect 62046 800 62338 856
rect 62506 800 62706 856
rect 62874 800 63074 856
rect 63242 800 63534 856
rect 63702 800 63902 856
rect 64070 800 64362 856
rect 64530 800 64730 856
rect 64898 800 65098 856
rect 65266 800 65558 856
rect 65726 800 65926 856
rect 66094 800 66386 856
rect 66554 800 66754 856
rect 66922 800 67214 856
rect 67382 800 67582 856
rect 67750 800 67950 856
rect 68118 800 68410 856
rect 68578 800 68778 856
rect 68946 800 69238 856
rect 69406 800 69606 856
rect 69774 800 70066 856
rect 70234 800 70434 856
rect 70602 800 70802 856
rect 70970 800 71262 856
rect 71430 800 71630 856
rect 71798 800 72090 856
rect 72258 800 72458 856
rect 72626 800 72826 856
rect 72994 800 73286 856
rect 73454 800 73654 856
rect 73822 800 74114 856
rect 74282 800 74482 856
rect 74650 800 74942 856
rect 75110 800 75310 856
rect 75478 800 75678 856
rect 75846 800 76138 856
rect 76306 800 76506 856
rect 76674 800 76966 856
rect 77134 800 77334 856
rect 77502 800 77702 856
rect 77870 800 78162 856
rect 78330 800 78530 856
rect 78698 800 78990 856
rect 79158 800 79358 856
rect 79526 800 79818 856
rect 79986 800 80186 856
rect 80354 800 80554 856
rect 80722 800 81014 856
rect 81182 800 81382 856
rect 81550 800 81842 856
rect 82010 800 82210 856
rect 82378 800 82578 856
rect 82746 800 83038 856
rect 83206 800 83406 856
rect 83574 800 83866 856
rect 84034 800 84234 856
rect 84402 800 84694 856
rect 84862 800 85062 856
rect 85230 800 85430 856
rect 85598 800 85890 856
rect 86058 800 86258 856
rect 86426 800 86718 856
rect 86886 800 87086 856
rect 87254 800 87546 856
rect 87714 800 87914 856
rect 88082 800 88282 856
rect 88450 800 88742 856
rect 88910 800 89110 856
rect 89278 800 89570 856
rect 89738 800 89938 856
rect 90106 800 90306 856
rect 90474 800 90766 856
rect 90934 800 91134 856
rect 91302 800 91594 856
rect 91762 800 91962 856
rect 92130 800 92422 856
rect 92590 800 92790 856
rect 92958 800 93158 856
rect 93326 800 93618 856
rect 93786 800 93986 856
rect 94154 800 94446 856
rect 94614 800 94814 856
rect 94982 800 95182 856
rect 95350 800 95642 856
rect 95810 800 96010 856
rect 96178 800 96470 856
rect 96638 800 96838 856
rect 97006 800 97298 856
rect 97466 800 97666 856
rect 97834 800 98034 856
rect 98202 800 98494 856
rect 98662 800 98862 856
rect 99030 800 99322 856
rect 99490 800 99690 856
rect 99858 800 100150 856
rect 100318 800 100518 856
rect 100686 800 100886 856
rect 101054 800 101346 856
rect 101514 800 101714 856
rect 101882 800 102174 856
rect 102342 800 102542 856
rect 102710 800 102910 856
rect 103078 800 103370 856
rect 103538 800 103738 856
rect 103906 800 104198 856
rect 104366 800 104566 856
rect 104734 800 105026 856
rect 105194 800 105394 856
rect 105562 800 105762 856
rect 105930 800 106222 856
rect 106390 800 106590 856
rect 106758 800 107050 856
rect 107218 800 107418 856
rect 107586 800 107786 856
rect 107954 800 108246 856
rect 108414 800 108614 856
rect 108782 800 109074 856
rect 109242 800 109442 856
rect 109610 800 109902 856
rect 110070 800 110270 856
rect 110438 800 110638 856
rect 110806 800 111098 856
rect 111266 800 111466 856
rect 111634 800 111926 856
rect 112094 800 112294 856
rect 112462 800 112662 856
rect 112830 800 113122 856
rect 113290 800 113490 856
rect 113658 800 113950 856
rect 114118 800 114318 856
rect 114486 800 114778 856
rect 114946 800 115146 856
rect 115314 800 115514 856
rect 115682 800 115974 856
rect 116142 800 116342 856
rect 116510 800 116802 856
rect 116970 800 117170 856
rect 117338 800 117630 856
rect 117798 800 117998 856
rect 118166 800 118366 856
rect 118534 800 118826 856
rect 118994 800 119194 856
rect 119362 800 119654 856
rect 119822 800 120022 856
rect 120190 800 120390 856
rect 120558 800 120850 856
rect 121018 800 121218 856
rect 121386 800 121678 856
rect 121846 800 122046 856
rect 122214 800 122506 856
rect 122674 800 122874 856
rect 123042 800 123242 856
rect 123410 800 123702 856
rect 123870 800 124070 856
rect 124238 800 124530 856
rect 124698 800 124898 856
rect 125066 800 125266 856
rect 125434 800 125726 856
rect 125894 800 126094 856
rect 126262 800 126554 856
rect 126722 800 126922 856
rect 127090 800 127382 856
rect 127550 800 127750 856
rect 127918 800 128118 856
rect 128286 800 128578 856
rect 128746 800 128946 856
rect 129114 800 129406 856
rect 129574 800 129774 856
rect 129942 800 130142 856
rect 130310 800 130602 856
rect 130770 800 130970 856
rect 131138 800 131430 856
rect 131598 800 131798 856
rect 131966 800 132258 856
rect 132426 800 132626 856
rect 132794 800 132994 856
rect 133162 800 133454 856
rect 133622 800 133822 856
rect 133990 800 134282 856
rect 134450 800 134650 856
rect 134818 800 135110 856
rect 135278 800 135478 856
rect 135646 800 135846 856
rect 136014 800 136306 856
rect 136474 800 136674 856
rect 136842 800 137134 856
rect 137302 800 137502 856
rect 137670 800 137870 856
rect 138038 800 138330 856
rect 138498 800 138698 856
rect 138866 800 139158 856
rect 139326 800 139526 856
rect 139694 800 139986 856
rect 140154 800 140354 856
rect 140522 800 140722 856
rect 140890 800 141182 856
rect 141350 800 141550 856
rect 141718 800 142010 856
rect 142178 800 142378 856
rect 142546 800 142746 856
rect 142914 800 143206 856
rect 143374 800 143574 856
rect 143742 800 144034 856
rect 144202 800 144402 856
rect 144570 800 144862 856
rect 145030 800 145230 856
rect 145398 800 145598 856
rect 145766 800 146058 856
rect 146226 800 146426 856
rect 146594 800 146886 856
rect 147054 800 147254 856
rect 147422 800 147622 856
rect 147790 800 148082 856
rect 148250 800 148450 856
rect 148618 800 148910 856
rect 149078 800 149278 856
rect 149446 800 149738 856
rect 149906 800 150106 856
rect 150274 800 150474 856
rect 150642 800 150934 856
rect 151102 800 151302 856
rect 151470 800 151762 856
rect 151930 800 152130 856
rect 152298 800 152590 856
rect 152758 800 152958 856
rect 153126 800 153326 856
rect 153494 800 153786 856
rect 153954 800 154154 856
rect 154322 800 154614 856
rect 154782 800 154982 856
rect 155150 800 155350 856
rect 155518 800 155810 856
rect 155978 800 156178 856
rect 156346 800 156638 856
rect 156806 800 157006 856
rect 157174 800 157466 856
rect 157634 800 157834 856
rect 158002 800 158202 856
rect 158370 800 158662 856
rect 158830 800 159030 856
rect 159198 800 159490 856
rect 159658 800 159858 856
rect 160026 800 160226 856
rect 160394 800 160686 856
rect 160854 800 161054 856
rect 161222 800 161514 856
rect 161682 800 161882 856
rect 162050 800 162342 856
rect 162510 800 162710 856
rect 162878 800 163078 856
rect 163246 800 163538 856
rect 163706 800 163906 856
rect 164074 800 164366 856
rect 164534 800 164734 856
rect 164902 800 165102 856
rect 165270 800 165562 856
rect 165730 800 165930 856
rect 166098 800 166390 856
rect 166558 800 166758 856
rect 166926 800 167218 856
rect 167386 800 167586 856
rect 167754 800 167954 856
rect 168122 800 168414 856
rect 168582 800 168782 856
rect 168950 800 169242 856
rect 169410 800 169610 856
rect 169778 800 170070 856
rect 170238 800 170438 856
rect 170606 800 170806 856
rect 170974 800 171266 856
rect 171434 800 171634 856
rect 171802 800 172094 856
rect 172262 800 172462 856
rect 172630 800 172830 856
rect 172998 800 173290 856
rect 173458 800 173658 856
rect 173826 800 174118 856
rect 174286 800 174486 856
rect 174654 800 174946 856
rect 175114 800 175314 856
rect 175482 800 175682 856
rect 175850 800 176142 856
rect 176310 800 176510 856
rect 176678 800 176970 856
rect 177138 800 177338 856
rect 177506 800 177706 856
rect 177874 800 178166 856
rect 178334 800 178534 856
rect 178702 800 178994 856
rect 179162 800 179362 856
rect 179530 800 179822 856
rect 179990 800 180190 856
rect 180358 800 180558 856
rect 180726 800 181018 856
rect 181186 800 181386 856
rect 181554 800 181846 856
rect 182014 800 182214 856
rect 182382 800 182582 856
rect 182750 800 183042 856
rect 183210 800 183410 856
rect 183578 800 183870 856
rect 184038 800 184238 856
rect 184406 800 184698 856
rect 184866 800 185066 856
rect 185234 800 185434 856
rect 185602 800 185894 856
rect 186062 800 186262 856
rect 186430 800 186722 856
rect 186890 800 187090 856
rect 187258 800 187550 856
rect 187718 800 187918 856
rect 188086 800 188286 856
rect 188454 800 188746 856
rect 188914 800 189114 856
rect 189282 800 189574 856
rect 189742 800 189942 856
rect 190110 800 190310 856
rect 190478 800 190770 856
rect 190938 800 191138 856
rect 191306 800 191598 856
rect 191766 800 191966 856
rect 192134 800 192426 856
rect 192594 800 192794 856
rect 192962 800 193162 856
rect 193330 800 193622 856
rect 193790 800 193990 856
rect 194158 800 194450 856
rect 194618 800 194818 856
rect 194986 800 195186 856
rect 195354 800 195646 856
rect 195814 800 196014 856
rect 196182 800 196474 856
rect 196642 800 196842 856
rect 197010 800 197302 856
rect 197470 800 197670 856
rect 197838 800 198038 856
rect 198206 800 198498 856
<< metal3 >>
rect 0 224952 800 225072
rect 0 74944 800 75064
rect 199200 224952 200000 225072
rect 199200 74944 200000 75064
<< obsm3 >>
rect 2405 851 188848 297601
<< metal4 >>
rect 4208 2128 4528 297616
rect 19568 2128 19888 297616
rect 34928 2128 35248 297616
rect 50288 2128 50608 297616
rect 65648 2128 65968 297616
rect 81008 2128 81328 297616
rect 96368 2128 96688 297616
rect 111728 2128 112048 297616
rect 127088 2128 127408 297616
rect 142448 2128 142768 297616
rect 157808 2128 158128 297616
rect 173168 2128 173488 297616
rect 188528 2128 188848 297616
<< obsm4 >>
rect 3187 4251 4128 293997
rect 4608 4251 19488 293997
rect 19968 4251 34848 293997
rect 35328 4251 50208 293997
rect 50688 4251 65568 293997
rect 66048 4251 80928 293997
rect 81408 4251 96288 293997
rect 96768 4251 111648 293997
rect 112128 4251 127008 293997
rect 127488 4251 139413 293997
<< labels >>
rlabel metal2 s 846 299200 902 300000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 52550 299200 52606 300000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 57702 299200 57758 300000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 62854 299200 62910 300000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 68006 299200 68062 300000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 73250 299200 73306 300000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 78402 299200 78458 300000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 83554 299200 83610 300000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 88706 299200 88762 300000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 93950 299200 94006 300000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 99102 299200 99158 300000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 5998 299200 6054 300000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 104254 299200 104310 300000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 109406 299200 109462 300000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 114558 299200 114614 300000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 119802 299200 119858 300000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 124954 299200 125010 300000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 130106 299200 130162 300000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 135258 299200 135314 300000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 140502 299200 140558 300000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 145654 299200 145710 300000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 150806 299200 150862 300000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 11150 299200 11206 300000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 155958 299200 156014 300000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 161110 299200 161166 300000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 166354 299200 166410 300000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 171506 299200 171562 300000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 176658 299200 176714 300000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 181810 299200 181866 300000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 187054 299200 187110 300000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 192206 299200 192262 300000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 16302 299200 16358 300000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 21454 299200 21510 300000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 26698 299200 26754 300000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 31850 299200 31906 300000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 37002 299200 37058 300000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 42154 299200 42210 300000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 47398 299200 47454 300000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 2502 299200 2558 300000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 54206 299200 54262 300000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 59450 299200 59506 300000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 64602 299200 64658 300000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 69754 299200 69810 300000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 74906 299200 74962 300000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 80150 299200 80206 300000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 85302 299200 85358 300000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 90454 299200 90510 300000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 95606 299200 95662 300000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 100850 299200 100906 300000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 7654 299200 7710 300000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 106002 299200 106058 300000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 111154 299200 111210 300000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 116306 299200 116362 300000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 121458 299200 121514 300000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 126702 299200 126758 300000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 131854 299200 131910 300000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 137006 299200 137062 300000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 142158 299200 142214 300000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 147402 299200 147458 300000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 152554 299200 152610 300000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 12898 299200 12954 300000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 157706 299200 157762 300000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 162858 299200 162914 300000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 168010 299200 168066 300000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 173254 299200 173310 300000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 178406 299200 178462 300000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 183558 299200 183614 300000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 188710 299200 188766 300000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 193954 299200 194010 300000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 18050 299200 18106 300000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 23202 299200 23258 300000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 28354 299200 28410 300000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 33598 299200 33654 300000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 38750 299200 38806 300000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 43902 299200 43958 300000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 49054 299200 49110 300000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 4250 299200 4306 300000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 55954 299200 56010 300000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 61106 299200 61162 300000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 66350 299200 66406 300000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 71502 299200 71558 300000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 76654 299200 76710 300000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 81806 299200 81862 300000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 87050 299200 87106 300000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 92202 299200 92258 300000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 97354 299200 97410 300000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 102506 299200 102562 300000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 9402 299200 9458 300000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 107658 299200 107714 300000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 112902 299200 112958 300000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 118054 299200 118110 300000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 123206 299200 123262 300000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 128358 299200 128414 300000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 133602 299200 133658 300000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 138754 299200 138810 300000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 143906 299200 143962 300000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 149058 299200 149114 300000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 154210 299200 154266 300000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 14554 299200 14610 300000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 159454 299200 159510 300000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 164606 299200 164662 300000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 169758 299200 169814 300000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 174910 299200 174966 300000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 180154 299200 180210 300000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 185306 299200 185362 300000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 190458 299200 190514 300000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 195610 299200 195666 300000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 19798 299200 19854 300000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 24950 299200 25006 300000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 30102 299200 30158 300000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 35254 299200 35310 300000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 40498 299200 40554 300000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 45650 299200 45706 300000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 50802 299200 50858 300000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 43258 0 43314 800 6 la_data_in[0]
port 115 nsew signal input
rlabel metal2 s 165158 0 165214 800 6 la_data_in[100]
port 116 nsew signal input
rlabel metal2 s 166446 0 166502 800 6 la_data_in[101]
port 117 nsew signal input
rlabel metal2 s 167642 0 167698 800 6 la_data_in[102]
port 118 nsew signal input
rlabel metal2 s 168838 0 168894 800 6 la_data_in[103]
port 119 nsew signal input
rlabel metal2 s 170126 0 170182 800 6 la_data_in[104]
port 120 nsew signal input
rlabel metal2 s 171322 0 171378 800 6 la_data_in[105]
port 121 nsew signal input
rlabel metal2 s 172518 0 172574 800 6 la_data_in[106]
port 122 nsew signal input
rlabel metal2 s 173714 0 173770 800 6 la_data_in[107]
port 123 nsew signal input
rlabel metal2 s 175002 0 175058 800 6 la_data_in[108]
port 124 nsew signal input
rlabel metal2 s 176198 0 176254 800 6 la_data_in[109]
port 125 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 la_data_in[10]
port 126 nsew signal input
rlabel metal2 s 177394 0 177450 800 6 la_data_in[110]
port 127 nsew signal input
rlabel metal2 s 178590 0 178646 800 6 la_data_in[111]
port 128 nsew signal input
rlabel metal2 s 179878 0 179934 800 6 la_data_in[112]
port 129 nsew signal input
rlabel metal2 s 181074 0 181130 800 6 la_data_in[113]
port 130 nsew signal input
rlabel metal2 s 182270 0 182326 800 6 la_data_in[114]
port 131 nsew signal input
rlabel metal2 s 183466 0 183522 800 6 la_data_in[115]
port 132 nsew signal input
rlabel metal2 s 184754 0 184810 800 6 la_data_in[116]
port 133 nsew signal input
rlabel metal2 s 185950 0 186006 800 6 la_data_in[117]
port 134 nsew signal input
rlabel metal2 s 187146 0 187202 800 6 la_data_in[118]
port 135 nsew signal input
rlabel metal2 s 188342 0 188398 800 6 la_data_in[119]
port 136 nsew signal input
rlabel metal2 s 56690 0 56746 800 6 la_data_in[11]
port 137 nsew signal input
rlabel metal2 s 189630 0 189686 800 6 la_data_in[120]
port 138 nsew signal input
rlabel metal2 s 190826 0 190882 800 6 la_data_in[121]
port 139 nsew signal input
rlabel metal2 s 192022 0 192078 800 6 la_data_in[122]
port 140 nsew signal input
rlabel metal2 s 193218 0 193274 800 6 la_data_in[123]
port 141 nsew signal input
rlabel metal2 s 194506 0 194562 800 6 la_data_in[124]
port 142 nsew signal input
rlabel metal2 s 195702 0 195758 800 6 la_data_in[125]
port 143 nsew signal input
rlabel metal2 s 196898 0 196954 800 6 la_data_in[126]
port 144 nsew signal input
rlabel metal2 s 198094 0 198150 800 6 la_data_in[127]
port 145 nsew signal input
rlabel metal2 s 57886 0 57942 800 6 la_data_in[12]
port 146 nsew signal input
rlabel metal2 s 59082 0 59138 800 6 la_data_in[13]
port 147 nsew signal input
rlabel metal2 s 60278 0 60334 800 6 la_data_in[14]
port 148 nsew signal input
rlabel metal2 s 61566 0 61622 800 6 la_data_in[15]
port 149 nsew signal input
rlabel metal2 s 62762 0 62818 800 6 la_data_in[16]
port 150 nsew signal input
rlabel metal2 s 63958 0 64014 800 6 la_data_in[17]
port 151 nsew signal input
rlabel metal2 s 65154 0 65210 800 6 la_data_in[18]
port 152 nsew signal input
rlabel metal2 s 66442 0 66498 800 6 la_data_in[19]
port 153 nsew signal input
rlabel metal2 s 44454 0 44510 800 6 la_data_in[1]
port 154 nsew signal input
rlabel metal2 s 67638 0 67694 800 6 la_data_in[20]
port 155 nsew signal input
rlabel metal2 s 68834 0 68890 800 6 la_data_in[21]
port 156 nsew signal input
rlabel metal2 s 70122 0 70178 800 6 la_data_in[22]
port 157 nsew signal input
rlabel metal2 s 71318 0 71374 800 6 la_data_in[23]
port 158 nsew signal input
rlabel metal2 s 72514 0 72570 800 6 la_data_in[24]
port 159 nsew signal input
rlabel metal2 s 73710 0 73766 800 6 la_data_in[25]
port 160 nsew signal input
rlabel metal2 s 74998 0 75054 800 6 la_data_in[26]
port 161 nsew signal input
rlabel metal2 s 76194 0 76250 800 6 la_data_in[27]
port 162 nsew signal input
rlabel metal2 s 77390 0 77446 800 6 la_data_in[28]
port 163 nsew signal input
rlabel metal2 s 78586 0 78642 800 6 la_data_in[29]
port 164 nsew signal input
rlabel metal2 s 45650 0 45706 800 6 la_data_in[2]
port 165 nsew signal input
rlabel metal2 s 79874 0 79930 800 6 la_data_in[30]
port 166 nsew signal input
rlabel metal2 s 81070 0 81126 800 6 la_data_in[31]
port 167 nsew signal input
rlabel metal2 s 82266 0 82322 800 6 la_data_in[32]
port 168 nsew signal input
rlabel metal2 s 83462 0 83518 800 6 la_data_in[33]
port 169 nsew signal input
rlabel metal2 s 84750 0 84806 800 6 la_data_in[34]
port 170 nsew signal input
rlabel metal2 s 85946 0 86002 800 6 la_data_in[35]
port 171 nsew signal input
rlabel metal2 s 87142 0 87198 800 6 la_data_in[36]
port 172 nsew signal input
rlabel metal2 s 88338 0 88394 800 6 la_data_in[37]
port 173 nsew signal input
rlabel metal2 s 89626 0 89682 800 6 la_data_in[38]
port 174 nsew signal input
rlabel metal2 s 90822 0 90878 800 6 la_data_in[39]
port 175 nsew signal input
rlabel metal2 s 46938 0 46994 800 6 la_data_in[3]
port 176 nsew signal input
rlabel metal2 s 92018 0 92074 800 6 la_data_in[40]
port 177 nsew signal input
rlabel metal2 s 93214 0 93270 800 6 la_data_in[41]
port 178 nsew signal input
rlabel metal2 s 94502 0 94558 800 6 la_data_in[42]
port 179 nsew signal input
rlabel metal2 s 95698 0 95754 800 6 la_data_in[43]
port 180 nsew signal input
rlabel metal2 s 96894 0 96950 800 6 la_data_in[44]
port 181 nsew signal input
rlabel metal2 s 98090 0 98146 800 6 la_data_in[45]
port 182 nsew signal input
rlabel metal2 s 99378 0 99434 800 6 la_data_in[46]
port 183 nsew signal input
rlabel metal2 s 100574 0 100630 800 6 la_data_in[47]
port 184 nsew signal input
rlabel metal2 s 101770 0 101826 800 6 la_data_in[48]
port 185 nsew signal input
rlabel metal2 s 102966 0 103022 800 6 la_data_in[49]
port 186 nsew signal input
rlabel metal2 s 48134 0 48190 800 6 la_data_in[4]
port 187 nsew signal input
rlabel metal2 s 104254 0 104310 800 6 la_data_in[50]
port 188 nsew signal input
rlabel metal2 s 105450 0 105506 800 6 la_data_in[51]
port 189 nsew signal input
rlabel metal2 s 106646 0 106702 800 6 la_data_in[52]
port 190 nsew signal input
rlabel metal2 s 107842 0 107898 800 6 la_data_in[53]
port 191 nsew signal input
rlabel metal2 s 109130 0 109186 800 6 la_data_in[54]
port 192 nsew signal input
rlabel metal2 s 110326 0 110382 800 6 la_data_in[55]
port 193 nsew signal input
rlabel metal2 s 111522 0 111578 800 6 la_data_in[56]
port 194 nsew signal input
rlabel metal2 s 112718 0 112774 800 6 la_data_in[57]
port 195 nsew signal input
rlabel metal2 s 114006 0 114062 800 6 la_data_in[58]
port 196 nsew signal input
rlabel metal2 s 115202 0 115258 800 6 la_data_in[59]
port 197 nsew signal input
rlabel metal2 s 49330 0 49386 800 6 la_data_in[5]
port 198 nsew signal input
rlabel metal2 s 116398 0 116454 800 6 la_data_in[60]
port 199 nsew signal input
rlabel metal2 s 117686 0 117742 800 6 la_data_in[61]
port 200 nsew signal input
rlabel metal2 s 118882 0 118938 800 6 la_data_in[62]
port 201 nsew signal input
rlabel metal2 s 120078 0 120134 800 6 la_data_in[63]
port 202 nsew signal input
rlabel metal2 s 121274 0 121330 800 6 la_data_in[64]
port 203 nsew signal input
rlabel metal2 s 122562 0 122618 800 6 la_data_in[65]
port 204 nsew signal input
rlabel metal2 s 123758 0 123814 800 6 la_data_in[66]
port 205 nsew signal input
rlabel metal2 s 124954 0 125010 800 6 la_data_in[67]
port 206 nsew signal input
rlabel metal2 s 126150 0 126206 800 6 la_data_in[68]
port 207 nsew signal input
rlabel metal2 s 127438 0 127494 800 6 la_data_in[69]
port 208 nsew signal input
rlabel metal2 s 50526 0 50582 800 6 la_data_in[6]
port 209 nsew signal input
rlabel metal2 s 128634 0 128690 800 6 la_data_in[70]
port 210 nsew signal input
rlabel metal2 s 129830 0 129886 800 6 la_data_in[71]
port 211 nsew signal input
rlabel metal2 s 131026 0 131082 800 6 la_data_in[72]
port 212 nsew signal input
rlabel metal2 s 132314 0 132370 800 6 la_data_in[73]
port 213 nsew signal input
rlabel metal2 s 133510 0 133566 800 6 la_data_in[74]
port 214 nsew signal input
rlabel metal2 s 134706 0 134762 800 6 la_data_in[75]
port 215 nsew signal input
rlabel metal2 s 135902 0 135958 800 6 la_data_in[76]
port 216 nsew signal input
rlabel metal2 s 137190 0 137246 800 6 la_data_in[77]
port 217 nsew signal input
rlabel metal2 s 138386 0 138442 800 6 la_data_in[78]
port 218 nsew signal input
rlabel metal2 s 139582 0 139638 800 6 la_data_in[79]
port 219 nsew signal input
rlabel metal2 s 51814 0 51870 800 6 la_data_in[7]
port 220 nsew signal input
rlabel metal2 s 140778 0 140834 800 6 la_data_in[80]
port 221 nsew signal input
rlabel metal2 s 142066 0 142122 800 6 la_data_in[81]
port 222 nsew signal input
rlabel metal2 s 143262 0 143318 800 6 la_data_in[82]
port 223 nsew signal input
rlabel metal2 s 144458 0 144514 800 6 la_data_in[83]
port 224 nsew signal input
rlabel metal2 s 145654 0 145710 800 6 la_data_in[84]
port 225 nsew signal input
rlabel metal2 s 146942 0 146998 800 6 la_data_in[85]
port 226 nsew signal input
rlabel metal2 s 148138 0 148194 800 6 la_data_in[86]
port 227 nsew signal input
rlabel metal2 s 149334 0 149390 800 6 la_data_in[87]
port 228 nsew signal input
rlabel metal2 s 150530 0 150586 800 6 la_data_in[88]
port 229 nsew signal input
rlabel metal2 s 151818 0 151874 800 6 la_data_in[89]
port 230 nsew signal input
rlabel metal2 s 53010 0 53066 800 6 la_data_in[8]
port 231 nsew signal input
rlabel metal2 s 153014 0 153070 800 6 la_data_in[90]
port 232 nsew signal input
rlabel metal2 s 154210 0 154266 800 6 la_data_in[91]
port 233 nsew signal input
rlabel metal2 s 155406 0 155462 800 6 la_data_in[92]
port 234 nsew signal input
rlabel metal2 s 156694 0 156750 800 6 la_data_in[93]
port 235 nsew signal input
rlabel metal2 s 157890 0 157946 800 6 la_data_in[94]
port 236 nsew signal input
rlabel metal2 s 159086 0 159142 800 6 la_data_in[95]
port 237 nsew signal input
rlabel metal2 s 160282 0 160338 800 6 la_data_in[96]
port 238 nsew signal input
rlabel metal2 s 161570 0 161626 800 6 la_data_in[97]
port 239 nsew signal input
rlabel metal2 s 162766 0 162822 800 6 la_data_in[98]
port 240 nsew signal input
rlabel metal2 s 163962 0 164018 800 6 la_data_in[99]
port 241 nsew signal input
rlabel metal2 s 54206 0 54262 800 6 la_data_in[9]
port 242 nsew signal input
rlabel metal2 s 43626 0 43682 800 6 la_data_out[0]
port 243 nsew signal output
rlabel metal2 s 165618 0 165674 800 6 la_data_out[100]
port 244 nsew signal output
rlabel metal2 s 166814 0 166870 800 6 la_data_out[101]
port 245 nsew signal output
rlabel metal2 s 168010 0 168066 800 6 la_data_out[102]
port 246 nsew signal output
rlabel metal2 s 169298 0 169354 800 6 la_data_out[103]
port 247 nsew signal output
rlabel metal2 s 170494 0 170550 800 6 la_data_out[104]
port 248 nsew signal output
rlabel metal2 s 171690 0 171746 800 6 la_data_out[105]
port 249 nsew signal output
rlabel metal2 s 172886 0 172942 800 6 la_data_out[106]
port 250 nsew signal output
rlabel metal2 s 174174 0 174230 800 6 la_data_out[107]
port 251 nsew signal output
rlabel metal2 s 175370 0 175426 800 6 la_data_out[108]
port 252 nsew signal output
rlabel metal2 s 176566 0 176622 800 6 la_data_out[109]
port 253 nsew signal output
rlabel metal2 s 55862 0 55918 800 6 la_data_out[10]
port 254 nsew signal output
rlabel metal2 s 177762 0 177818 800 6 la_data_out[110]
port 255 nsew signal output
rlabel metal2 s 179050 0 179106 800 6 la_data_out[111]
port 256 nsew signal output
rlabel metal2 s 180246 0 180302 800 6 la_data_out[112]
port 257 nsew signal output
rlabel metal2 s 181442 0 181498 800 6 la_data_out[113]
port 258 nsew signal output
rlabel metal2 s 182638 0 182694 800 6 la_data_out[114]
port 259 nsew signal output
rlabel metal2 s 183926 0 183982 800 6 la_data_out[115]
port 260 nsew signal output
rlabel metal2 s 185122 0 185178 800 6 la_data_out[116]
port 261 nsew signal output
rlabel metal2 s 186318 0 186374 800 6 la_data_out[117]
port 262 nsew signal output
rlabel metal2 s 187606 0 187662 800 6 la_data_out[118]
port 263 nsew signal output
rlabel metal2 s 188802 0 188858 800 6 la_data_out[119]
port 264 nsew signal output
rlabel metal2 s 57058 0 57114 800 6 la_data_out[11]
port 265 nsew signal output
rlabel metal2 s 189998 0 190054 800 6 la_data_out[120]
port 266 nsew signal output
rlabel metal2 s 191194 0 191250 800 6 la_data_out[121]
port 267 nsew signal output
rlabel metal2 s 192482 0 192538 800 6 la_data_out[122]
port 268 nsew signal output
rlabel metal2 s 193678 0 193734 800 6 la_data_out[123]
port 269 nsew signal output
rlabel metal2 s 194874 0 194930 800 6 la_data_out[124]
port 270 nsew signal output
rlabel metal2 s 196070 0 196126 800 6 la_data_out[125]
port 271 nsew signal output
rlabel metal2 s 197358 0 197414 800 6 la_data_out[126]
port 272 nsew signal output
rlabel metal2 s 198554 0 198610 800 6 la_data_out[127]
port 273 nsew signal output
rlabel metal2 s 58254 0 58310 800 6 la_data_out[12]
port 274 nsew signal output
rlabel metal2 s 59542 0 59598 800 6 la_data_out[13]
port 275 nsew signal output
rlabel metal2 s 60738 0 60794 800 6 la_data_out[14]
port 276 nsew signal output
rlabel metal2 s 61934 0 61990 800 6 la_data_out[15]
port 277 nsew signal output
rlabel metal2 s 63130 0 63186 800 6 la_data_out[16]
port 278 nsew signal output
rlabel metal2 s 64418 0 64474 800 6 la_data_out[17]
port 279 nsew signal output
rlabel metal2 s 65614 0 65670 800 6 la_data_out[18]
port 280 nsew signal output
rlabel metal2 s 66810 0 66866 800 6 la_data_out[19]
port 281 nsew signal output
rlabel metal2 s 44914 0 44970 800 6 la_data_out[1]
port 282 nsew signal output
rlabel metal2 s 68006 0 68062 800 6 la_data_out[20]
port 283 nsew signal output
rlabel metal2 s 69294 0 69350 800 6 la_data_out[21]
port 284 nsew signal output
rlabel metal2 s 70490 0 70546 800 6 la_data_out[22]
port 285 nsew signal output
rlabel metal2 s 71686 0 71742 800 6 la_data_out[23]
port 286 nsew signal output
rlabel metal2 s 72882 0 72938 800 6 la_data_out[24]
port 287 nsew signal output
rlabel metal2 s 74170 0 74226 800 6 la_data_out[25]
port 288 nsew signal output
rlabel metal2 s 75366 0 75422 800 6 la_data_out[26]
port 289 nsew signal output
rlabel metal2 s 76562 0 76618 800 6 la_data_out[27]
port 290 nsew signal output
rlabel metal2 s 77758 0 77814 800 6 la_data_out[28]
port 291 nsew signal output
rlabel metal2 s 79046 0 79102 800 6 la_data_out[29]
port 292 nsew signal output
rlabel metal2 s 46110 0 46166 800 6 la_data_out[2]
port 293 nsew signal output
rlabel metal2 s 80242 0 80298 800 6 la_data_out[30]
port 294 nsew signal output
rlabel metal2 s 81438 0 81494 800 6 la_data_out[31]
port 295 nsew signal output
rlabel metal2 s 82634 0 82690 800 6 la_data_out[32]
port 296 nsew signal output
rlabel metal2 s 83922 0 83978 800 6 la_data_out[33]
port 297 nsew signal output
rlabel metal2 s 85118 0 85174 800 6 la_data_out[34]
port 298 nsew signal output
rlabel metal2 s 86314 0 86370 800 6 la_data_out[35]
port 299 nsew signal output
rlabel metal2 s 87602 0 87658 800 6 la_data_out[36]
port 300 nsew signal output
rlabel metal2 s 88798 0 88854 800 6 la_data_out[37]
port 301 nsew signal output
rlabel metal2 s 89994 0 90050 800 6 la_data_out[38]
port 302 nsew signal output
rlabel metal2 s 91190 0 91246 800 6 la_data_out[39]
port 303 nsew signal output
rlabel metal2 s 47306 0 47362 800 6 la_data_out[3]
port 304 nsew signal output
rlabel metal2 s 92478 0 92534 800 6 la_data_out[40]
port 305 nsew signal output
rlabel metal2 s 93674 0 93730 800 6 la_data_out[41]
port 306 nsew signal output
rlabel metal2 s 94870 0 94926 800 6 la_data_out[42]
port 307 nsew signal output
rlabel metal2 s 96066 0 96122 800 6 la_data_out[43]
port 308 nsew signal output
rlabel metal2 s 97354 0 97410 800 6 la_data_out[44]
port 309 nsew signal output
rlabel metal2 s 98550 0 98606 800 6 la_data_out[45]
port 310 nsew signal output
rlabel metal2 s 99746 0 99802 800 6 la_data_out[46]
port 311 nsew signal output
rlabel metal2 s 100942 0 100998 800 6 la_data_out[47]
port 312 nsew signal output
rlabel metal2 s 102230 0 102286 800 6 la_data_out[48]
port 313 nsew signal output
rlabel metal2 s 103426 0 103482 800 6 la_data_out[49]
port 314 nsew signal output
rlabel metal2 s 48502 0 48558 800 6 la_data_out[4]
port 315 nsew signal output
rlabel metal2 s 104622 0 104678 800 6 la_data_out[50]
port 316 nsew signal output
rlabel metal2 s 105818 0 105874 800 6 la_data_out[51]
port 317 nsew signal output
rlabel metal2 s 107106 0 107162 800 6 la_data_out[52]
port 318 nsew signal output
rlabel metal2 s 108302 0 108358 800 6 la_data_out[53]
port 319 nsew signal output
rlabel metal2 s 109498 0 109554 800 6 la_data_out[54]
port 320 nsew signal output
rlabel metal2 s 110694 0 110750 800 6 la_data_out[55]
port 321 nsew signal output
rlabel metal2 s 111982 0 112038 800 6 la_data_out[56]
port 322 nsew signal output
rlabel metal2 s 113178 0 113234 800 6 la_data_out[57]
port 323 nsew signal output
rlabel metal2 s 114374 0 114430 800 6 la_data_out[58]
port 324 nsew signal output
rlabel metal2 s 115570 0 115626 800 6 la_data_out[59]
port 325 nsew signal output
rlabel metal2 s 49790 0 49846 800 6 la_data_out[5]
port 326 nsew signal output
rlabel metal2 s 116858 0 116914 800 6 la_data_out[60]
port 327 nsew signal output
rlabel metal2 s 118054 0 118110 800 6 la_data_out[61]
port 328 nsew signal output
rlabel metal2 s 119250 0 119306 800 6 la_data_out[62]
port 329 nsew signal output
rlabel metal2 s 120446 0 120502 800 6 la_data_out[63]
port 330 nsew signal output
rlabel metal2 s 121734 0 121790 800 6 la_data_out[64]
port 331 nsew signal output
rlabel metal2 s 122930 0 122986 800 6 la_data_out[65]
port 332 nsew signal output
rlabel metal2 s 124126 0 124182 800 6 la_data_out[66]
port 333 nsew signal output
rlabel metal2 s 125322 0 125378 800 6 la_data_out[67]
port 334 nsew signal output
rlabel metal2 s 126610 0 126666 800 6 la_data_out[68]
port 335 nsew signal output
rlabel metal2 s 127806 0 127862 800 6 la_data_out[69]
port 336 nsew signal output
rlabel metal2 s 50986 0 51042 800 6 la_data_out[6]
port 337 nsew signal output
rlabel metal2 s 129002 0 129058 800 6 la_data_out[70]
port 338 nsew signal output
rlabel metal2 s 130198 0 130254 800 6 la_data_out[71]
port 339 nsew signal output
rlabel metal2 s 131486 0 131542 800 6 la_data_out[72]
port 340 nsew signal output
rlabel metal2 s 132682 0 132738 800 6 la_data_out[73]
port 341 nsew signal output
rlabel metal2 s 133878 0 133934 800 6 la_data_out[74]
port 342 nsew signal output
rlabel metal2 s 135166 0 135222 800 6 la_data_out[75]
port 343 nsew signal output
rlabel metal2 s 136362 0 136418 800 6 la_data_out[76]
port 344 nsew signal output
rlabel metal2 s 137558 0 137614 800 6 la_data_out[77]
port 345 nsew signal output
rlabel metal2 s 138754 0 138810 800 6 la_data_out[78]
port 346 nsew signal output
rlabel metal2 s 140042 0 140098 800 6 la_data_out[79]
port 347 nsew signal output
rlabel metal2 s 52182 0 52238 800 6 la_data_out[7]
port 348 nsew signal output
rlabel metal2 s 141238 0 141294 800 6 la_data_out[80]
port 349 nsew signal output
rlabel metal2 s 142434 0 142490 800 6 la_data_out[81]
port 350 nsew signal output
rlabel metal2 s 143630 0 143686 800 6 la_data_out[82]
port 351 nsew signal output
rlabel metal2 s 144918 0 144974 800 6 la_data_out[83]
port 352 nsew signal output
rlabel metal2 s 146114 0 146170 800 6 la_data_out[84]
port 353 nsew signal output
rlabel metal2 s 147310 0 147366 800 6 la_data_out[85]
port 354 nsew signal output
rlabel metal2 s 148506 0 148562 800 6 la_data_out[86]
port 355 nsew signal output
rlabel metal2 s 149794 0 149850 800 6 la_data_out[87]
port 356 nsew signal output
rlabel metal2 s 150990 0 151046 800 6 la_data_out[88]
port 357 nsew signal output
rlabel metal2 s 152186 0 152242 800 6 la_data_out[89]
port 358 nsew signal output
rlabel metal2 s 53378 0 53434 800 6 la_data_out[8]
port 359 nsew signal output
rlabel metal2 s 153382 0 153438 800 6 la_data_out[90]
port 360 nsew signal output
rlabel metal2 s 154670 0 154726 800 6 la_data_out[91]
port 361 nsew signal output
rlabel metal2 s 155866 0 155922 800 6 la_data_out[92]
port 362 nsew signal output
rlabel metal2 s 157062 0 157118 800 6 la_data_out[93]
port 363 nsew signal output
rlabel metal2 s 158258 0 158314 800 6 la_data_out[94]
port 364 nsew signal output
rlabel metal2 s 159546 0 159602 800 6 la_data_out[95]
port 365 nsew signal output
rlabel metal2 s 160742 0 160798 800 6 la_data_out[96]
port 366 nsew signal output
rlabel metal2 s 161938 0 161994 800 6 la_data_out[97]
port 367 nsew signal output
rlabel metal2 s 163134 0 163190 800 6 la_data_out[98]
port 368 nsew signal output
rlabel metal2 s 164422 0 164478 800 6 la_data_out[99]
port 369 nsew signal output
rlabel metal2 s 54666 0 54722 800 6 la_data_out[9]
port 370 nsew signal output
rlabel metal2 s 44086 0 44142 800 6 la_oen[0]
port 371 nsew signal input
rlabel metal2 s 165986 0 166042 800 6 la_oen[100]
port 372 nsew signal input
rlabel metal2 s 167274 0 167330 800 6 la_oen[101]
port 373 nsew signal input
rlabel metal2 s 168470 0 168526 800 6 la_oen[102]
port 374 nsew signal input
rlabel metal2 s 169666 0 169722 800 6 la_oen[103]
port 375 nsew signal input
rlabel metal2 s 170862 0 170918 800 6 la_oen[104]
port 376 nsew signal input
rlabel metal2 s 172150 0 172206 800 6 la_oen[105]
port 377 nsew signal input
rlabel metal2 s 173346 0 173402 800 6 la_oen[106]
port 378 nsew signal input
rlabel metal2 s 174542 0 174598 800 6 la_oen[107]
port 379 nsew signal input
rlabel metal2 s 175738 0 175794 800 6 la_oen[108]
port 380 nsew signal input
rlabel metal2 s 177026 0 177082 800 6 la_oen[109]
port 381 nsew signal input
rlabel metal2 s 56230 0 56286 800 6 la_oen[10]
port 382 nsew signal input
rlabel metal2 s 178222 0 178278 800 6 la_oen[110]
port 383 nsew signal input
rlabel metal2 s 179418 0 179474 800 6 la_oen[111]
port 384 nsew signal input
rlabel metal2 s 180614 0 180670 800 6 la_oen[112]
port 385 nsew signal input
rlabel metal2 s 181902 0 181958 800 6 la_oen[113]
port 386 nsew signal input
rlabel metal2 s 183098 0 183154 800 6 la_oen[114]
port 387 nsew signal input
rlabel metal2 s 184294 0 184350 800 6 la_oen[115]
port 388 nsew signal input
rlabel metal2 s 185490 0 185546 800 6 la_oen[116]
port 389 nsew signal input
rlabel metal2 s 186778 0 186834 800 6 la_oen[117]
port 390 nsew signal input
rlabel metal2 s 187974 0 188030 800 6 la_oen[118]
port 391 nsew signal input
rlabel metal2 s 189170 0 189226 800 6 la_oen[119]
port 392 nsew signal input
rlabel metal2 s 57518 0 57574 800 6 la_oen[11]
port 393 nsew signal input
rlabel metal2 s 190366 0 190422 800 6 la_oen[120]
port 394 nsew signal input
rlabel metal2 s 191654 0 191710 800 6 la_oen[121]
port 395 nsew signal input
rlabel metal2 s 192850 0 192906 800 6 la_oen[122]
port 396 nsew signal input
rlabel metal2 s 194046 0 194102 800 6 la_oen[123]
port 397 nsew signal input
rlabel metal2 s 195242 0 195298 800 6 la_oen[124]
port 398 nsew signal input
rlabel metal2 s 196530 0 196586 800 6 la_oen[125]
port 399 nsew signal input
rlabel metal2 s 197726 0 197782 800 6 la_oen[126]
port 400 nsew signal input
rlabel metal2 s 198922 0 198978 800 6 la_oen[127]
port 401 nsew signal input
rlabel metal2 s 58714 0 58770 800 6 la_oen[12]
port 402 nsew signal input
rlabel metal2 s 59910 0 59966 800 6 la_oen[13]
port 403 nsew signal input
rlabel metal2 s 61106 0 61162 800 6 la_oen[14]
port 404 nsew signal input
rlabel metal2 s 62394 0 62450 800 6 la_oen[15]
port 405 nsew signal input
rlabel metal2 s 63590 0 63646 800 6 la_oen[16]
port 406 nsew signal input
rlabel metal2 s 64786 0 64842 800 6 la_oen[17]
port 407 nsew signal input
rlabel metal2 s 65982 0 66038 800 6 la_oen[18]
port 408 nsew signal input
rlabel metal2 s 67270 0 67326 800 6 la_oen[19]
port 409 nsew signal input
rlabel metal2 s 45282 0 45338 800 6 la_oen[1]
port 410 nsew signal input
rlabel metal2 s 68466 0 68522 800 6 la_oen[20]
port 411 nsew signal input
rlabel metal2 s 69662 0 69718 800 6 la_oen[21]
port 412 nsew signal input
rlabel metal2 s 70858 0 70914 800 6 la_oen[22]
port 413 nsew signal input
rlabel metal2 s 72146 0 72202 800 6 la_oen[23]
port 414 nsew signal input
rlabel metal2 s 73342 0 73398 800 6 la_oen[24]
port 415 nsew signal input
rlabel metal2 s 74538 0 74594 800 6 la_oen[25]
port 416 nsew signal input
rlabel metal2 s 75734 0 75790 800 6 la_oen[26]
port 417 nsew signal input
rlabel metal2 s 77022 0 77078 800 6 la_oen[27]
port 418 nsew signal input
rlabel metal2 s 78218 0 78274 800 6 la_oen[28]
port 419 nsew signal input
rlabel metal2 s 79414 0 79470 800 6 la_oen[29]
port 420 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 la_oen[2]
port 421 nsew signal input
rlabel metal2 s 80610 0 80666 800 6 la_oen[30]
port 422 nsew signal input
rlabel metal2 s 81898 0 81954 800 6 la_oen[31]
port 423 nsew signal input
rlabel metal2 s 83094 0 83150 800 6 la_oen[32]
port 424 nsew signal input
rlabel metal2 s 84290 0 84346 800 6 la_oen[33]
port 425 nsew signal input
rlabel metal2 s 85486 0 85542 800 6 la_oen[34]
port 426 nsew signal input
rlabel metal2 s 86774 0 86830 800 6 la_oen[35]
port 427 nsew signal input
rlabel metal2 s 87970 0 88026 800 6 la_oen[36]
port 428 nsew signal input
rlabel metal2 s 89166 0 89222 800 6 la_oen[37]
port 429 nsew signal input
rlabel metal2 s 90362 0 90418 800 6 la_oen[38]
port 430 nsew signal input
rlabel metal2 s 91650 0 91706 800 6 la_oen[39]
port 431 nsew signal input
rlabel metal2 s 47674 0 47730 800 6 la_oen[3]
port 432 nsew signal input
rlabel metal2 s 92846 0 92902 800 6 la_oen[40]
port 433 nsew signal input
rlabel metal2 s 94042 0 94098 800 6 la_oen[41]
port 434 nsew signal input
rlabel metal2 s 95238 0 95294 800 6 la_oen[42]
port 435 nsew signal input
rlabel metal2 s 96526 0 96582 800 6 la_oen[43]
port 436 nsew signal input
rlabel metal2 s 97722 0 97778 800 6 la_oen[44]
port 437 nsew signal input
rlabel metal2 s 98918 0 98974 800 6 la_oen[45]
port 438 nsew signal input
rlabel metal2 s 100206 0 100262 800 6 la_oen[46]
port 439 nsew signal input
rlabel metal2 s 101402 0 101458 800 6 la_oen[47]
port 440 nsew signal input
rlabel metal2 s 102598 0 102654 800 6 la_oen[48]
port 441 nsew signal input
rlabel metal2 s 103794 0 103850 800 6 la_oen[49]
port 442 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 la_oen[4]
port 443 nsew signal input
rlabel metal2 s 105082 0 105138 800 6 la_oen[50]
port 444 nsew signal input
rlabel metal2 s 106278 0 106334 800 6 la_oen[51]
port 445 nsew signal input
rlabel metal2 s 107474 0 107530 800 6 la_oen[52]
port 446 nsew signal input
rlabel metal2 s 108670 0 108726 800 6 la_oen[53]
port 447 nsew signal input
rlabel metal2 s 109958 0 110014 800 6 la_oen[54]
port 448 nsew signal input
rlabel metal2 s 111154 0 111210 800 6 la_oen[55]
port 449 nsew signal input
rlabel metal2 s 112350 0 112406 800 6 la_oen[56]
port 450 nsew signal input
rlabel metal2 s 113546 0 113602 800 6 la_oen[57]
port 451 nsew signal input
rlabel metal2 s 114834 0 114890 800 6 la_oen[58]
port 452 nsew signal input
rlabel metal2 s 116030 0 116086 800 6 la_oen[59]
port 453 nsew signal input
rlabel metal2 s 50158 0 50214 800 6 la_oen[5]
port 454 nsew signal input
rlabel metal2 s 117226 0 117282 800 6 la_oen[60]
port 455 nsew signal input
rlabel metal2 s 118422 0 118478 800 6 la_oen[61]
port 456 nsew signal input
rlabel metal2 s 119710 0 119766 800 6 la_oen[62]
port 457 nsew signal input
rlabel metal2 s 120906 0 120962 800 6 la_oen[63]
port 458 nsew signal input
rlabel metal2 s 122102 0 122158 800 6 la_oen[64]
port 459 nsew signal input
rlabel metal2 s 123298 0 123354 800 6 la_oen[65]
port 460 nsew signal input
rlabel metal2 s 124586 0 124642 800 6 la_oen[66]
port 461 nsew signal input
rlabel metal2 s 125782 0 125838 800 6 la_oen[67]
port 462 nsew signal input
rlabel metal2 s 126978 0 127034 800 6 la_oen[68]
port 463 nsew signal input
rlabel metal2 s 128174 0 128230 800 6 la_oen[69]
port 464 nsew signal input
rlabel metal2 s 51354 0 51410 800 6 la_oen[6]
port 465 nsew signal input
rlabel metal2 s 129462 0 129518 800 6 la_oen[70]
port 466 nsew signal input
rlabel metal2 s 130658 0 130714 800 6 la_oen[71]
port 467 nsew signal input
rlabel metal2 s 131854 0 131910 800 6 la_oen[72]
port 468 nsew signal input
rlabel metal2 s 133050 0 133106 800 6 la_oen[73]
port 469 nsew signal input
rlabel metal2 s 134338 0 134394 800 6 la_oen[74]
port 470 nsew signal input
rlabel metal2 s 135534 0 135590 800 6 la_oen[75]
port 471 nsew signal input
rlabel metal2 s 136730 0 136786 800 6 la_oen[76]
port 472 nsew signal input
rlabel metal2 s 137926 0 137982 800 6 la_oen[77]
port 473 nsew signal input
rlabel metal2 s 139214 0 139270 800 6 la_oen[78]
port 474 nsew signal input
rlabel metal2 s 140410 0 140466 800 6 la_oen[79]
port 475 nsew signal input
rlabel metal2 s 52642 0 52698 800 6 la_oen[7]
port 476 nsew signal input
rlabel metal2 s 141606 0 141662 800 6 la_oen[80]
port 477 nsew signal input
rlabel metal2 s 142802 0 142858 800 6 la_oen[81]
port 478 nsew signal input
rlabel metal2 s 144090 0 144146 800 6 la_oen[82]
port 479 nsew signal input
rlabel metal2 s 145286 0 145342 800 6 la_oen[83]
port 480 nsew signal input
rlabel metal2 s 146482 0 146538 800 6 la_oen[84]
port 481 nsew signal input
rlabel metal2 s 147678 0 147734 800 6 la_oen[85]
port 482 nsew signal input
rlabel metal2 s 148966 0 149022 800 6 la_oen[86]
port 483 nsew signal input
rlabel metal2 s 150162 0 150218 800 6 la_oen[87]
port 484 nsew signal input
rlabel metal2 s 151358 0 151414 800 6 la_oen[88]
port 485 nsew signal input
rlabel metal2 s 152646 0 152702 800 6 la_oen[89]
port 486 nsew signal input
rlabel metal2 s 53838 0 53894 800 6 la_oen[8]
port 487 nsew signal input
rlabel metal2 s 153842 0 153898 800 6 la_oen[90]
port 488 nsew signal input
rlabel metal2 s 155038 0 155094 800 6 la_oen[91]
port 489 nsew signal input
rlabel metal2 s 156234 0 156290 800 6 la_oen[92]
port 490 nsew signal input
rlabel metal2 s 157522 0 157578 800 6 la_oen[93]
port 491 nsew signal input
rlabel metal2 s 158718 0 158774 800 6 la_oen[94]
port 492 nsew signal input
rlabel metal2 s 159914 0 159970 800 6 la_oen[95]
port 493 nsew signal input
rlabel metal2 s 161110 0 161166 800 6 la_oen[96]
port 494 nsew signal input
rlabel metal2 s 162398 0 162454 800 6 la_oen[97]
port 495 nsew signal input
rlabel metal2 s 163594 0 163650 800 6 la_oen[98]
port 496 nsew signal input
rlabel metal2 s 164790 0 164846 800 6 la_oen[99]
port 497 nsew signal input
rlabel metal2 s 55034 0 55090 800 6 la_oen[9]
port 498 nsew signal input
rlabel metal3 s 199200 74944 200000 75064 6 vccd1
port 499 nsew signal bidirectional
rlabel metal2 s 197358 299200 197414 300000 6 vccd2
port 500 nsew signal bidirectional
rlabel metal3 s 0 74944 800 75064 6 vdda1
port 501 nsew signal bidirectional
rlabel metal2 s 199382 0 199438 800 6 vdda2
port 502 nsew signal bidirectional
rlabel metal3 s 0 224952 800 225072 6 vssa1
port 503 nsew signal bidirectional
rlabel metal3 s 199200 224952 200000 225072 6 vssa2
port 504 nsew signal bidirectional
rlabel metal2 s 199750 0 199806 800 6 vssd1
port 505 nsew signal bidirectional
rlabel metal2 s 199106 299200 199162 300000 6 vssd2
port 506 nsew signal bidirectional
rlabel metal2 s 202 0 258 800 6 wb_clk_i
port 507 nsew signal input
rlabel metal2 s 570 0 626 800 6 wb_rst_i
port 508 nsew signal input
rlabel metal2 s 938 0 994 800 6 wbs_ack_o
port 509 nsew signal output
rlabel metal2 s 2594 0 2650 800 6 wbs_adr_i[0]
port 510 nsew signal input
rlabel metal2 s 16394 0 16450 800 6 wbs_adr_i[10]
port 511 nsew signal input
rlabel metal2 s 17682 0 17738 800 6 wbs_adr_i[11]
port 512 nsew signal input
rlabel metal2 s 18878 0 18934 800 6 wbs_adr_i[12]
port 513 nsew signal input
rlabel metal2 s 20074 0 20130 800 6 wbs_adr_i[13]
port 514 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 wbs_adr_i[14]
port 515 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 wbs_adr_i[15]
port 516 nsew signal input
rlabel metal2 s 23754 0 23810 800 6 wbs_adr_i[16]
port 517 nsew signal input
rlabel metal2 s 24950 0 25006 800 6 wbs_adr_i[17]
port 518 nsew signal input
rlabel metal2 s 26146 0 26202 800 6 wbs_adr_i[18]
port 519 nsew signal input
rlabel metal2 s 27434 0 27490 800 6 wbs_adr_i[19]
port 520 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 wbs_adr_i[1]
port 521 nsew signal input
rlabel metal2 s 28630 0 28686 800 6 wbs_adr_i[20]
port 522 nsew signal input
rlabel metal2 s 29826 0 29882 800 6 wbs_adr_i[21]
port 523 nsew signal input
rlabel metal2 s 31022 0 31078 800 6 wbs_adr_i[22]
port 524 nsew signal input
rlabel metal2 s 32310 0 32366 800 6 wbs_adr_i[23]
port 525 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 wbs_adr_i[24]
port 526 nsew signal input
rlabel metal2 s 34702 0 34758 800 6 wbs_adr_i[25]
port 527 nsew signal input
rlabel metal2 s 35898 0 35954 800 6 wbs_adr_i[26]
port 528 nsew signal input
rlabel metal2 s 37186 0 37242 800 6 wbs_adr_i[27]
port 529 nsew signal input
rlabel metal2 s 38382 0 38438 800 6 wbs_adr_i[28]
port 530 nsew signal input
rlabel metal2 s 39578 0 39634 800 6 wbs_adr_i[29]
port 531 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 wbs_adr_i[2]
port 532 nsew signal input
rlabel metal2 s 40774 0 40830 800 6 wbs_adr_i[30]
port 533 nsew signal input
rlabel metal2 s 42062 0 42118 800 6 wbs_adr_i[31]
port 534 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 wbs_adr_i[3]
port 535 nsew signal input
rlabel metal2 s 9126 0 9182 800 6 wbs_adr_i[4]
port 536 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 wbs_adr_i[5]
port 537 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 wbs_adr_i[6]
port 538 nsew signal input
rlabel metal2 s 12714 0 12770 800 6 wbs_adr_i[7]
port 539 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 wbs_adr_i[8]
port 540 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 wbs_adr_i[9]
port 541 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 wbs_cyc_i
port 542 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 wbs_dat_i[0]
port 543 nsew signal input
rlabel metal2 s 16854 0 16910 800 6 wbs_dat_i[10]
port 544 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 wbs_dat_i[11]
port 545 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 wbs_dat_i[12]
port 546 nsew signal input
rlabel metal2 s 20442 0 20498 800 6 wbs_dat_i[13]
port 547 nsew signal input
rlabel metal2 s 21730 0 21786 800 6 wbs_dat_i[14]
port 548 nsew signal input
rlabel metal2 s 22926 0 22982 800 6 wbs_dat_i[15]
port 549 nsew signal input
rlabel metal2 s 24122 0 24178 800 6 wbs_dat_i[16]
port 550 nsew signal input
rlabel metal2 s 25318 0 25374 800 6 wbs_dat_i[17]
port 551 nsew signal input
rlabel metal2 s 26606 0 26662 800 6 wbs_dat_i[18]
port 552 nsew signal input
rlabel metal2 s 27802 0 27858 800 6 wbs_dat_i[19]
port 553 nsew signal input
rlabel metal2 s 4618 0 4674 800 6 wbs_dat_i[1]
port 554 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 wbs_dat_i[20]
port 555 nsew signal input
rlabel metal2 s 30194 0 30250 800 6 wbs_dat_i[21]
port 556 nsew signal input
rlabel metal2 s 31482 0 31538 800 6 wbs_dat_i[22]
port 557 nsew signal input
rlabel metal2 s 32678 0 32734 800 6 wbs_dat_i[23]
port 558 nsew signal input
rlabel metal2 s 33874 0 33930 800 6 wbs_dat_i[24]
port 559 nsew signal input
rlabel metal2 s 35162 0 35218 800 6 wbs_dat_i[25]
port 560 nsew signal input
rlabel metal2 s 36358 0 36414 800 6 wbs_dat_i[26]
port 561 nsew signal input
rlabel metal2 s 37554 0 37610 800 6 wbs_dat_i[27]
port 562 nsew signal input
rlabel metal2 s 38750 0 38806 800 6 wbs_dat_i[28]
port 563 nsew signal input
rlabel metal2 s 40038 0 40094 800 6 wbs_dat_i[29]
port 564 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 wbs_dat_i[2]
port 565 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 wbs_dat_i[30]
port 566 nsew signal input
rlabel metal2 s 42430 0 42486 800 6 wbs_dat_i[31]
port 567 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 wbs_dat_i[3]
port 568 nsew signal input
rlabel metal2 s 9494 0 9550 800 6 wbs_dat_i[4]
port 569 nsew signal input
rlabel metal2 s 10690 0 10746 800 6 wbs_dat_i[5]
port 570 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 wbs_dat_i[6]
port 571 nsew signal input
rlabel metal2 s 13174 0 13230 800 6 wbs_dat_i[7]
port 572 nsew signal input
rlabel metal2 s 14370 0 14426 800 6 wbs_dat_i[8]
port 573 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 wbs_dat_i[9]
port 574 nsew signal input
rlabel metal2 s 3422 0 3478 800 6 wbs_dat_o[0]
port 575 nsew signal output
rlabel metal2 s 17222 0 17278 800 6 wbs_dat_o[10]
port 576 nsew signal output
rlabel metal2 s 18418 0 18474 800 6 wbs_dat_o[11]
port 577 nsew signal output
rlabel metal2 s 19706 0 19762 800 6 wbs_dat_o[12]
port 578 nsew signal output
rlabel metal2 s 20902 0 20958 800 6 wbs_dat_o[13]
port 579 nsew signal output
rlabel metal2 s 22098 0 22154 800 6 wbs_dat_o[14]
port 580 nsew signal output
rlabel metal2 s 23294 0 23350 800 6 wbs_dat_o[15]
port 581 nsew signal output
rlabel metal2 s 24582 0 24638 800 6 wbs_dat_o[16]
port 582 nsew signal output
rlabel metal2 s 25778 0 25834 800 6 wbs_dat_o[17]
port 583 nsew signal output
rlabel metal2 s 26974 0 27030 800 6 wbs_dat_o[18]
port 584 nsew signal output
rlabel metal2 s 28170 0 28226 800 6 wbs_dat_o[19]
port 585 nsew signal output
rlabel metal2 s 5078 0 5134 800 6 wbs_dat_o[1]
port 586 nsew signal output
rlabel metal2 s 29458 0 29514 800 6 wbs_dat_o[20]
port 587 nsew signal output
rlabel metal2 s 30654 0 30710 800 6 wbs_dat_o[21]
port 588 nsew signal output
rlabel metal2 s 31850 0 31906 800 6 wbs_dat_o[22]
port 589 nsew signal output
rlabel metal2 s 33046 0 33102 800 6 wbs_dat_o[23]
port 590 nsew signal output
rlabel metal2 s 34334 0 34390 800 6 wbs_dat_o[24]
port 591 nsew signal output
rlabel metal2 s 35530 0 35586 800 6 wbs_dat_o[25]
port 592 nsew signal output
rlabel metal2 s 36726 0 36782 800 6 wbs_dat_o[26]
port 593 nsew signal output
rlabel metal2 s 37922 0 37978 800 6 wbs_dat_o[27]
port 594 nsew signal output
rlabel metal2 s 39210 0 39266 800 6 wbs_dat_o[28]
port 595 nsew signal output
rlabel metal2 s 40406 0 40462 800 6 wbs_dat_o[29]
port 596 nsew signal output
rlabel metal2 s 6642 0 6698 800 6 wbs_dat_o[2]
port 597 nsew signal output
rlabel metal2 s 41602 0 41658 800 6 wbs_dat_o[30]
port 598 nsew signal output
rlabel metal2 s 42798 0 42854 800 6 wbs_dat_o[31]
port 599 nsew signal output
rlabel metal2 s 8298 0 8354 800 6 wbs_dat_o[3]
port 600 nsew signal output
rlabel metal2 s 9954 0 10010 800 6 wbs_dat_o[4]
port 601 nsew signal output
rlabel metal2 s 11150 0 11206 800 6 wbs_dat_o[5]
port 602 nsew signal output
rlabel metal2 s 12346 0 12402 800 6 wbs_dat_o[6]
port 603 nsew signal output
rlabel metal2 s 13542 0 13598 800 6 wbs_dat_o[7]
port 604 nsew signal output
rlabel metal2 s 14830 0 14886 800 6 wbs_dat_o[8]
port 605 nsew signal output
rlabel metal2 s 16026 0 16082 800 6 wbs_dat_o[9]
port 606 nsew signal output
rlabel metal2 s 3790 0 3846 800 6 wbs_sel_i[0]
port 607 nsew signal input
rlabel metal2 s 5446 0 5502 800 6 wbs_sel_i[1]
port 608 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 wbs_sel_i[2]
port 609 nsew signal input
rlabel metal2 s 8666 0 8722 800 6 wbs_sel_i[3]
port 610 nsew signal input
rlabel metal2 s 1766 0 1822 800 6 wbs_stb_i
port 611 nsew signal input
rlabel metal2 s 2226 0 2282 800 6 wbs_we_i
port 612 nsew signal input
rlabel metal4 s 188528 2128 188848 297616 6 VPWR
port 613 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 297616 6 VPWR
port 614 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 297616 6 VPWR
port 615 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 297616 6 VPWR
port 616 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 297616 6 VPWR
port 617 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 297616 6 VPWR
port 618 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 297616 6 VPWR
port 619 nsew power bidirectional
rlabel metal4 s 173168 2128 173488 297616 6 VGND
port 620 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 297616 6 VGND
port 621 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 297616 6 VGND
port 622 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 297616 6 VGND
port 623 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 297616 6 VGND
port 624 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 297616 6 VGND
port 625 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 200000 300000
string LEFview TRUE
<< end >>
