magic
tech sky130A
magscale 1 2
timestamp 1611867494
<< obsli1 >>
rect 1104 2159 398820 497777
<< obsm1 >>
rect 382 1232 398820 497808
<< metal2 >>
rect 1674 499200 1730 500000
rect 5078 499200 5134 500000
rect 8482 499200 8538 500000
rect 11886 499200 11942 500000
rect 15290 499200 15346 500000
rect 18694 499200 18750 500000
rect 22098 499200 22154 500000
rect 25594 499200 25650 500000
rect 28998 499200 29054 500000
rect 32402 499200 32458 500000
rect 35806 499200 35862 500000
rect 39210 499200 39266 500000
rect 42614 499200 42670 500000
rect 46110 499200 46166 500000
rect 49514 499200 49570 500000
rect 52918 499200 52974 500000
rect 56322 499200 56378 500000
rect 59726 499200 59782 500000
rect 63130 499200 63186 500000
rect 66626 499200 66682 500000
rect 70030 499200 70086 500000
rect 73434 499200 73490 500000
rect 76838 499200 76894 500000
rect 80242 499200 80298 500000
rect 83646 499200 83702 500000
rect 87142 499200 87198 500000
rect 90546 499200 90602 500000
rect 93950 499200 94006 500000
rect 97354 499200 97410 500000
rect 100758 499200 100814 500000
rect 104162 499200 104218 500000
rect 107658 499200 107714 500000
rect 111062 499200 111118 500000
rect 114466 499200 114522 500000
rect 117870 499200 117926 500000
rect 121274 499200 121330 500000
rect 124678 499200 124734 500000
rect 128174 499200 128230 500000
rect 131578 499200 131634 500000
rect 134982 499200 135038 500000
rect 138386 499200 138442 500000
rect 141790 499200 141846 500000
rect 145194 499200 145250 500000
rect 148598 499200 148654 500000
rect 152094 499200 152150 500000
rect 155498 499200 155554 500000
rect 158902 499200 158958 500000
rect 162306 499200 162362 500000
rect 165710 499200 165766 500000
rect 169114 499200 169170 500000
rect 172610 499200 172666 500000
rect 176014 499200 176070 500000
rect 179418 499200 179474 500000
rect 182822 499200 182878 500000
rect 186226 499200 186282 500000
rect 189630 499200 189686 500000
rect 193126 499200 193182 500000
rect 196530 499200 196586 500000
rect 199934 499200 199990 500000
rect 203338 499200 203394 500000
rect 206742 499200 206798 500000
rect 210146 499200 210202 500000
rect 213642 499200 213698 500000
rect 217046 499200 217102 500000
rect 220450 499200 220506 500000
rect 223854 499200 223910 500000
rect 227258 499200 227314 500000
rect 230662 499200 230718 500000
rect 234158 499200 234214 500000
rect 237562 499200 237618 500000
rect 240966 499200 241022 500000
rect 244370 499200 244426 500000
rect 247774 499200 247830 500000
rect 251178 499200 251234 500000
rect 254674 499200 254730 500000
rect 258078 499200 258134 500000
rect 261482 499200 261538 500000
rect 264886 499200 264942 500000
rect 268290 499200 268346 500000
rect 271694 499200 271750 500000
rect 275098 499200 275154 500000
rect 278594 499200 278650 500000
rect 281998 499200 282054 500000
rect 285402 499200 285458 500000
rect 288806 499200 288862 500000
rect 292210 499200 292266 500000
rect 295614 499200 295670 500000
rect 299110 499200 299166 500000
rect 302514 499200 302570 500000
rect 305918 499200 305974 500000
rect 309322 499200 309378 500000
rect 312726 499200 312782 500000
rect 316130 499200 316186 500000
rect 319626 499200 319682 500000
rect 323030 499200 323086 500000
rect 326434 499200 326490 500000
rect 329838 499200 329894 500000
rect 333242 499200 333298 500000
rect 336646 499200 336702 500000
rect 340142 499200 340198 500000
rect 343546 499200 343602 500000
rect 346950 499200 347006 500000
rect 350354 499200 350410 500000
rect 353758 499200 353814 500000
rect 357162 499200 357218 500000
rect 360658 499200 360714 500000
rect 364062 499200 364118 500000
rect 367466 499200 367522 500000
rect 370870 499200 370926 500000
rect 374274 499200 374330 500000
rect 377678 499200 377734 500000
rect 381174 499200 381230 500000
rect 384578 499200 384634 500000
rect 387982 499200 388038 500000
rect 391386 499200 391442 500000
rect 394790 499200 394846 500000
rect 398194 499200 398250 500000
rect 386 0 442 800
rect 1122 0 1178 800
rect 1950 0 2006 800
rect 2778 0 2834 800
rect 3606 0 3662 800
rect 4434 0 4490 800
rect 5262 0 5318 800
rect 5998 0 6054 800
rect 6826 0 6882 800
rect 7654 0 7710 800
rect 8482 0 8538 800
rect 9310 0 9366 800
rect 10138 0 10194 800
rect 10874 0 10930 800
rect 11702 0 11758 800
rect 12530 0 12586 800
rect 13358 0 13414 800
rect 14186 0 14242 800
rect 15014 0 15070 800
rect 15750 0 15806 800
rect 16578 0 16634 800
rect 17406 0 17462 800
rect 18234 0 18290 800
rect 19062 0 19118 800
rect 19890 0 19946 800
rect 20626 0 20682 800
rect 21454 0 21510 800
rect 22282 0 22338 800
rect 23110 0 23166 800
rect 23938 0 23994 800
rect 24766 0 24822 800
rect 25502 0 25558 800
rect 26330 0 26386 800
rect 27158 0 27214 800
rect 27986 0 28042 800
rect 28814 0 28870 800
rect 29642 0 29698 800
rect 30378 0 30434 800
rect 31206 0 31262 800
rect 32034 0 32090 800
rect 32862 0 32918 800
rect 33690 0 33746 800
rect 34518 0 34574 800
rect 35346 0 35402 800
rect 36082 0 36138 800
rect 36910 0 36966 800
rect 37738 0 37794 800
rect 38566 0 38622 800
rect 39394 0 39450 800
rect 40222 0 40278 800
rect 40958 0 41014 800
rect 41786 0 41842 800
rect 42614 0 42670 800
rect 43442 0 43498 800
rect 44270 0 44326 800
rect 45098 0 45154 800
rect 45834 0 45890 800
rect 46662 0 46718 800
rect 47490 0 47546 800
rect 48318 0 48374 800
rect 49146 0 49202 800
rect 49974 0 50030 800
rect 50710 0 50766 800
rect 51538 0 51594 800
rect 52366 0 52422 800
rect 53194 0 53250 800
rect 54022 0 54078 800
rect 54850 0 54906 800
rect 55586 0 55642 800
rect 56414 0 56470 800
rect 57242 0 57298 800
rect 58070 0 58126 800
rect 58898 0 58954 800
rect 59726 0 59782 800
rect 60462 0 60518 800
rect 61290 0 61346 800
rect 62118 0 62174 800
rect 62946 0 63002 800
rect 63774 0 63830 800
rect 64602 0 64658 800
rect 65338 0 65394 800
rect 66166 0 66222 800
rect 66994 0 67050 800
rect 67822 0 67878 800
rect 68650 0 68706 800
rect 69478 0 69534 800
rect 70306 0 70362 800
rect 71042 0 71098 800
rect 71870 0 71926 800
rect 72698 0 72754 800
rect 73526 0 73582 800
rect 74354 0 74410 800
rect 75182 0 75238 800
rect 75918 0 75974 800
rect 76746 0 76802 800
rect 77574 0 77630 800
rect 78402 0 78458 800
rect 79230 0 79286 800
rect 80058 0 80114 800
rect 80794 0 80850 800
rect 81622 0 81678 800
rect 82450 0 82506 800
rect 83278 0 83334 800
rect 84106 0 84162 800
rect 84934 0 84990 800
rect 85670 0 85726 800
rect 86498 0 86554 800
rect 87326 0 87382 800
rect 88154 0 88210 800
rect 88982 0 89038 800
rect 89810 0 89866 800
rect 90546 0 90602 800
rect 91374 0 91430 800
rect 92202 0 92258 800
rect 93030 0 93086 800
rect 93858 0 93914 800
rect 94686 0 94742 800
rect 95422 0 95478 800
rect 96250 0 96306 800
rect 97078 0 97134 800
rect 97906 0 97962 800
rect 98734 0 98790 800
rect 99562 0 99618 800
rect 100390 0 100446 800
rect 101126 0 101182 800
rect 101954 0 102010 800
rect 102782 0 102838 800
rect 103610 0 103666 800
rect 104438 0 104494 800
rect 105266 0 105322 800
rect 106002 0 106058 800
rect 106830 0 106886 800
rect 107658 0 107714 800
rect 108486 0 108542 800
rect 109314 0 109370 800
rect 110142 0 110198 800
rect 110878 0 110934 800
rect 111706 0 111762 800
rect 112534 0 112590 800
rect 113362 0 113418 800
rect 114190 0 114246 800
rect 115018 0 115074 800
rect 115754 0 115810 800
rect 116582 0 116638 800
rect 117410 0 117466 800
rect 118238 0 118294 800
rect 119066 0 119122 800
rect 119894 0 119950 800
rect 120630 0 120686 800
rect 121458 0 121514 800
rect 122286 0 122342 800
rect 123114 0 123170 800
rect 123942 0 123998 800
rect 124770 0 124826 800
rect 125506 0 125562 800
rect 126334 0 126390 800
rect 127162 0 127218 800
rect 127990 0 128046 800
rect 128818 0 128874 800
rect 129646 0 129702 800
rect 130382 0 130438 800
rect 131210 0 131266 800
rect 132038 0 132094 800
rect 132866 0 132922 800
rect 133694 0 133750 800
rect 134522 0 134578 800
rect 135350 0 135406 800
rect 136086 0 136142 800
rect 136914 0 136970 800
rect 137742 0 137798 800
rect 138570 0 138626 800
rect 139398 0 139454 800
rect 140226 0 140282 800
rect 140962 0 141018 800
rect 141790 0 141846 800
rect 142618 0 142674 800
rect 143446 0 143502 800
rect 144274 0 144330 800
rect 145102 0 145158 800
rect 145838 0 145894 800
rect 146666 0 146722 800
rect 147494 0 147550 800
rect 148322 0 148378 800
rect 149150 0 149206 800
rect 149978 0 150034 800
rect 150714 0 150770 800
rect 151542 0 151598 800
rect 152370 0 152426 800
rect 153198 0 153254 800
rect 154026 0 154082 800
rect 154854 0 154910 800
rect 155590 0 155646 800
rect 156418 0 156474 800
rect 157246 0 157302 800
rect 158074 0 158130 800
rect 158902 0 158958 800
rect 159730 0 159786 800
rect 160466 0 160522 800
rect 161294 0 161350 800
rect 162122 0 162178 800
rect 162950 0 163006 800
rect 163778 0 163834 800
rect 164606 0 164662 800
rect 165342 0 165398 800
rect 166170 0 166226 800
rect 166998 0 167054 800
rect 167826 0 167882 800
rect 168654 0 168710 800
rect 169482 0 169538 800
rect 170310 0 170366 800
rect 171046 0 171102 800
rect 171874 0 171930 800
rect 172702 0 172758 800
rect 173530 0 173586 800
rect 174358 0 174414 800
rect 175186 0 175242 800
rect 175922 0 175978 800
rect 176750 0 176806 800
rect 177578 0 177634 800
rect 178406 0 178462 800
rect 179234 0 179290 800
rect 180062 0 180118 800
rect 180798 0 180854 800
rect 181626 0 181682 800
rect 182454 0 182510 800
rect 183282 0 183338 800
rect 184110 0 184166 800
rect 184938 0 184994 800
rect 185674 0 185730 800
rect 186502 0 186558 800
rect 187330 0 187386 800
rect 188158 0 188214 800
rect 188986 0 189042 800
rect 189814 0 189870 800
rect 190550 0 190606 800
rect 191378 0 191434 800
rect 192206 0 192262 800
rect 193034 0 193090 800
rect 193862 0 193918 800
rect 194690 0 194746 800
rect 195426 0 195482 800
rect 196254 0 196310 800
rect 197082 0 197138 800
rect 197910 0 197966 800
rect 198738 0 198794 800
rect 199566 0 199622 800
rect 200394 0 200450 800
rect 201130 0 201186 800
rect 201958 0 202014 800
rect 202786 0 202842 800
rect 203614 0 203670 800
rect 204442 0 204498 800
rect 205270 0 205326 800
rect 206006 0 206062 800
rect 206834 0 206890 800
rect 207662 0 207718 800
rect 208490 0 208546 800
rect 209318 0 209374 800
rect 210146 0 210202 800
rect 210882 0 210938 800
rect 211710 0 211766 800
rect 212538 0 212594 800
rect 213366 0 213422 800
rect 214194 0 214250 800
rect 215022 0 215078 800
rect 215758 0 215814 800
rect 216586 0 216642 800
rect 217414 0 217470 800
rect 218242 0 218298 800
rect 219070 0 219126 800
rect 219898 0 219954 800
rect 220634 0 220690 800
rect 221462 0 221518 800
rect 222290 0 222346 800
rect 223118 0 223174 800
rect 223946 0 224002 800
rect 224774 0 224830 800
rect 225510 0 225566 800
rect 226338 0 226394 800
rect 227166 0 227222 800
rect 227994 0 228050 800
rect 228822 0 228878 800
rect 229650 0 229706 800
rect 230386 0 230442 800
rect 231214 0 231270 800
rect 232042 0 232098 800
rect 232870 0 232926 800
rect 233698 0 233754 800
rect 234526 0 234582 800
rect 235354 0 235410 800
rect 236090 0 236146 800
rect 236918 0 236974 800
rect 237746 0 237802 800
rect 238574 0 238630 800
rect 239402 0 239458 800
rect 240230 0 240286 800
rect 240966 0 241022 800
rect 241794 0 241850 800
rect 242622 0 242678 800
rect 243450 0 243506 800
rect 244278 0 244334 800
rect 245106 0 245162 800
rect 245842 0 245898 800
rect 246670 0 246726 800
rect 247498 0 247554 800
rect 248326 0 248382 800
rect 249154 0 249210 800
rect 249982 0 250038 800
rect 250718 0 250774 800
rect 251546 0 251602 800
rect 252374 0 252430 800
rect 253202 0 253258 800
rect 254030 0 254086 800
rect 254858 0 254914 800
rect 255594 0 255650 800
rect 256422 0 256478 800
rect 257250 0 257306 800
rect 258078 0 258134 800
rect 258906 0 258962 800
rect 259734 0 259790 800
rect 260470 0 260526 800
rect 261298 0 261354 800
rect 262126 0 262182 800
rect 262954 0 263010 800
rect 263782 0 263838 800
rect 264610 0 264666 800
rect 265346 0 265402 800
rect 266174 0 266230 800
rect 267002 0 267058 800
rect 267830 0 267886 800
rect 268658 0 268714 800
rect 269486 0 269542 800
rect 270314 0 270370 800
rect 271050 0 271106 800
rect 271878 0 271934 800
rect 272706 0 272762 800
rect 273534 0 273590 800
rect 274362 0 274418 800
rect 275190 0 275246 800
rect 275926 0 275982 800
rect 276754 0 276810 800
rect 277582 0 277638 800
rect 278410 0 278466 800
rect 279238 0 279294 800
rect 280066 0 280122 800
rect 280802 0 280858 800
rect 281630 0 281686 800
rect 282458 0 282514 800
rect 283286 0 283342 800
rect 284114 0 284170 800
rect 284942 0 284998 800
rect 285678 0 285734 800
rect 286506 0 286562 800
rect 287334 0 287390 800
rect 288162 0 288218 800
rect 288990 0 289046 800
rect 289818 0 289874 800
rect 290554 0 290610 800
rect 291382 0 291438 800
rect 292210 0 292266 800
rect 293038 0 293094 800
rect 293866 0 293922 800
rect 294694 0 294750 800
rect 295430 0 295486 800
rect 296258 0 296314 800
rect 297086 0 297142 800
rect 297914 0 297970 800
rect 298742 0 298798 800
rect 299570 0 299626 800
rect 300398 0 300454 800
rect 301134 0 301190 800
rect 301962 0 302018 800
rect 302790 0 302846 800
rect 303618 0 303674 800
rect 304446 0 304502 800
rect 305274 0 305330 800
rect 306010 0 306066 800
rect 306838 0 306894 800
rect 307666 0 307722 800
rect 308494 0 308550 800
rect 309322 0 309378 800
rect 310150 0 310206 800
rect 310886 0 310942 800
rect 311714 0 311770 800
rect 312542 0 312598 800
rect 313370 0 313426 800
rect 314198 0 314254 800
rect 315026 0 315082 800
rect 315762 0 315818 800
rect 316590 0 316646 800
rect 317418 0 317474 800
rect 318246 0 318302 800
rect 319074 0 319130 800
rect 319902 0 319958 800
rect 320638 0 320694 800
rect 321466 0 321522 800
rect 322294 0 322350 800
rect 323122 0 323178 800
rect 323950 0 324006 800
rect 324778 0 324834 800
rect 325514 0 325570 800
rect 326342 0 326398 800
rect 327170 0 327226 800
rect 327998 0 328054 800
rect 328826 0 328882 800
rect 329654 0 329710 800
rect 330390 0 330446 800
rect 331218 0 331274 800
rect 332046 0 332102 800
rect 332874 0 332930 800
rect 333702 0 333758 800
rect 334530 0 334586 800
rect 335358 0 335414 800
rect 336094 0 336150 800
rect 336922 0 336978 800
rect 337750 0 337806 800
rect 338578 0 338634 800
rect 339406 0 339462 800
rect 340234 0 340290 800
rect 340970 0 341026 800
rect 341798 0 341854 800
rect 342626 0 342682 800
rect 343454 0 343510 800
rect 344282 0 344338 800
rect 345110 0 345166 800
rect 345846 0 345902 800
rect 346674 0 346730 800
rect 347502 0 347558 800
rect 348330 0 348386 800
rect 349158 0 349214 800
rect 349986 0 350042 800
rect 350722 0 350778 800
rect 351550 0 351606 800
rect 352378 0 352434 800
rect 353206 0 353262 800
rect 354034 0 354090 800
rect 354862 0 354918 800
rect 355598 0 355654 800
rect 356426 0 356482 800
rect 357254 0 357310 800
rect 358082 0 358138 800
rect 358910 0 358966 800
rect 359738 0 359794 800
rect 360474 0 360530 800
rect 361302 0 361358 800
rect 362130 0 362186 800
rect 362958 0 363014 800
rect 363786 0 363842 800
rect 364614 0 364670 800
rect 365350 0 365406 800
rect 366178 0 366234 800
rect 367006 0 367062 800
rect 367834 0 367890 800
rect 368662 0 368718 800
rect 369490 0 369546 800
rect 370318 0 370374 800
rect 371054 0 371110 800
rect 371882 0 371938 800
rect 372710 0 372766 800
rect 373538 0 373594 800
rect 374366 0 374422 800
rect 375194 0 375250 800
rect 375930 0 375986 800
rect 376758 0 376814 800
rect 377586 0 377642 800
rect 378414 0 378470 800
rect 379242 0 379298 800
rect 380070 0 380126 800
rect 380806 0 380862 800
rect 381634 0 381690 800
rect 382462 0 382518 800
rect 383290 0 383346 800
rect 384118 0 384174 800
rect 384946 0 385002 800
rect 385682 0 385738 800
rect 386510 0 386566 800
rect 387338 0 387394 800
rect 388166 0 388222 800
rect 388994 0 389050 800
rect 389822 0 389878 800
rect 390558 0 390614 800
rect 391386 0 391442 800
rect 392214 0 392270 800
rect 393042 0 393098 800
rect 393870 0 393926 800
rect 394698 0 394754 800
rect 395434 0 395490 800
rect 396262 0 396318 800
rect 397090 0 397146 800
rect 397918 0 397974 800
rect 398746 0 398802 800
rect 399574 0 399630 800
<< obsm2 >>
rect 388 499144 1618 499200
rect 1786 499144 5022 499200
rect 5190 499144 8426 499200
rect 8594 499144 11830 499200
rect 11998 499144 15234 499200
rect 15402 499144 18638 499200
rect 18806 499144 22042 499200
rect 22210 499144 25538 499200
rect 25706 499144 28942 499200
rect 29110 499144 32346 499200
rect 32514 499144 35750 499200
rect 35918 499144 39154 499200
rect 39322 499144 42558 499200
rect 42726 499144 46054 499200
rect 46222 499144 49458 499200
rect 49626 499144 52862 499200
rect 53030 499144 56266 499200
rect 56434 499144 59670 499200
rect 59838 499144 63074 499200
rect 63242 499144 66570 499200
rect 66738 499144 69974 499200
rect 70142 499144 73378 499200
rect 73546 499144 76782 499200
rect 76950 499144 80186 499200
rect 80354 499144 83590 499200
rect 83758 499144 87086 499200
rect 87254 499144 90490 499200
rect 90658 499144 93894 499200
rect 94062 499144 97298 499200
rect 97466 499144 100702 499200
rect 100870 499144 104106 499200
rect 104274 499144 107602 499200
rect 107770 499144 111006 499200
rect 111174 499144 114410 499200
rect 114578 499144 117814 499200
rect 117982 499144 121218 499200
rect 121386 499144 124622 499200
rect 124790 499144 128118 499200
rect 128286 499144 131522 499200
rect 131690 499144 134926 499200
rect 135094 499144 138330 499200
rect 138498 499144 141734 499200
rect 141902 499144 145138 499200
rect 145306 499144 148542 499200
rect 148710 499144 152038 499200
rect 152206 499144 155442 499200
rect 155610 499144 158846 499200
rect 159014 499144 162250 499200
rect 162418 499144 165654 499200
rect 165822 499144 169058 499200
rect 169226 499144 172554 499200
rect 172722 499144 175958 499200
rect 176126 499144 179362 499200
rect 179530 499144 182766 499200
rect 182934 499144 186170 499200
rect 186338 499144 189574 499200
rect 189742 499144 193070 499200
rect 193238 499144 196474 499200
rect 196642 499144 199878 499200
rect 200046 499144 203282 499200
rect 203450 499144 206686 499200
rect 206854 499144 210090 499200
rect 210258 499144 213586 499200
rect 213754 499144 216990 499200
rect 217158 499144 220394 499200
rect 220562 499144 223798 499200
rect 223966 499144 227202 499200
rect 227370 499144 230606 499200
rect 230774 499144 234102 499200
rect 234270 499144 237506 499200
rect 237674 499144 240910 499200
rect 241078 499144 244314 499200
rect 244482 499144 247718 499200
rect 247886 499144 251122 499200
rect 251290 499144 254618 499200
rect 254786 499144 258022 499200
rect 258190 499144 261426 499200
rect 261594 499144 264830 499200
rect 264998 499144 268234 499200
rect 268402 499144 271638 499200
rect 271806 499144 275042 499200
rect 275210 499144 278538 499200
rect 278706 499144 281942 499200
rect 282110 499144 285346 499200
rect 285514 499144 288750 499200
rect 288918 499144 292154 499200
rect 292322 499144 295558 499200
rect 295726 499144 299054 499200
rect 299222 499144 302458 499200
rect 302626 499144 305862 499200
rect 306030 499144 309266 499200
rect 309434 499144 312670 499200
rect 312838 499144 316074 499200
rect 316242 499144 319570 499200
rect 319738 499144 322974 499200
rect 323142 499144 326378 499200
rect 326546 499144 329782 499200
rect 329950 499144 333186 499200
rect 333354 499144 336590 499200
rect 336758 499144 340086 499200
rect 340254 499144 343490 499200
rect 343658 499144 346894 499200
rect 347062 499144 350298 499200
rect 350466 499144 353702 499200
rect 353870 499144 357106 499200
rect 357274 499144 360602 499200
rect 360770 499144 364006 499200
rect 364174 499144 367410 499200
rect 367578 499144 370814 499200
rect 370982 499144 374218 499200
rect 374386 499144 377622 499200
rect 377790 499144 381118 499200
rect 381286 499144 384522 499200
rect 384690 499144 387926 499200
rect 388094 499144 391330 499200
rect 391498 499144 394734 499200
rect 394902 499144 397144 499200
rect 388 856 397144 499144
rect 498 800 1066 856
rect 1234 800 1894 856
rect 2062 800 2722 856
rect 2890 800 3550 856
rect 3718 800 4378 856
rect 4546 800 5206 856
rect 5374 800 5942 856
rect 6110 800 6770 856
rect 6938 800 7598 856
rect 7766 800 8426 856
rect 8594 800 9254 856
rect 9422 800 10082 856
rect 10250 800 10818 856
rect 10986 800 11646 856
rect 11814 800 12474 856
rect 12642 800 13302 856
rect 13470 800 14130 856
rect 14298 800 14958 856
rect 15126 800 15694 856
rect 15862 800 16522 856
rect 16690 800 17350 856
rect 17518 800 18178 856
rect 18346 800 19006 856
rect 19174 800 19834 856
rect 20002 800 20570 856
rect 20738 800 21398 856
rect 21566 800 22226 856
rect 22394 800 23054 856
rect 23222 800 23882 856
rect 24050 800 24710 856
rect 24878 800 25446 856
rect 25614 800 26274 856
rect 26442 800 27102 856
rect 27270 800 27930 856
rect 28098 800 28758 856
rect 28926 800 29586 856
rect 29754 800 30322 856
rect 30490 800 31150 856
rect 31318 800 31978 856
rect 32146 800 32806 856
rect 32974 800 33634 856
rect 33802 800 34462 856
rect 34630 800 35290 856
rect 35458 800 36026 856
rect 36194 800 36854 856
rect 37022 800 37682 856
rect 37850 800 38510 856
rect 38678 800 39338 856
rect 39506 800 40166 856
rect 40334 800 40902 856
rect 41070 800 41730 856
rect 41898 800 42558 856
rect 42726 800 43386 856
rect 43554 800 44214 856
rect 44382 800 45042 856
rect 45210 800 45778 856
rect 45946 800 46606 856
rect 46774 800 47434 856
rect 47602 800 48262 856
rect 48430 800 49090 856
rect 49258 800 49918 856
rect 50086 800 50654 856
rect 50822 800 51482 856
rect 51650 800 52310 856
rect 52478 800 53138 856
rect 53306 800 53966 856
rect 54134 800 54794 856
rect 54962 800 55530 856
rect 55698 800 56358 856
rect 56526 800 57186 856
rect 57354 800 58014 856
rect 58182 800 58842 856
rect 59010 800 59670 856
rect 59838 800 60406 856
rect 60574 800 61234 856
rect 61402 800 62062 856
rect 62230 800 62890 856
rect 63058 800 63718 856
rect 63886 800 64546 856
rect 64714 800 65282 856
rect 65450 800 66110 856
rect 66278 800 66938 856
rect 67106 800 67766 856
rect 67934 800 68594 856
rect 68762 800 69422 856
rect 69590 800 70250 856
rect 70418 800 70986 856
rect 71154 800 71814 856
rect 71982 800 72642 856
rect 72810 800 73470 856
rect 73638 800 74298 856
rect 74466 800 75126 856
rect 75294 800 75862 856
rect 76030 800 76690 856
rect 76858 800 77518 856
rect 77686 800 78346 856
rect 78514 800 79174 856
rect 79342 800 80002 856
rect 80170 800 80738 856
rect 80906 800 81566 856
rect 81734 800 82394 856
rect 82562 800 83222 856
rect 83390 800 84050 856
rect 84218 800 84878 856
rect 85046 800 85614 856
rect 85782 800 86442 856
rect 86610 800 87270 856
rect 87438 800 88098 856
rect 88266 800 88926 856
rect 89094 800 89754 856
rect 89922 800 90490 856
rect 90658 800 91318 856
rect 91486 800 92146 856
rect 92314 800 92974 856
rect 93142 800 93802 856
rect 93970 800 94630 856
rect 94798 800 95366 856
rect 95534 800 96194 856
rect 96362 800 97022 856
rect 97190 800 97850 856
rect 98018 800 98678 856
rect 98846 800 99506 856
rect 99674 800 100334 856
rect 100502 800 101070 856
rect 101238 800 101898 856
rect 102066 800 102726 856
rect 102894 800 103554 856
rect 103722 800 104382 856
rect 104550 800 105210 856
rect 105378 800 105946 856
rect 106114 800 106774 856
rect 106942 800 107602 856
rect 107770 800 108430 856
rect 108598 800 109258 856
rect 109426 800 110086 856
rect 110254 800 110822 856
rect 110990 800 111650 856
rect 111818 800 112478 856
rect 112646 800 113306 856
rect 113474 800 114134 856
rect 114302 800 114962 856
rect 115130 800 115698 856
rect 115866 800 116526 856
rect 116694 800 117354 856
rect 117522 800 118182 856
rect 118350 800 119010 856
rect 119178 800 119838 856
rect 120006 800 120574 856
rect 120742 800 121402 856
rect 121570 800 122230 856
rect 122398 800 123058 856
rect 123226 800 123886 856
rect 124054 800 124714 856
rect 124882 800 125450 856
rect 125618 800 126278 856
rect 126446 800 127106 856
rect 127274 800 127934 856
rect 128102 800 128762 856
rect 128930 800 129590 856
rect 129758 800 130326 856
rect 130494 800 131154 856
rect 131322 800 131982 856
rect 132150 800 132810 856
rect 132978 800 133638 856
rect 133806 800 134466 856
rect 134634 800 135294 856
rect 135462 800 136030 856
rect 136198 800 136858 856
rect 137026 800 137686 856
rect 137854 800 138514 856
rect 138682 800 139342 856
rect 139510 800 140170 856
rect 140338 800 140906 856
rect 141074 800 141734 856
rect 141902 800 142562 856
rect 142730 800 143390 856
rect 143558 800 144218 856
rect 144386 800 145046 856
rect 145214 800 145782 856
rect 145950 800 146610 856
rect 146778 800 147438 856
rect 147606 800 148266 856
rect 148434 800 149094 856
rect 149262 800 149922 856
rect 150090 800 150658 856
rect 150826 800 151486 856
rect 151654 800 152314 856
rect 152482 800 153142 856
rect 153310 800 153970 856
rect 154138 800 154798 856
rect 154966 800 155534 856
rect 155702 800 156362 856
rect 156530 800 157190 856
rect 157358 800 158018 856
rect 158186 800 158846 856
rect 159014 800 159674 856
rect 159842 800 160410 856
rect 160578 800 161238 856
rect 161406 800 162066 856
rect 162234 800 162894 856
rect 163062 800 163722 856
rect 163890 800 164550 856
rect 164718 800 165286 856
rect 165454 800 166114 856
rect 166282 800 166942 856
rect 167110 800 167770 856
rect 167938 800 168598 856
rect 168766 800 169426 856
rect 169594 800 170254 856
rect 170422 800 170990 856
rect 171158 800 171818 856
rect 171986 800 172646 856
rect 172814 800 173474 856
rect 173642 800 174302 856
rect 174470 800 175130 856
rect 175298 800 175866 856
rect 176034 800 176694 856
rect 176862 800 177522 856
rect 177690 800 178350 856
rect 178518 800 179178 856
rect 179346 800 180006 856
rect 180174 800 180742 856
rect 180910 800 181570 856
rect 181738 800 182398 856
rect 182566 800 183226 856
rect 183394 800 184054 856
rect 184222 800 184882 856
rect 185050 800 185618 856
rect 185786 800 186446 856
rect 186614 800 187274 856
rect 187442 800 188102 856
rect 188270 800 188930 856
rect 189098 800 189758 856
rect 189926 800 190494 856
rect 190662 800 191322 856
rect 191490 800 192150 856
rect 192318 800 192978 856
rect 193146 800 193806 856
rect 193974 800 194634 856
rect 194802 800 195370 856
rect 195538 800 196198 856
rect 196366 800 197026 856
rect 197194 800 197854 856
rect 198022 800 198682 856
rect 198850 800 199510 856
rect 199678 800 200338 856
rect 200506 800 201074 856
rect 201242 800 201902 856
rect 202070 800 202730 856
rect 202898 800 203558 856
rect 203726 800 204386 856
rect 204554 800 205214 856
rect 205382 800 205950 856
rect 206118 800 206778 856
rect 206946 800 207606 856
rect 207774 800 208434 856
rect 208602 800 209262 856
rect 209430 800 210090 856
rect 210258 800 210826 856
rect 210994 800 211654 856
rect 211822 800 212482 856
rect 212650 800 213310 856
rect 213478 800 214138 856
rect 214306 800 214966 856
rect 215134 800 215702 856
rect 215870 800 216530 856
rect 216698 800 217358 856
rect 217526 800 218186 856
rect 218354 800 219014 856
rect 219182 800 219842 856
rect 220010 800 220578 856
rect 220746 800 221406 856
rect 221574 800 222234 856
rect 222402 800 223062 856
rect 223230 800 223890 856
rect 224058 800 224718 856
rect 224886 800 225454 856
rect 225622 800 226282 856
rect 226450 800 227110 856
rect 227278 800 227938 856
rect 228106 800 228766 856
rect 228934 800 229594 856
rect 229762 800 230330 856
rect 230498 800 231158 856
rect 231326 800 231986 856
rect 232154 800 232814 856
rect 232982 800 233642 856
rect 233810 800 234470 856
rect 234638 800 235298 856
rect 235466 800 236034 856
rect 236202 800 236862 856
rect 237030 800 237690 856
rect 237858 800 238518 856
rect 238686 800 239346 856
rect 239514 800 240174 856
rect 240342 800 240910 856
rect 241078 800 241738 856
rect 241906 800 242566 856
rect 242734 800 243394 856
rect 243562 800 244222 856
rect 244390 800 245050 856
rect 245218 800 245786 856
rect 245954 800 246614 856
rect 246782 800 247442 856
rect 247610 800 248270 856
rect 248438 800 249098 856
rect 249266 800 249926 856
rect 250094 800 250662 856
rect 250830 800 251490 856
rect 251658 800 252318 856
rect 252486 800 253146 856
rect 253314 800 253974 856
rect 254142 800 254802 856
rect 254970 800 255538 856
rect 255706 800 256366 856
rect 256534 800 257194 856
rect 257362 800 258022 856
rect 258190 800 258850 856
rect 259018 800 259678 856
rect 259846 800 260414 856
rect 260582 800 261242 856
rect 261410 800 262070 856
rect 262238 800 262898 856
rect 263066 800 263726 856
rect 263894 800 264554 856
rect 264722 800 265290 856
rect 265458 800 266118 856
rect 266286 800 266946 856
rect 267114 800 267774 856
rect 267942 800 268602 856
rect 268770 800 269430 856
rect 269598 800 270258 856
rect 270426 800 270994 856
rect 271162 800 271822 856
rect 271990 800 272650 856
rect 272818 800 273478 856
rect 273646 800 274306 856
rect 274474 800 275134 856
rect 275302 800 275870 856
rect 276038 800 276698 856
rect 276866 800 277526 856
rect 277694 800 278354 856
rect 278522 800 279182 856
rect 279350 800 280010 856
rect 280178 800 280746 856
rect 280914 800 281574 856
rect 281742 800 282402 856
rect 282570 800 283230 856
rect 283398 800 284058 856
rect 284226 800 284886 856
rect 285054 800 285622 856
rect 285790 800 286450 856
rect 286618 800 287278 856
rect 287446 800 288106 856
rect 288274 800 288934 856
rect 289102 800 289762 856
rect 289930 800 290498 856
rect 290666 800 291326 856
rect 291494 800 292154 856
rect 292322 800 292982 856
rect 293150 800 293810 856
rect 293978 800 294638 856
rect 294806 800 295374 856
rect 295542 800 296202 856
rect 296370 800 297030 856
rect 297198 800 297858 856
rect 298026 800 298686 856
rect 298854 800 299514 856
rect 299682 800 300342 856
rect 300510 800 301078 856
rect 301246 800 301906 856
rect 302074 800 302734 856
rect 302902 800 303562 856
rect 303730 800 304390 856
rect 304558 800 305218 856
rect 305386 800 305954 856
rect 306122 800 306782 856
rect 306950 800 307610 856
rect 307778 800 308438 856
rect 308606 800 309266 856
rect 309434 800 310094 856
rect 310262 800 310830 856
rect 310998 800 311658 856
rect 311826 800 312486 856
rect 312654 800 313314 856
rect 313482 800 314142 856
rect 314310 800 314970 856
rect 315138 800 315706 856
rect 315874 800 316534 856
rect 316702 800 317362 856
rect 317530 800 318190 856
rect 318358 800 319018 856
rect 319186 800 319846 856
rect 320014 800 320582 856
rect 320750 800 321410 856
rect 321578 800 322238 856
rect 322406 800 323066 856
rect 323234 800 323894 856
rect 324062 800 324722 856
rect 324890 800 325458 856
rect 325626 800 326286 856
rect 326454 800 327114 856
rect 327282 800 327942 856
rect 328110 800 328770 856
rect 328938 800 329598 856
rect 329766 800 330334 856
rect 330502 800 331162 856
rect 331330 800 331990 856
rect 332158 800 332818 856
rect 332986 800 333646 856
rect 333814 800 334474 856
rect 334642 800 335302 856
rect 335470 800 336038 856
rect 336206 800 336866 856
rect 337034 800 337694 856
rect 337862 800 338522 856
rect 338690 800 339350 856
rect 339518 800 340178 856
rect 340346 800 340914 856
rect 341082 800 341742 856
rect 341910 800 342570 856
rect 342738 800 343398 856
rect 343566 800 344226 856
rect 344394 800 345054 856
rect 345222 800 345790 856
rect 345958 800 346618 856
rect 346786 800 347446 856
rect 347614 800 348274 856
rect 348442 800 349102 856
rect 349270 800 349930 856
rect 350098 800 350666 856
rect 350834 800 351494 856
rect 351662 800 352322 856
rect 352490 800 353150 856
rect 353318 800 353978 856
rect 354146 800 354806 856
rect 354974 800 355542 856
rect 355710 800 356370 856
rect 356538 800 357198 856
rect 357366 800 358026 856
rect 358194 800 358854 856
rect 359022 800 359682 856
rect 359850 800 360418 856
rect 360586 800 361246 856
rect 361414 800 362074 856
rect 362242 800 362902 856
rect 363070 800 363730 856
rect 363898 800 364558 856
rect 364726 800 365294 856
rect 365462 800 366122 856
rect 366290 800 366950 856
rect 367118 800 367778 856
rect 367946 800 368606 856
rect 368774 800 369434 856
rect 369602 800 370262 856
rect 370430 800 370998 856
rect 371166 800 371826 856
rect 371994 800 372654 856
rect 372822 800 373482 856
rect 373650 800 374310 856
rect 374478 800 375138 856
rect 375306 800 375874 856
rect 376042 800 376702 856
rect 376870 800 377530 856
rect 377698 800 378358 856
rect 378526 800 379186 856
rect 379354 800 380014 856
rect 380182 800 380750 856
rect 380918 800 381578 856
rect 381746 800 382406 856
rect 382574 800 383234 856
rect 383402 800 384062 856
rect 384230 800 384890 856
rect 385058 800 385626 856
rect 385794 800 386454 856
rect 386622 800 387282 856
rect 387450 800 388110 856
rect 388278 800 388938 856
rect 389106 800 389766 856
rect 389934 800 390502 856
rect 390670 800 391330 856
rect 391498 800 392158 856
rect 392326 800 392986 856
rect 393154 800 393814 856
rect 393982 800 394642 856
rect 394810 800 395378 856
rect 395546 800 396206 856
rect 396374 800 397034 856
<< metal3 >>
rect 0 374960 800 375080
rect 0 124992 800 125112
rect 399200 249976 400000 250096
<< obsm3 >>
rect 2405 2143 388528 497793
<< metal4 >>
rect 4208 2128 4528 497808
rect 19568 2128 19888 497808
rect 34928 2128 35248 497808
rect 50288 2128 50608 497808
rect 65648 2128 65968 497808
rect 81008 2128 81328 497808
rect 96368 2128 96688 497808
rect 111728 2128 112048 497808
rect 127088 2128 127408 497808
rect 142448 2128 142768 497808
rect 157808 2128 158128 497808
rect 173168 2128 173488 497808
rect 188528 2128 188848 497808
rect 203888 2128 204208 497808
rect 219248 2128 219568 497808
rect 234608 2128 234928 497808
rect 249968 2128 250288 497808
rect 265328 2128 265648 497808
rect 280688 2128 281008 497808
rect 296048 2128 296368 497808
rect 311408 2128 311728 497808
rect 326768 2128 327088 497808
rect 342128 2128 342448 497808
rect 357488 2128 357808 497808
rect 372848 2128 373168 497808
rect 388208 2128 388528 497808
<< labels >>
rlabel metal2 s 1674 499200 1730 500000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 104162 499200 104218 500000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 114466 499200 114522 500000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 124678 499200 124734 500000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 134982 499200 135038 500000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 145194 499200 145250 500000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 155498 499200 155554 500000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 165710 499200 165766 500000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 176014 499200 176070 500000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 186226 499200 186282 500000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 196530 499200 196586 500000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 11886 499200 11942 500000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 206742 499200 206798 500000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 217046 499200 217102 500000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 227258 499200 227314 500000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 237562 499200 237618 500000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 247774 499200 247830 500000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 258078 499200 258134 500000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 268290 499200 268346 500000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 278594 499200 278650 500000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 288806 499200 288862 500000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 299110 499200 299166 500000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 22098 499200 22154 500000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 309322 499200 309378 500000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 319626 499200 319682 500000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 329838 499200 329894 500000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 340142 499200 340198 500000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 350354 499200 350410 500000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 360658 499200 360714 500000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 370870 499200 370926 500000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 381174 499200 381230 500000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 32402 499200 32458 500000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 42614 499200 42670 500000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 52918 499200 52974 500000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 63130 499200 63186 500000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 73434 499200 73490 500000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 83646 499200 83702 500000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 93950 499200 94006 500000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 5078 499200 5134 500000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 107658 499200 107714 500000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 117870 499200 117926 500000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 128174 499200 128230 500000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 138386 499200 138442 500000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 148598 499200 148654 500000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 158902 499200 158958 500000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 169114 499200 169170 500000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 179418 499200 179474 500000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 189630 499200 189686 500000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 199934 499200 199990 500000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 15290 499200 15346 500000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 210146 499200 210202 500000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 220450 499200 220506 500000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 230662 499200 230718 500000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 240966 499200 241022 500000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 251178 499200 251234 500000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 261482 499200 261538 500000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 271694 499200 271750 500000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 281998 499200 282054 500000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 292210 499200 292266 500000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 302514 499200 302570 500000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 25594 499200 25650 500000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 312726 499200 312782 500000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 323030 499200 323086 500000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 333242 499200 333298 500000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 343546 499200 343602 500000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 353758 499200 353814 500000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 364062 499200 364118 500000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 374274 499200 374330 500000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 384578 499200 384634 500000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 35806 499200 35862 500000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 46110 499200 46166 500000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 56322 499200 56378 500000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 66626 499200 66682 500000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 76838 499200 76894 500000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 87142 499200 87198 500000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 97354 499200 97410 500000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 8482 499200 8538 500000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 111062 499200 111118 500000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 121274 499200 121330 500000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 131578 499200 131634 500000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 141790 499200 141846 500000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 152094 499200 152150 500000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 162306 499200 162362 500000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 172610 499200 172666 500000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 182822 499200 182878 500000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 193126 499200 193182 500000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 203338 499200 203394 500000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 18694 499200 18750 500000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 213642 499200 213698 500000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 223854 499200 223910 500000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 234158 499200 234214 500000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 244370 499200 244426 500000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 254674 499200 254730 500000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 264886 499200 264942 500000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 275098 499200 275154 500000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 285402 499200 285458 500000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 295614 499200 295670 500000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 305918 499200 305974 500000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 28998 499200 29054 500000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 316130 499200 316186 500000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 326434 499200 326490 500000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 336646 499200 336702 500000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 346950 499200 347006 500000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 357162 499200 357218 500000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 367466 499200 367522 500000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 377678 499200 377734 500000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 387982 499200 388038 500000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 39210 499200 39266 500000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 49514 499200 49570 500000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 59726 499200 59782 500000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 70030 499200 70086 500000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 80242 499200 80298 500000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 90546 499200 90602 500000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 100758 499200 100814 500000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 86498 0 86554 800 6 la_data_in[0]
port 115 nsew signal input
rlabel metal2 s 330390 0 330446 800 6 la_data_in[100]
port 116 nsew signal input
rlabel metal2 s 332874 0 332930 800 6 la_data_in[101]
port 117 nsew signal input
rlabel metal2 s 335358 0 335414 800 6 la_data_in[102]
port 118 nsew signal input
rlabel metal2 s 337750 0 337806 800 6 la_data_in[103]
port 119 nsew signal input
rlabel metal2 s 340234 0 340290 800 6 la_data_in[104]
port 120 nsew signal input
rlabel metal2 s 342626 0 342682 800 6 la_data_in[105]
port 121 nsew signal input
rlabel metal2 s 345110 0 345166 800 6 la_data_in[106]
port 122 nsew signal input
rlabel metal2 s 347502 0 347558 800 6 la_data_in[107]
port 123 nsew signal input
rlabel metal2 s 349986 0 350042 800 6 la_data_in[108]
port 124 nsew signal input
rlabel metal2 s 352378 0 352434 800 6 la_data_in[109]
port 125 nsew signal input
rlabel metal2 s 110878 0 110934 800 6 la_data_in[10]
port 126 nsew signal input
rlabel metal2 s 354862 0 354918 800 6 la_data_in[110]
port 127 nsew signal input
rlabel metal2 s 357254 0 357310 800 6 la_data_in[111]
port 128 nsew signal input
rlabel metal2 s 359738 0 359794 800 6 la_data_in[112]
port 129 nsew signal input
rlabel metal2 s 362130 0 362186 800 6 la_data_in[113]
port 130 nsew signal input
rlabel metal2 s 364614 0 364670 800 6 la_data_in[114]
port 131 nsew signal input
rlabel metal2 s 367006 0 367062 800 6 la_data_in[115]
port 132 nsew signal input
rlabel metal2 s 369490 0 369546 800 6 la_data_in[116]
port 133 nsew signal input
rlabel metal2 s 371882 0 371938 800 6 la_data_in[117]
port 134 nsew signal input
rlabel metal2 s 374366 0 374422 800 6 la_data_in[118]
port 135 nsew signal input
rlabel metal2 s 376758 0 376814 800 6 la_data_in[119]
port 136 nsew signal input
rlabel metal2 s 113362 0 113418 800 6 la_data_in[11]
port 137 nsew signal input
rlabel metal2 s 379242 0 379298 800 6 la_data_in[120]
port 138 nsew signal input
rlabel metal2 s 381634 0 381690 800 6 la_data_in[121]
port 139 nsew signal input
rlabel metal2 s 384118 0 384174 800 6 la_data_in[122]
port 140 nsew signal input
rlabel metal2 s 386510 0 386566 800 6 la_data_in[123]
port 141 nsew signal input
rlabel metal2 s 388994 0 389050 800 6 la_data_in[124]
port 142 nsew signal input
rlabel metal2 s 391386 0 391442 800 6 la_data_in[125]
port 143 nsew signal input
rlabel metal2 s 393870 0 393926 800 6 la_data_in[126]
port 144 nsew signal input
rlabel metal2 s 396262 0 396318 800 6 la_data_in[127]
port 145 nsew signal input
rlabel metal2 s 115754 0 115810 800 6 la_data_in[12]
port 146 nsew signal input
rlabel metal2 s 118238 0 118294 800 6 la_data_in[13]
port 147 nsew signal input
rlabel metal2 s 120630 0 120686 800 6 la_data_in[14]
port 148 nsew signal input
rlabel metal2 s 123114 0 123170 800 6 la_data_in[15]
port 149 nsew signal input
rlabel metal2 s 125506 0 125562 800 6 la_data_in[16]
port 150 nsew signal input
rlabel metal2 s 127990 0 128046 800 6 la_data_in[17]
port 151 nsew signal input
rlabel metal2 s 130382 0 130438 800 6 la_data_in[18]
port 152 nsew signal input
rlabel metal2 s 132866 0 132922 800 6 la_data_in[19]
port 153 nsew signal input
rlabel metal2 s 88982 0 89038 800 6 la_data_in[1]
port 154 nsew signal input
rlabel metal2 s 135350 0 135406 800 6 la_data_in[20]
port 155 nsew signal input
rlabel metal2 s 137742 0 137798 800 6 la_data_in[21]
port 156 nsew signal input
rlabel metal2 s 140226 0 140282 800 6 la_data_in[22]
port 157 nsew signal input
rlabel metal2 s 142618 0 142674 800 6 la_data_in[23]
port 158 nsew signal input
rlabel metal2 s 145102 0 145158 800 6 la_data_in[24]
port 159 nsew signal input
rlabel metal2 s 147494 0 147550 800 6 la_data_in[25]
port 160 nsew signal input
rlabel metal2 s 149978 0 150034 800 6 la_data_in[26]
port 161 nsew signal input
rlabel metal2 s 152370 0 152426 800 6 la_data_in[27]
port 162 nsew signal input
rlabel metal2 s 154854 0 154910 800 6 la_data_in[28]
port 163 nsew signal input
rlabel metal2 s 157246 0 157302 800 6 la_data_in[29]
port 164 nsew signal input
rlabel metal2 s 91374 0 91430 800 6 la_data_in[2]
port 165 nsew signal input
rlabel metal2 s 159730 0 159786 800 6 la_data_in[30]
port 166 nsew signal input
rlabel metal2 s 162122 0 162178 800 6 la_data_in[31]
port 167 nsew signal input
rlabel metal2 s 164606 0 164662 800 6 la_data_in[32]
port 168 nsew signal input
rlabel metal2 s 166998 0 167054 800 6 la_data_in[33]
port 169 nsew signal input
rlabel metal2 s 169482 0 169538 800 6 la_data_in[34]
port 170 nsew signal input
rlabel metal2 s 171874 0 171930 800 6 la_data_in[35]
port 171 nsew signal input
rlabel metal2 s 174358 0 174414 800 6 la_data_in[36]
port 172 nsew signal input
rlabel metal2 s 176750 0 176806 800 6 la_data_in[37]
port 173 nsew signal input
rlabel metal2 s 179234 0 179290 800 6 la_data_in[38]
port 174 nsew signal input
rlabel metal2 s 181626 0 181682 800 6 la_data_in[39]
port 175 nsew signal input
rlabel metal2 s 93858 0 93914 800 6 la_data_in[3]
port 176 nsew signal input
rlabel metal2 s 184110 0 184166 800 6 la_data_in[40]
port 177 nsew signal input
rlabel metal2 s 186502 0 186558 800 6 la_data_in[41]
port 178 nsew signal input
rlabel metal2 s 188986 0 189042 800 6 la_data_in[42]
port 179 nsew signal input
rlabel metal2 s 191378 0 191434 800 6 la_data_in[43]
port 180 nsew signal input
rlabel metal2 s 193862 0 193918 800 6 la_data_in[44]
port 181 nsew signal input
rlabel metal2 s 196254 0 196310 800 6 la_data_in[45]
port 182 nsew signal input
rlabel metal2 s 198738 0 198794 800 6 la_data_in[46]
port 183 nsew signal input
rlabel metal2 s 201130 0 201186 800 6 la_data_in[47]
port 184 nsew signal input
rlabel metal2 s 203614 0 203670 800 6 la_data_in[48]
port 185 nsew signal input
rlabel metal2 s 206006 0 206062 800 6 la_data_in[49]
port 186 nsew signal input
rlabel metal2 s 96250 0 96306 800 6 la_data_in[4]
port 187 nsew signal input
rlabel metal2 s 208490 0 208546 800 6 la_data_in[50]
port 188 nsew signal input
rlabel metal2 s 210882 0 210938 800 6 la_data_in[51]
port 189 nsew signal input
rlabel metal2 s 213366 0 213422 800 6 la_data_in[52]
port 190 nsew signal input
rlabel metal2 s 215758 0 215814 800 6 la_data_in[53]
port 191 nsew signal input
rlabel metal2 s 218242 0 218298 800 6 la_data_in[54]
port 192 nsew signal input
rlabel metal2 s 220634 0 220690 800 6 la_data_in[55]
port 193 nsew signal input
rlabel metal2 s 223118 0 223174 800 6 la_data_in[56]
port 194 nsew signal input
rlabel metal2 s 225510 0 225566 800 6 la_data_in[57]
port 195 nsew signal input
rlabel metal2 s 227994 0 228050 800 6 la_data_in[58]
port 196 nsew signal input
rlabel metal2 s 230386 0 230442 800 6 la_data_in[59]
port 197 nsew signal input
rlabel metal2 s 98734 0 98790 800 6 la_data_in[5]
port 198 nsew signal input
rlabel metal2 s 232870 0 232926 800 6 la_data_in[60]
port 199 nsew signal input
rlabel metal2 s 235354 0 235410 800 6 la_data_in[61]
port 200 nsew signal input
rlabel metal2 s 237746 0 237802 800 6 la_data_in[62]
port 201 nsew signal input
rlabel metal2 s 240230 0 240286 800 6 la_data_in[63]
port 202 nsew signal input
rlabel metal2 s 242622 0 242678 800 6 la_data_in[64]
port 203 nsew signal input
rlabel metal2 s 245106 0 245162 800 6 la_data_in[65]
port 204 nsew signal input
rlabel metal2 s 247498 0 247554 800 6 la_data_in[66]
port 205 nsew signal input
rlabel metal2 s 249982 0 250038 800 6 la_data_in[67]
port 206 nsew signal input
rlabel metal2 s 252374 0 252430 800 6 la_data_in[68]
port 207 nsew signal input
rlabel metal2 s 254858 0 254914 800 6 la_data_in[69]
port 208 nsew signal input
rlabel metal2 s 101126 0 101182 800 6 la_data_in[6]
port 209 nsew signal input
rlabel metal2 s 257250 0 257306 800 6 la_data_in[70]
port 210 nsew signal input
rlabel metal2 s 259734 0 259790 800 6 la_data_in[71]
port 211 nsew signal input
rlabel metal2 s 262126 0 262182 800 6 la_data_in[72]
port 212 nsew signal input
rlabel metal2 s 264610 0 264666 800 6 la_data_in[73]
port 213 nsew signal input
rlabel metal2 s 267002 0 267058 800 6 la_data_in[74]
port 214 nsew signal input
rlabel metal2 s 269486 0 269542 800 6 la_data_in[75]
port 215 nsew signal input
rlabel metal2 s 271878 0 271934 800 6 la_data_in[76]
port 216 nsew signal input
rlabel metal2 s 274362 0 274418 800 6 la_data_in[77]
port 217 nsew signal input
rlabel metal2 s 276754 0 276810 800 6 la_data_in[78]
port 218 nsew signal input
rlabel metal2 s 279238 0 279294 800 6 la_data_in[79]
port 219 nsew signal input
rlabel metal2 s 103610 0 103666 800 6 la_data_in[7]
port 220 nsew signal input
rlabel metal2 s 281630 0 281686 800 6 la_data_in[80]
port 221 nsew signal input
rlabel metal2 s 284114 0 284170 800 6 la_data_in[81]
port 222 nsew signal input
rlabel metal2 s 286506 0 286562 800 6 la_data_in[82]
port 223 nsew signal input
rlabel metal2 s 288990 0 289046 800 6 la_data_in[83]
port 224 nsew signal input
rlabel metal2 s 291382 0 291438 800 6 la_data_in[84]
port 225 nsew signal input
rlabel metal2 s 293866 0 293922 800 6 la_data_in[85]
port 226 nsew signal input
rlabel metal2 s 296258 0 296314 800 6 la_data_in[86]
port 227 nsew signal input
rlabel metal2 s 298742 0 298798 800 6 la_data_in[87]
port 228 nsew signal input
rlabel metal2 s 301134 0 301190 800 6 la_data_in[88]
port 229 nsew signal input
rlabel metal2 s 303618 0 303674 800 6 la_data_in[89]
port 230 nsew signal input
rlabel metal2 s 106002 0 106058 800 6 la_data_in[8]
port 231 nsew signal input
rlabel metal2 s 306010 0 306066 800 6 la_data_in[90]
port 232 nsew signal input
rlabel metal2 s 308494 0 308550 800 6 la_data_in[91]
port 233 nsew signal input
rlabel metal2 s 310886 0 310942 800 6 la_data_in[92]
port 234 nsew signal input
rlabel metal2 s 313370 0 313426 800 6 la_data_in[93]
port 235 nsew signal input
rlabel metal2 s 315762 0 315818 800 6 la_data_in[94]
port 236 nsew signal input
rlabel metal2 s 318246 0 318302 800 6 la_data_in[95]
port 237 nsew signal input
rlabel metal2 s 320638 0 320694 800 6 la_data_in[96]
port 238 nsew signal input
rlabel metal2 s 323122 0 323178 800 6 la_data_in[97]
port 239 nsew signal input
rlabel metal2 s 325514 0 325570 800 6 la_data_in[98]
port 240 nsew signal input
rlabel metal2 s 327998 0 328054 800 6 la_data_in[99]
port 241 nsew signal input
rlabel metal2 s 108486 0 108542 800 6 la_data_in[9]
port 242 nsew signal input
rlabel metal2 s 87326 0 87382 800 6 la_data_out[0]
port 243 nsew signal output
rlabel metal2 s 331218 0 331274 800 6 la_data_out[100]
port 244 nsew signal output
rlabel metal2 s 333702 0 333758 800 6 la_data_out[101]
port 245 nsew signal output
rlabel metal2 s 336094 0 336150 800 6 la_data_out[102]
port 246 nsew signal output
rlabel metal2 s 338578 0 338634 800 6 la_data_out[103]
port 247 nsew signal output
rlabel metal2 s 340970 0 341026 800 6 la_data_out[104]
port 248 nsew signal output
rlabel metal2 s 343454 0 343510 800 6 la_data_out[105]
port 249 nsew signal output
rlabel metal2 s 345846 0 345902 800 6 la_data_out[106]
port 250 nsew signal output
rlabel metal2 s 348330 0 348386 800 6 la_data_out[107]
port 251 nsew signal output
rlabel metal2 s 350722 0 350778 800 6 la_data_out[108]
port 252 nsew signal output
rlabel metal2 s 353206 0 353262 800 6 la_data_out[109]
port 253 nsew signal output
rlabel metal2 s 111706 0 111762 800 6 la_data_out[10]
port 254 nsew signal output
rlabel metal2 s 355598 0 355654 800 6 la_data_out[110]
port 255 nsew signal output
rlabel metal2 s 358082 0 358138 800 6 la_data_out[111]
port 256 nsew signal output
rlabel metal2 s 360474 0 360530 800 6 la_data_out[112]
port 257 nsew signal output
rlabel metal2 s 362958 0 363014 800 6 la_data_out[113]
port 258 nsew signal output
rlabel metal2 s 365350 0 365406 800 6 la_data_out[114]
port 259 nsew signal output
rlabel metal2 s 367834 0 367890 800 6 la_data_out[115]
port 260 nsew signal output
rlabel metal2 s 370318 0 370374 800 6 la_data_out[116]
port 261 nsew signal output
rlabel metal2 s 372710 0 372766 800 6 la_data_out[117]
port 262 nsew signal output
rlabel metal2 s 375194 0 375250 800 6 la_data_out[118]
port 263 nsew signal output
rlabel metal2 s 377586 0 377642 800 6 la_data_out[119]
port 264 nsew signal output
rlabel metal2 s 114190 0 114246 800 6 la_data_out[11]
port 265 nsew signal output
rlabel metal2 s 380070 0 380126 800 6 la_data_out[120]
port 266 nsew signal output
rlabel metal2 s 382462 0 382518 800 6 la_data_out[121]
port 267 nsew signal output
rlabel metal2 s 384946 0 385002 800 6 la_data_out[122]
port 268 nsew signal output
rlabel metal2 s 387338 0 387394 800 6 la_data_out[123]
port 269 nsew signal output
rlabel metal2 s 389822 0 389878 800 6 la_data_out[124]
port 270 nsew signal output
rlabel metal2 s 392214 0 392270 800 6 la_data_out[125]
port 271 nsew signal output
rlabel metal2 s 394698 0 394754 800 6 la_data_out[126]
port 272 nsew signal output
rlabel metal2 s 397090 0 397146 800 6 la_data_out[127]
port 273 nsew signal output
rlabel metal2 s 116582 0 116638 800 6 la_data_out[12]
port 274 nsew signal output
rlabel metal2 s 119066 0 119122 800 6 la_data_out[13]
port 275 nsew signal output
rlabel metal2 s 121458 0 121514 800 6 la_data_out[14]
port 276 nsew signal output
rlabel metal2 s 123942 0 123998 800 6 la_data_out[15]
port 277 nsew signal output
rlabel metal2 s 126334 0 126390 800 6 la_data_out[16]
port 278 nsew signal output
rlabel metal2 s 128818 0 128874 800 6 la_data_out[17]
port 279 nsew signal output
rlabel metal2 s 131210 0 131266 800 6 la_data_out[18]
port 280 nsew signal output
rlabel metal2 s 133694 0 133750 800 6 la_data_out[19]
port 281 nsew signal output
rlabel metal2 s 89810 0 89866 800 6 la_data_out[1]
port 282 nsew signal output
rlabel metal2 s 136086 0 136142 800 6 la_data_out[20]
port 283 nsew signal output
rlabel metal2 s 138570 0 138626 800 6 la_data_out[21]
port 284 nsew signal output
rlabel metal2 s 140962 0 141018 800 6 la_data_out[22]
port 285 nsew signal output
rlabel metal2 s 143446 0 143502 800 6 la_data_out[23]
port 286 nsew signal output
rlabel metal2 s 145838 0 145894 800 6 la_data_out[24]
port 287 nsew signal output
rlabel metal2 s 148322 0 148378 800 6 la_data_out[25]
port 288 nsew signal output
rlabel metal2 s 150714 0 150770 800 6 la_data_out[26]
port 289 nsew signal output
rlabel metal2 s 153198 0 153254 800 6 la_data_out[27]
port 290 nsew signal output
rlabel metal2 s 155590 0 155646 800 6 la_data_out[28]
port 291 nsew signal output
rlabel metal2 s 158074 0 158130 800 6 la_data_out[29]
port 292 nsew signal output
rlabel metal2 s 92202 0 92258 800 6 la_data_out[2]
port 293 nsew signal output
rlabel metal2 s 160466 0 160522 800 6 la_data_out[30]
port 294 nsew signal output
rlabel metal2 s 162950 0 163006 800 6 la_data_out[31]
port 295 nsew signal output
rlabel metal2 s 165342 0 165398 800 6 la_data_out[32]
port 296 nsew signal output
rlabel metal2 s 167826 0 167882 800 6 la_data_out[33]
port 297 nsew signal output
rlabel metal2 s 170310 0 170366 800 6 la_data_out[34]
port 298 nsew signal output
rlabel metal2 s 172702 0 172758 800 6 la_data_out[35]
port 299 nsew signal output
rlabel metal2 s 175186 0 175242 800 6 la_data_out[36]
port 300 nsew signal output
rlabel metal2 s 177578 0 177634 800 6 la_data_out[37]
port 301 nsew signal output
rlabel metal2 s 180062 0 180118 800 6 la_data_out[38]
port 302 nsew signal output
rlabel metal2 s 182454 0 182510 800 6 la_data_out[39]
port 303 nsew signal output
rlabel metal2 s 94686 0 94742 800 6 la_data_out[3]
port 304 nsew signal output
rlabel metal2 s 184938 0 184994 800 6 la_data_out[40]
port 305 nsew signal output
rlabel metal2 s 187330 0 187386 800 6 la_data_out[41]
port 306 nsew signal output
rlabel metal2 s 189814 0 189870 800 6 la_data_out[42]
port 307 nsew signal output
rlabel metal2 s 192206 0 192262 800 6 la_data_out[43]
port 308 nsew signal output
rlabel metal2 s 194690 0 194746 800 6 la_data_out[44]
port 309 nsew signal output
rlabel metal2 s 197082 0 197138 800 6 la_data_out[45]
port 310 nsew signal output
rlabel metal2 s 199566 0 199622 800 6 la_data_out[46]
port 311 nsew signal output
rlabel metal2 s 201958 0 202014 800 6 la_data_out[47]
port 312 nsew signal output
rlabel metal2 s 204442 0 204498 800 6 la_data_out[48]
port 313 nsew signal output
rlabel metal2 s 206834 0 206890 800 6 la_data_out[49]
port 314 nsew signal output
rlabel metal2 s 97078 0 97134 800 6 la_data_out[4]
port 315 nsew signal output
rlabel metal2 s 209318 0 209374 800 6 la_data_out[50]
port 316 nsew signal output
rlabel metal2 s 211710 0 211766 800 6 la_data_out[51]
port 317 nsew signal output
rlabel metal2 s 214194 0 214250 800 6 la_data_out[52]
port 318 nsew signal output
rlabel metal2 s 216586 0 216642 800 6 la_data_out[53]
port 319 nsew signal output
rlabel metal2 s 219070 0 219126 800 6 la_data_out[54]
port 320 nsew signal output
rlabel metal2 s 221462 0 221518 800 6 la_data_out[55]
port 321 nsew signal output
rlabel metal2 s 223946 0 224002 800 6 la_data_out[56]
port 322 nsew signal output
rlabel metal2 s 226338 0 226394 800 6 la_data_out[57]
port 323 nsew signal output
rlabel metal2 s 228822 0 228878 800 6 la_data_out[58]
port 324 nsew signal output
rlabel metal2 s 231214 0 231270 800 6 la_data_out[59]
port 325 nsew signal output
rlabel metal2 s 99562 0 99618 800 6 la_data_out[5]
port 326 nsew signal output
rlabel metal2 s 233698 0 233754 800 6 la_data_out[60]
port 327 nsew signal output
rlabel metal2 s 236090 0 236146 800 6 la_data_out[61]
port 328 nsew signal output
rlabel metal2 s 238574 0 238630 800 6 la_data_out[62]
port 329 nsew signal output
rlabel metal2 s 240966 0 241022 800 6 la_data_out[63]
port 330 nsew signal output
rlabel metal2 s 243450 0 243506 800 6 la_data_out[64]
port 331 nsew signal output
rlabel metal2 s 245842 0 245898 800 6 la_data_out[65]
port 332 nsew signal output
rlabel metal2 s 248326 0 248382 800 6 la_data_out[66]
port 333 nsew signal output
rlabel metal2 s 250718 0 250774 800 6 la_data_out[67]
port 334 nsew signal output
rlabel metal2 s 253202 0 253258 800 6 la_data_out[68]
port 335 nsew signal output
rlabel metal2 s 255594 0 255650 800 6 la_data_out[69]
port 336 nsew signal output
rlabel metal2 s 101954 0 102010 800 6 la_data_out[6]
port 337 nsew signal output
rlabel metal2 s 258078 0 258134 800 6 la_data_out[70]
port 338 nsew signal output
rlabel metal2 s 260470 0 260526 800 6 la_data_out[71]
port 339 nsew signal output
rlabel metal2 s 262954 0 263010 800 6 la_data_out[72]
port 340 nsew signal output
rlabel metal2 s 265346 0 265402 800 6 la_data_out[73]
port 341 nsew signal output
rlabel metal2 s 267830 0 267886 800 6 la_data_out[74]
port 342 nsew signal output
rlabel metal2 s 270314 0 270370 800 6 la_data_out[75]
port 343 nsew signal output
rlabel metal2 s 272706 0 272762 800 6 la_data_out[76]
port 344 nsew signal output
rlabel metal2 s 275190 0 275246 800 6 la_data_out[77]
port 345 nsew signal output
rlabel metal2 s 277582 0 277638 800 6 la_data_out[78]
port 346 nsew signal output
rlabel metal2 s 280066 0 280122 800 6 la_data_out[79]
port 347 nsew signal output
rlabel metal2 s 104438 0 104494 800 6 la_data_out[7]
port 348 nsew signal output
rlabel metal2 s 282458 0 282514 800 6 la_data_out[80]
port 349 nsew signal output
rlabel metal2 s 284942 0 284998 800 6 la_data_out[81]
port 350 nsew signal output
rlabel metal2 s 287334 0 287390 800 6 la_data_out[82]
port 351 nsew signal output
rlabel metal2 s 289818 0 289874 800 6 la_data_out[83]
port 352 nsew signal output
rlabel metal2 s 292210 0 292266 800 6 la_data_out[84]
port 353 nsew signal output
rlabel metal2 s 294694 0 294750 800 6 la_data_out[85]
port 354 nsew signal output
rlabel metal2 s 297086 0 297142 800 6 la_data_out[86]
port 355 nsew signal output
rlabel metal2 s 299570 0 299626 800 6 la_data_out[87]
port 356 nsew signal output
rlabel metal2 s 301962 0 302018 800 6 la_data_out[88]
port 357 nsew signal output
rlabel metal2 s 304446 0 304502 800 6 la_data_out[89]
port 358 nsew signal output
rlabel metal2 s 106830 0 106886 800 6 la_data_out[8]
port 359 nsew signal output
rlabel metal2 s 306838 0 306894 800 6 la_data_out[90]
port 360 nsew signal output
rlabel metal2 s 309322 0 309378 800 6 la_data_out[91]
port 361 nsew signal output
rlabel metal2 s 311714 0 311770 800 6 la_data_out[92]
port 362 nsew signal output
rlabel metal2 s 314198 0 314254 800 6 la_data_out[93]
port 363 nsew signal output
rlabel metal2 s 316590 0 316646 800 6 la_data_out[94]
port 364 nsew signal output
rlabel metal2 s 319074 0 319130 800 6 la_data_out[95]
port 365 nsew signal output
rlabel metal2 s 321466 0 321522 800 6 la_data_out[96]
port 366 nsew signal output
rlabel metal2 s 323950 0 324006 800 6 la_data_out[97]
port 367 nsew signal output
rlabel metal2 s 326342 0 326398 800 6 la_data_out[98]
port 368 nsew signal output
rlabel metal2 s 328826 0 328882 800 6 la_data_out[99]
port 369 nsew signal output
rlabel metal2 s 109314 0 109370 800 6 la_data_out[9]
port 370 nsew signal output
rlabel metal2 s 88154 0 88210 800 6 la_oen[0]
port 371 nsew signal input
rlabel metal2 s 332046 0 332102 800 6 la_oen[100]
port 372 nsew signal input
rlabel metal2 s 334530 0 334586 800 6 la_oen[101]
port 373 nsew signal input
rlabel metal2 s 336922 0 336978 800 6 la_oen[102]
port 374 nsew signal input
rlabel metal2 s 339406 0 339462 800 6 la_oen[103]
port 375 nsew signal input
rlabel metal2 s 341798 0 341854 800 6 la_oen[104]
port 376 nsew signal input
rlabel metal2 s 344282 0 344338 800 6 la_oen[105]
port 377 nsew signal input
rlabel metal2 s 346674 0 346730 800 6 la_oen[106]
port 378 nsew signal input
rlabel metal2 s 349158 0 349214 800 6 la_oen[107]
port 379 nsew signal input
rlabel metal2 s 351550 0 351606 800 6 la_oen[108]
port 380 nsew signal input
rlabel metal2 s 354034 0 354090 800 6 la_oen[109]
port 381 nsew signal input
rlabel metal2 s 112534 0 112590 800 6 la_oen[10]
port 382 nsew signal input
rlabel metal2 s 356426 0 356482 800 6 la_oen[110]
port 383 nsew signal input
rlabel metal2 s 358910 0 358966 800 6 la_oen[111]
port 384 nsew signal input
rlabel metal2 s 361302 0 361358 800 6 la_oen[112]
port 385 nsew signal input
rlabel metal2 s 363786 0 363842 800 6 la_oen[113]
port 386 nsew signal input
rlabel metal2 s 366178 0 366234 800 6 la_oen[114]
port 387 nsew signal input
rlabel metal2 s 368662 0 368718 800 6 la_oen[115]
port 388 nsew signal input
rlabel metal2 s 371054 0 371110 800 6 la_oen[116]
port 389 nsew signal input
rlabel metal2 s 373538 0 373594 800 6 la_oen[117]
port 390 nsew signal input
rlabel metal2 s 375930 0 375986 800 6 la_oen[118]
port 391 nsew signal input
rlabel metal2 s 378414 0 378470 800 6 la_oen[119]
port 392 nsew signal input
rlabel metal2 s 115018 0 115074 800 6 la_oen[11]
port 393 nsew signal input
rlabel metal2 s 380806 0 380862 800 6 la_oen[120]
port 394 nsew signal input
rlabel metal2 s 383290 0 383346 800 6 la_oen[121]
port 395 nsew signal input
rlabel metal2 s 385682 0 385738 800 6 la_oen[122]
port 396 nsew signal input
rlabel metal2 s 388166 0 388222 800 6 la_oen[123]
port 397 nsew signal input
rlabel metal2 s 390558 0 390614 800 6 la_oen[124]
port 398 nsew signal input
rlabel metal2 s 393042 0 393098 800 6 la_oen[125]
port 399 nsew signal input
rlabel metal2 s 395434 0 395490 800 6 la_oen[126]
port 400 nsew signal input
rlabel metal2 s 397918 0 397974 800 6 la_oen[127]
port 401 nsew signal input
rlabel metal2 s 117410 0 117466 800 6 la_oen[12]
port 402 nsew signal input
rlabel metal2 s 119894 0 119950 800 6 la_oen[13]
port 403 nsew signal input
rlabel metal2 s 122286 0 122342 800 6 la_oen[14]
port 404 nsew signal input
rlabel metal2 s 124770 0 124826 800 6 la_oen[15]
port 405 nsew signal input
rlabel metal2 s 127162 0 127218 800 6 la_oen[16]
port 406 nsew signal input
rlabel metal2 s 129646 0 129702 800 6 la_oen[17]
port 407 nsew signal input
rlabel metal2 s 132038 0 132094 800 6 la_oen[18]
port 408 nsew signal input
rlabel metal2 s 134522 0 134578 800 6 la_oen[19]
port 409 nsew signal input
rlabel metal2 s 90546 0 90602 800 6 la_oen[1]
port 410 nsew signal input
rlabel metal2 s 136914 0 136970 800 6 la_oen[20]
port 411 nsew signal input
rlabel metal2 s 139398 0 139454 800 6 la_oen[21]
port 412 nsew signal input
rlabel metal2 s 141790 0 141846 800 6 la_oen[22]
port 413 nsew signal input
rlabel metal2 s 144274 0 144330 800 6 la_oen[23]
port 414 nsew signal input
rlabel metal2 s 146666 0 146722 800 6 la_oen[24]
port 415 nsew signal input
rlabel metal2 s 149150 0 149206 800 6 la_oen[25]
port 416 nsew signal input
rlabel metal2 s 151542 0 151598 800 6 la_oen[26]
port 417 nsew signal input
rlabel metal2 s 154026 0 154082 800 6 la_oen[27]
port 418 nsew signal input
rlabel metal2 s 156418 0 156474 800 6 la_oen[28]
port 419 nsew signal input
rlabel metal2 s 158902 0 158958 800 6 la_oen[29]
port 420 nsew signal input
rlabel metal2 s 93030 0 93086 800 6 la_oen[2]
port 421 nsew signal input
rlabel metal2 s 161294 0 161350 800 6 la_oen[30]
port 422 nsew signal input
rlabel metal2 s 163778 0 163834 800 6 la_oen[31]
port 423 nsew signal input
rlabel metal2 s 166170 0 166226 800 6 la_oen[32]
port 424 nsew signal input
rlabel metal2 s 168654 0 168710 800 6 la_oen[33]
port 425 nsew signal input
rlabel metal2 s 171046 0 171102 800 6 la_oen[34]
port 426 nsew signal input
rlabel metal2 s 173530 0 173586 800 6 la_oen[35]
port 427 nsew signal input
rlabel metal2 s 175922 0 175978 800 6 la_oen[36]
port 428 nsew signal input
rlabel metal2 s 178406 0 178462 800 6 la_oen[37]
port 429 nsew signal input
rlabel metal2 s 180798 0 180854 800 6 la_oen[38]
port 430 nsew signal input
rlabel metal2 s 183282 0 183338 800 6 la_oen[39]
port 431 nsew signal input
rlabel metal2 s 95422 0 95478 800 6 la_oen[3]
port 432 nsew signal input
rlabel metal2 s 185674 0 185730 800 6 la_oen[40]
port 433 nsew signal input
rlabel metal2 s 188158 0 188214 800 6 la_oen[41]
port 434 nsew signal input
rlabel metal2 s 190550 0 190606 800 6 la_oen[42]
port 435 nsew signal input
rlabel metal2 s 193034 0 193090 800 6 la_oen[43]
port 436 nsew signal input
rlabel metal2 s 195426 0 195482 800 6 la_oen[44]
port 437 nsew signal input
rlabel metal2 s 197910 0 197966 800 6 la_oen[45]
port 438 nsew signal input
rlabel metal2 s 200394 0 200450 800 6 la_oen[46]
port 439 nsew signal input
rlabel metal2 s 202786 0 202842 800 6 la_oen[47]
port 440 nsew signal input
rlabel metal2 s 205270 0 205326 800 6 la_oen[48]
port 441 nsew signal input
rlabel metal2 s 207662 0 207718 800 6 la_oen[49]
port 442 nsew signal input
rlabel metal2 s 97906 0 97962 800 6 la_oen[4]
port 443 nsew signal input
rlabel metal2 s 210146 0 210202 800 6 la_oen[50]
port 444 nsew signal input
rlabel metal2 s 212538 0 212594 800 6 la_oen[51]
port 445 nsew signal input
rlabel metal2 s 215022 0 215078 800 6 la_oen[52]
port 446 nsew signal input
rlabel metal2 s 217414 0 217470 800 6 la_oen[53]
port 447 nsew signal input
rlabel metal2 s 219898 0 219954 800 6 la_oen[54]
port 448 nsew signal input
rlabel metal2 s 222290 0 222346 800 6 la_oen[55]
port 449 nsew signal input
rlabel metal2 s 224774 0 224830 800 6 la_oen[56]
port 450 nsew signal input
rlabel metal2 s 227166 0 227222 800 6 la_oen[57]
port 451 nsew signal input
rlabel metal2 s 229650 0 229706 800 6 la_oen[58]
port 452 nsew signal input
rlabel metal2 s 232042 0 232098 800 6 la_oen[59]
port 453 nsew signal input
rlabel metal2 s 100390 0 100446 800 6 la_oen[5]
port 454 nsew signal input
rlabel metal2 s 234526 0 234582 800 6 la_oen[60]
port 455 nsew signal input
rlabel metal2 s 236918 0 236974 800 6 la_oen[61]
port 456 nsew signal input
rlabel metal2 s 239402 0 239458 800 6 la_oen[62]
port 457 nsew signal input
rlabel metal2 s 241794 0 241850 800 6 la_oen[63]
port 458 nsew signal input
rlabel metal2 s 244278 0 244334 800 6 la_oen[64]
port 459 nsew signal input
rlabel metal2 s 246670 0 246726 800 6 la_oen[65]
port 460 nsew signal input
rlabel metal2 s 249154 0 249210 800 6 la_oen[66]
port 461 nsew signal input
rlabel metal2 s 251546 0 251602 800 6 la_oen[67]
port 462 nsew signal input
rlabel metal2 s 254030 0 254086 800 6 la_oen[68]
port 463 nsew signal input
rlabel metal2 s 256422 0 256478 800 6 la_oen[69]
port 464 nsew signal input
rlabel metal2 s 102782 0 102838 800 6 la_oen[6]
port 465 nsew signal input
rlabel metal2 s 258906 0 258962 800 6 la_oen[70]
port 466 nsew signal input
rlabel metal2 s 261298 0 261354 800 6 la_oen[71]
port 467 nsew signal input
rlabel metal2 s 263782 0 263838 800 6 la_oen[72]
port 468 nsew signal input
rlabel metal2 s 266174 0 266230 800 6 la_oen[73]
port 469 nsew signal input
rlabel metal2 s 268658 0 268714 800 6 la_oen[74]
port 470 nsew signal input
rlabel metal2 s 271050 0 271106 800 6 la_oen[75]
port 471 nsew signal input
rlabel metal2 s 273534 0 273590 800 6 la_oen[76]
port 472 nsew signal input
rlabel metal2 s 275926 0 275982 800 6 la_oen[77]
port 473 nsew signal input
rlabel metal2 s 278410 0 278466 800 6 la_oen[78]
port 474 nsew signal input
rlabel metal2 s 280802 0 280858 800 6 la_oen[79]
port 475 nsew signal input
rlabel metal2 s 105266 0 105322 800 6 la_oen[7]
port 476 nsew signal input
rlabel metal2 s 283286 0 283342 800 6 la_oen[80]
port 477 nsew signal input
rlabel metal2 s 285678 0 285734 800 6 la_oen[81]
port 478 nsew signal input
rlabel metal2 s 288162 0 288218 800 6 la_oen[82]
port 479 nsew signal input
rlabel metal2 s 290554 0 290610 800 6 la_oen[83]
port 480 nsew signal input
rlabel metal2 s 293038 0 293094 800 6 la_oen[84]
port 481 nsew signal input
rlabel metal2 s 295430 0 295486 800 6 la_oen[85]
port 482 nsew signal input
rlabel metal2 s 297914 0 297970 800 6 la_oen[86]
port 483 nsew signal input
rlabel metal2 s 300398 0 300454 800 6 la_oen[87]
port 484 nsew signal input
rlabel metal2 s 302790 0 302846 800 6 la_oen[88]
port 485 nsew signal input
rlabel metal2 s 305274 0 305330 800 6 la_oen[89]
port 486 nsew signal input
rlabel metal2 s 107658 0 107714 800 6 la_oen[8]
port 487 nsew signal input
rlabel metal2 s 307666 0 307722 800 6 la_oen[90]
port 488 nsew signal input
rlabel metal2 s 310150 0 310206 800 6 la_oen[91]
port 489 nsew signal input
rlabel metal2 s 312542 0 312598 800 6 la_oen[92]
port 490 nsew signal input
rlabel metal2 s 315026 0 315082 800 6 la_oen[93]
port 491 nsew signal input
rlabel metal2 s 317418 0 317474 800 6 la_oen[94]
port 492 nsew signal input
rlabel metal2 s 319902 0 319958 800 6 la_oen[95]
port 493 nsew signal input
rlabel metal2 s 322294 0 322350 800 6 la_oen[96]
port 494 nsew signal input
rlabel metal2 s 324778 0 324834 800 6 la_oen[97]
port 495 nsew signal input
rlabel metal2 s 327170 0 327226 800 6 la_oen[98]
port 496 nsew signal input
rlabel metal2 s 329654 0 329710 800 6 la_oen[99]
port 497 nsew signal input
rlabel metal2 s 110142 0 110198 800 6 la_oen[9]
port 498 nsew signal input
rlabel metal3 s 0 124992 800 125112 6 vccd1
port 499 nsew signal bidirectional
rlabel metal2 s 391386 499200 391442 500000 6 vccd2
port 500 nsew signal bidirectional
rlabel metal2 s 394790 499200 394846 500000 6 vdda1
port 501 nsew signal bidirectional
rlabel metal2 s 398746 0 398802 800 6 vdda2
port 502 nsew signal bidirectional
rlabel metal3 s 0 374960 800 375080 6 vssa1
port 503 nsew signal bidirectional
rlabel metal3 s 399200 249976 400000 250096 6 vssa2
port 504 nsew signal bidirectional
rlabel metal2 s 399574 0 399630 800 6 vssd1
port 505 nsew signal bidirectional
rlabel metal2 s 398194 499200 398250 500000 6 vssd2
port 506 nsew signal bidirectional
rlabel metal2 s 386 0 442 800 6 wb_clk_i
port 507 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 wb_rst_i
port 508 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 wbs_ack_o
port 509 nsew signal output
rlabel metal2 s 5262 0 5318 800 6 wbs_adr_i[0]
port 510 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 wbs_adr_i[10]
port 511 nsew signal input
rlabel metal2 s 35346 0 35402 800 6 wbs_adr_i[11]
port 512 nsew signal input
rlabel metal2 s 37738 0 37794 800 6 wbs_adr_i[12]
port 513 nsew signal input
rlabel metal2 s 40222 0 40278 800 6 wbs_adr_i[13]
port 514 nsew signal input
rlabel metal2 s 42614 0 42670 800 6 wbs_adr_i[14]
port 515 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 wbs_adr_i[15]
port 516 nsew signal input
rlabel metal2 s 47490 0 47546 800 6 wbs_adr_i[16]
port 517 nsew signal input
rlabel metal2 s 49974 0 50030 800 6 wbs_adr_i[17]
port 518 nsew signal input
rlabel metal2 s 52366 0 52422 800 6 wbs_adr_i[18]
port 519 nsew signal input
rlabel metal2 s 54850 0 54906 800 6 wbs_adr_i[19]
port 520 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 wbs_adr_i[1]
port 521 nsew signal input
rlabel metal2 s 57242 0 57298 800 6 wbs_adr_i[20]
port 522 nsew signal input
rlabel metal2 s 59726 0 59782 800 6 wbs_adr_i[21]
port 523 nsew signal input
rlabel metal2 s 62118 0 62174 800 6 wbs_adr_i[22]
port 524 nsew signal input
rlabel metal2 s 64602 0 64658 800 6 wbs_adr_i[23]
port 525 nsew signal input
rlabel metal2 s 66994 0 67050 800 6 wbs_adr_i[24]
port 526 nsew signal input
rlabel metal2 s 69478 0 69534 800 6 wbs_adr_i[25]
port 527 nsew signal input
rlabel metal2 s 71870 0 71926 800 6 wbs_adr_i[26]
port 528 nsew signal input
rlabel metal2 s 74354 0 74410 800 6 wbs_adr_i[27]
port 529 nsew signal input
rlabel metal2 s 76746 0 76802 800 6 wbs_adr_i[28]
port 530 nsew signal input
rlabel metal2 s 79230 0 79286 800 6 wbs_adr_i[29]
port 531 nsew signal input
rlabel metal2 s 11702 0 11758 800 6 wbs_adr_i[2]
port 532 nsew signal input
rlabel metal2 s 81622 0 81678 800 6 wbs_adr_i[30]
port 533 nsew signal input
rlabel metal2 s 84106 0 84162 800 6 wbs_adr_i[31]
port 534 nsew signal input
rlabel metal2 s 15014 0 15070 800 6 wbs_adr_i[3]
port 535 nsew signal input
rlabel metal2 s 18234 0 18290 800 6 wbs_adr_i[4]
port 536 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 wbs_adr_i[5]
port 537 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 wbs_adr_i[6]
port 538 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 wbs_adr_i[7]
port 539 nsew signal input
rlabel metal2 s 27986 0 28042 800 6 wbs_adr_i[8]
port 540 nsew signal input
rlabel metal2 s 30378 0 30434 800 6 wbs_adr_i[9]
port 541 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 wbs_cyc_i
port 542 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 wbs_dat_i[0]
port 543 nsew signal input
rlabel metal2 s 33690 0 33746 800 6 wbs_dat_i[10]
port 544 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 wbs_dat_i[11]
port 545 nsew signal input
rlabel metal2 s 38566 0 38622 800 6 wbs_dat_i[12]
port 546 nsew signal input
rlabel metal2 s 40958 0 41014 800 6 wbs_dat_i[13]
port 547 nsew signal input
rlabel metal2 s 43442 0 43498 800 6 wbs_dat_i[14]
port 548 nsew signal input
rlabel metal2 s 45834 0 45890 800 6 wbs_dat_i[15]
port 549 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 wbs_dat_i[16]
port 550 nsew signal input
rlabel metal2 s 50710 0 50766 800 6 wbs_dat_i[17]
port 551 nsew signal input
rlabel metal2 s 53194 0 53250 800 6 wbs_dat_i[18]
port 552 nsew signal input
rlabel metal2 s 55586 0 55642 800 6 wbs_dat_i[19]
port 553 nsew signal input
rlabel metal2 s 9310 0 9366 800 6 wbs_dat_i[1]
port 554 nsew signal input
rlabel metal2 s 58070 0 58126 800 6 wbs_dat_i[20]
port 555 nsew signal input
rlabel metal2 s 60462 0 60518 800 6 wbs_dat_i[21]
port 556 nsew signal input
rlabel metal2 s 62946 0 63002 800 6 wbs_dat_i[22]
port 557 nsew signal input
rlabel metal2 s 65338 0 65394 800 6 wbs_dat_i[23]
port 558 nsew signal input
rlabel metal2 s 67822 0 67878 800 6 wbs_dat_i[24]
port 559 nsew signal input
rlabel metal2 s 70306 0 70362 800 6 wbs_dat_i[25]
port 560 nsew signal input
rlabel metal2 s 72698 0 72754 800 6 wbs_dat_i[26]
port 561 nsew signal input
rlabel metal2 s 75182 0 75238 800 6 wbs_dat_i[27]
port 562 nsew signal input
rlabel metal2 s 77574 0 77630 800 6 wbs_dat_i[28]
port 563 nsew signal input
rlabel metal2 s 80058 0 80114 800 6 wbs_dat_i[29]
port 564 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 wbs_dat_i[2]
port 565 nsew signal input
rlabel metal2 s 82450 0 82506 800 6 wbs_dat_i[30]
port 566 nsew signal input
rlabel metal2 s 84934 0 84990 800 6 wbs_dat_i[31]
port 567 nsew signal input
rlabel metal2 s 15750 0 15806 800 6 wbs_dat_i[3]
port 568 nsew signal input
rlabel metal2 s 19062 0 19118 800 6 wbs_dat_i[4]
port 569 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 wbs_dat_i[5]
port 570 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 wbs_dat_i[6]
port 571 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 wbs_dat_i[7]
port 572 nsew signal input
rlabel metal2 s 28814 0 28870 800 6 wbs_dat_i[8]
port 573 nsew signal input
rlabel metal2 s 31206 0 31262 800 6 wbs_dat_i[9]
port 574 nsew signal input
rlabel metal2 s 6826 0 6882 800 6 wbs_dat_o[0]
port 575 nsew signal output
rlabel metal2 s 34518 0 34574 800 6 wbs_dat_o[10]
port 576 nsew signal output
rlabel metal2 s 36910 0 36966 800 6 wbs_dat_o[11]
port 577 nsew signal output
rlabel metal2 s 39394 0 39450 800 6 wbs_dat_o[12]
port 578 nsew signal output
rlabel metal2 s 41786 0 41842 800 6 wbs_dat_o[13]
port 579 nsew signal output
rlabel metal2 s 44270 0 44326 800 6 wbs_dat_o[14]
port 580 nsew signal output
rlabel metal2 s 46662 0 46718 800 6 wbs_dat_o[15]
port 581 nsew signal output
rlabel metal2 s 49146 0 49202 800 6 wbs_dat_o[16]
port 582 nsew signal output
rlabel metal2 s 51538 0 51594 800 6 wbs_dat_o[17]
port 583 nsew signal output
rlabel metal2 s 54022 0 54078 800 6 wbs_dat_o[18]
port 584 nsew signal output
rlabel metal2 s 56414 0 56470 800 6 wbs_dat_o[19]
port 585 nsew signal output
rlabel metal2 s 10138 0 10194 800 6 wbs_dat_o[1]
port 586 nsew signal output
rlabel metal2 s 58898 0 58954 800 6 wbs_dat_o[20]
port 587 nsew signal output
rlabel metal2 s 61290 0 61346 800 6 wbs_dat_o[21]
port 588 nsew signal output
rlabel metal2 s 63774 0 63830 800 6 wbs_dat_o[22]
port 589 nsew signal output
rlabel metal2 s 66166 0 66222 800 6 wbs_dat_o[23]
port 590 nsew signal output
rlabel metal2 s 68650 0 68706 800 6 wbs_dat_o[24]
port 591 nsew signal output
rlabel metal2 s 71042 0 71098 800 6 wbs_dat_o[25]
port 592 nsew signal output
rlabel metal2 s 73526 0 73582 800 6 wbs_dat_o[26]
port 593 nsew signal output
rlabel metal2 s 75918 0 75974 800 6 wbs_dat_o[27]
port 594 nsew signal output
rlabel metal2 s 78402 0 78458 800 6 wbs_dat_o[28]
port 595 nsew signal output
rlabel metal2 s 80794 0 80850 800 6 wbs_dat_o[29]
port 596 nsew signal output
rlabel metal2 s 13358 0 13414 800 6 wbs_dat_o[2]
port 597 nsew signal output
rlabel metal2 s 83278 0 83334 800 6 wbs_dat_o[30]
port 598 nsew signal output
rlabel metal2 s 85670 0 85726 800 6 wbs_dat_o[31]
port 599 nsew signal output
rlabel metal2 s 16578 0 16634 800 6 wbs_dat_o[3]
port 600 nsew signal output
rlabel metal2 s 19890 0 19946 800 6 wbs_dat_o[4]
port 601 nsew signal output
rlabel metal2 s 22282 0 22338 800 6 wbs_dat_o[5]
port 602 nsew signal output
rlabel metal2 s 24766 0 24822 800 6 wbs_dat_o[6]
port 603 nsew signal output
rlabel metal2 s 27158 0 27214 800 6 wbs_dat_o[7]
port 604 nsew signal output
rlabel metal2 s 29642 0 29698 800 6 wbs_dat_o[8]
port 605 nsew signal output
rlabel metal2 s 32034 0 32090 800 6 wbs_dat_o[9]
port 606 nsew signal output
rlabel metal2 s 7654 0 7710 800 6 wbs_sel_i[0]
port 607 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 wbs_sel_i[1]
port 608 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 wbs_sel_i[2]
port 609 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 wbs_sel_i[3]
port 610 nsew signal input
rlabel metal2 s 3606 0 3662 800 6 wbs_stb_i
port 611 nsew signal input
rlabel metal2 s 4434 0 4490 800 6 wbs_we_i
port 612 nsew signal input
rlabel metal4 s 372848 2128 373168 497808 6 VPWR
port 613 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 497808 6 VPWR
port 614 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 497808 6 VPWR
port 615 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 497808 6 VPWR
port 616 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 497808 6 VPWR
port 617 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 497808 6 VPWR
port 618 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 497808 6 VPWR
port 619 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 497808 6 VPWR
port 620 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 497808 6 VPWR
port 621 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 497808 6 VPWR
port 622 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 497808 6 VPWR
port 623 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 497808 6 VPWR
port 624 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 497808 6 VPWR
port 625 nsew power bidirectional
rlabel metal4 s 388208 2128 388528 497808 6 VGND
port 626 nsew ground bidirectional
rlabel metal4 s 357488 2128 357808 497808 6 VGND
port 627 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 497808 6 VGND
port 628 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 497808 6 VGND
port 629 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 497808 6 VGND
port 630 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 497808 6 VGND
port 631 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 497808 6 VGND
port 632 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 497808 6 VGND
port 633 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 497808 6 VGND
port 634 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 497808 6 VGND
port 635 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 497808 6 VGND
port 636 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 497808 6 VGND
port 637 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 497808 6 VGND
port 638 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 400000 500000
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj_aes/runs/user_proj_aes/results/magic/user_proj_aes.gds
string GDS_END 94485806
string GDS_START 270814
<< end >>

