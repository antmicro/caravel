magic
tech sky130A
magscale 1 2
timestamp 1607420573
<< locali >>
rect 269405 699703 269439 700009
rect 291393 698207 291427 700417
rect 267565 685967 267599 688721
rect 269221 685967 269255 695453
rect 287161 688347 287195 695453
rect 289921 688619 289955 695453
rect 291393 688619 291427 695453
rect 252385 676243 252419 685797
rect 267565 682975 267599 684437
rect 269221 676243 269255 684437
rect 252385 656931 252419 666485
rect 267381 665295 267415 674781
rect 287161 666587 287195 676141
rect 299857 666587 299891 684437
rect 494069 666587 494103 676141
rect 559297 666587 559331 684437
rect 267565 659583 267599 665125
rect 252385 637619 252419 647173
rect 267473 645915 267507 650165
rect 269405 649927 269439 663697
rect 276121 656931 276155 666485
rect 289829 656931 289863 666485
rect 289829 637619 289863 647173
rect 267473 626671 267507 630853
rect 291301 627963 291335 637517
rect 289921 618307 289955 627861
rect 291301 608651 291335 618205
rect 287161 598995 287195 608549
rect 267289 589407 267323 592093
rect 269129 589339 269163 598893
rect 276213 591991 276247 598893
rect 291301 597567 291335 607121
rect 299673 601715 299707 608549
rect 559113 601715 559147 608549
rect 299765 589339 299799 598893
rect 559297 589339 559331 598893
rect 269221 582403 269255 587809
rect 276213 582267 276247 589237
rect 291393 569959 291427 579581
rect 494161 563091 494195 569857
rect 559021 550647 559055 560201
rect 287161 531335 287195 534089
rect 276247 521645 276489 521679
rect 287103 521645 287345 521679
rect 17141 519095 17175 519605
rect 17233 519231 17267 519537
rect 17325 518959 17359 519673
rect 22753 519231 22787 519537
rect 26801 518959 26835 519673
rect 26893 519095 26927 519605
rect 36461 519095 36495 519605
rect 36553 519231 36587 519537
rect 36645 518959 36679 519673
rect 42073 519231 42107 519537
rect 46121 518959 46155 519673
rect 46213 519095 46247 519605
rect 55781 519095 55815 519605
rect 55873 519231 55907 519537
rect 55965 518959 55999 519673
rect 61393 519231 61427 519537
rect 65441 518959 65475 519673
rect 65533 519095 65567 519605
rect 75101 519095 75135 519605
rect 75193 519231 75227 519537
rect 75285 518959 75319 519673
rect 80713 519231 80747 519537
rect 84761 518959 84795 519673
rect 84853 519095 84887 519605
rect 94421 519095 94455 519605
rect 94513 519231 94547 519537
rect 94605 518959 94639 519673
rect 100033 519231 100067 519537
rect 104081 518959 104115 519673
rect 104173 519095 104207 519605
rect 113741 519095 113775 519605
rect 113833 519231 113867 519537
rect 113925 518959 113959 519673
rect 119353 519231 119387 519537
rect 123401 518959 123435 519673
rect 123493 519095 123527 519605
rect 133061 519095 133095 519605
rect 133153 519231 133187 519537
rect 133245 518959 133279 519673
rect 138673 519231 138707 519537
rect 142721 518959 142755 519673
rect 142813 519095 142847 519605
rect 152381 519095 152415 519605
rect 152473 519231 152507 519537
rect 152565 518959 152599 519673
rect 157993 519231 158027 519537
rect 162041 518959 162075 519673
rect 162133 519095 162167 519605
rect 171701 519095 171735 519673
rect 171793 519231 171827 519605
rect 171885 518959 171919 519741
rect 179429 518211 179463 519537
rect 181361 519095 181395 519673
rect 181453 519231 181487 519605
rect 181545 518959 181579 519741
rect 188353 518959 188387 519673
rect 190009 519231 190043 519537
rect 191113 519095 191147 519605
rect 195989 519231 196023 519537
rect 200681 518959 200715 519673
rect 200773 519095 200807 519605
rect 209789 519231 209823 519605
rect 209881 519095 209915 519673
rect 209823 519061 209915 519095
rect 209973 518959 210007 519741
rect 209823 518925 210007 518959
rect 219173 518959 219207 519741
rect 219265 519095 219299 519673
rect 219357 519231 219391 519605
rect 305377 519231 305411 519605
rect 316877 519231 316911 519605
rect 325709 519231 325743 519333
rect 306883 519129 307033 519163
rect 316785 519095 316819 519197
rect 325801 519095 325835 519401
rect 219265 519061 219357 519095
rect 306849 519061 307125 519095
rect 325743 519061 325835 519095
rect 306849 518959 306883 519061
rect 219173 518925 219357 518959
rect 316693 518959 316727 519061
rect 325893 518959 325927 519469
rect 325743 518925 325927 518959
rect 335185 518959 335219 519469
rect 335277 519095 335311 519401
rect 345121 518959 345155 519129
rect 349997 519095 350031 519265
rect 335185 518925 335277 518959
rect 345063 518925 345155 518959
rect 351837 518279 351871 519265
rect 355149 519027 355183 519265
rect 275879 217957 275937 217991
rect 329297 217923 329331 218025
rect 281549 217719 281583 217821
rect 170873 217515 170907 217685
rect 168297 217447 168331 217481
rect 170781 217447 170815 217481
rect 170965 217447 170999 217685
rect 167009 217413 167193 217447
rect 168297 217413 168481 217447
rect 170781 217413 170999 217447
rect 167009 217379 167043 217413
rect 167101 217311 167135 217345
rect 167101 217277 167285 217311
rect 180165 212551 180199 217685
rect 181453 216699 181487 217277
rect 212365 212551 212399 217685
rect 281733 217447 281767 217821
rect 281825 217175 281859 217413
rect 282009 216903 282043 217073
rect 282929 216767 282963 217345
rect 283113 216835 283147 217889
rect 292623 217685 292715 217719
rect 292681 217447 292715 217685
rect 289829 216699 289863 216869
rect 291209 216767 291243 217277
rect 295349 217039 295383 217617
rect 321569 217515 321603 217889
rect 323593 217515 323627 217889
rect 332333 217855 332367 218025
rect 320005 217243 320039 217481
rect 302157 216835 302191 217073
rect 319913 217039 319947 217209
rect 216965 212551 216999 215305
rect 291945 215203 291979 216801
rect 307217 216835 307251 217005
rect 308447 216869 308689 216903
rect 299397 216699 299431 216801
rect 311909 216767 311943 216937
rect 331137 216699 331171 217549
rect 332425 217379 332459 217821
rect 335369 217447 335403 217821
rect 337485 217821 337853 217855
rect 337485 217719 337519 217821
rect 336657 217447 336691 217685
rect 339417 217379 339451 218161
rect 340613 217855 340647 218025
rect 340739 217957 340831 217991
rect 339509 217447 339543 217685
rect 340521 217413 340705 217447
rect 340521 217311 340555 217413
rect 340797 217379 340831 217957
rect 350549 217787 350583 217889
rect 369777 216767 369811 217685
rect 211905 202895 211939 212449
rect 217057 201535 217091 211089
rect 219817 202895 219851 205649
rect 258273 202895 258307 207689
rect 262597 205615 262631 211089
rect 315865 202895 315899 205649
rect 328101 205615 328135 211089
rect 329389 201467 329423 209729
rect 343281 205615 343315 211089
rect 344569 205615 344603 211089
rect 171517 193239 171551 195993
rect 192125 193171 192159 201433
rect 179981 179435 180015 188989
rect 182189 182223 182223 186337
rect 262505 186303 262539 191777
rect 277225 183583 277259 200073
rect 282837 193171 282871 201433
rect 315773 191879 315807 196061
rect 315681 182223 315715 191709
rect 328193 186303 328227 193069
rect 362509 191879 362543 201433
rect 176945 173179 176979 179333
rect 181085 169779 181119 179333
rect 182189 176579 182223 181985
rect 192217 176103 192251 182121
rect 217333 171139 217367 180761
rect 224049 172567 224083 182121
rect 262597 172567 262631 182053
rect 177129 158763 177163 168317
rect 182189 161483 182223 171037
rect 181085 151827 181119 161381
rect 182189 156723 182223 161313
rect 192217 153255 192251 156757
rect 177129 139519 177163 149005
rect 178141 139519 178175 149005
rect 203165 144891 203199 161381
rect 211905 154615 211939 171037
rect 212457 154615 212491 164169
rect 225429 162707 225463 172465
rect 229385 164203 229419 172465
rect 275845 171139 275879 180761
rect 277133 172567 277167 182121
rect 217149 151827 217183 161381
rect 225613 150331 225647 158661
rect 177129 129795 177163 139349
rect 178141 129795 178175 139349
rect 179981 131223 180015 140709
rect 181085 132583 181119 142069
rect 171425 115991 171459 125545
rect 173081 115991 173115 125545
rect 181085 122859 181119 132413
rect 182189 124219 182223 142069
rect 194885 131155 194919 140709
rect 211905 135303 211939 144857
rect 201785 124219 201819 133841
rect 203073 132515 203107 133977
rect 212273 131155 212307 140709
rect 228189 139451 228223 157301
rect 229293 153255 229327 162809
rect 236377 160191 236411 171037
rect 285229 166923 285263 182121
rect 329573 181611 329607 191777
rect 354229 183515 354263 191777
rect 354321 176579 354355 182121
rect 355609 176647 355643 182121
rect 362417 171207 362451 182121
rect 318441 164271 318475 169133
rect 258273 157335 258307 164169
rect 344569 162911 344603 167501
rect 355609 164271 355643 167025
rect 261125 153255 261159 162809
rect 286701 153255 286735 162809
rect 317153 157335 317187 162809
rect 318441 157335 318475 162809
rect 230949 144891 230983 153153
rect 291945 145027 291979 154513
rect 341993 153255 342027 162809
rect 299213 144959 299247 147781
rect 300501 144959 300535 147781
rect 181177 121431 181211 122689
rect 178325 110483 178359 120037
rect 180993 111911 181027 121397
rect 182189 118031 182223 122757
rect 171425 96679 171459 106233
rect 173081 96679 173115 106233
rect 181085 102255 181119 111741
rect 184029 108851 184063 115889
rect 192309 110415 192343 122757
rect 200313 115855 200347 124117
rect 203073 114563 203107 124117
rect 211905 115991 211939 125545
rect 194885 104907 194919 114461
rect 201877 104907 201911 114461
rect 212273 113135 212307 121397
rect 229201 118031 229235 122757
rect 231041 114563 231075 124117
rect 232237 113203 232271 122757
rect 236285 120683 236319 142069
rect 258273 137955 258307 144857
rect 317245 143599 317279 147645
rect 328285 144959 328319 147645
rect 261125 133943 261159 143497
rect 275845 133943 275879 143497
rect 285321 137955 285355 143497
rect 286609 137955 286643 143497
rect 289369 137955 289403 143497
rect 235273 115991 235307 118677
rect 258273 118643 258307 125545
rect 277225 124219 277259 133841
rect 315865 132515 315899 142069
rect 318441 134011 318475 143497
rect 329573 135303 329607 144857
rect 341993 140811 342027 142137
rect 343281 140811 343315 158661
rect 345673 151827 345707 161381
rect 354321 157335 354355 162809
rect 355517 153255 355551 162809
rect 362417 161483 362451 171037
rect 361221 150535 361255 160021
rect 362417 144891 362451 156621
rect 299213 124219 299247 128469
rect 300501 124219 300535 128469
rect 318441 125579 318475 133841
rect 341717 129795 341751 139349
rect 361405 132515 361439 142069
rect 328285 124219 328319 128333
rect 261125 114563 261159 124117
rect 177037 92531 177071 102085
rect 178049 91103 178083 95081
rect 179981 92531 180015 102085
rect 182189 99331 182223 104737
rect 211905 100079 211939 106233
rect 217057 102187 217091 111673
rect 219817 103615 219851 113101
rect 273085 106335 273119 115889
rect 277225 114563 277259 118745
rect 282745 114563 282779 115957
rect 291945 114563 291979 124117
rect 315865 114563 315899 118745
rect 318533 114563 318567 124117
rect 329573 115991 329607 125545
rect 343281 121499 343315 131053
rect 345581 122859 345615 132413
rect 354413 124219 354447 128333
rect 355701 124219 355735 128333
rect 362325 115923 362359 121397
rect 171425 77299 171459 86921
rect 173081 77299 173115 86921
rect 182189 84235 182223 93789
rect 194885 85595 194919 95149
rect 171425 57987 171459 67541
rect 173081 57987 173115 67541
rect 178141 63563 178175 81345
rect 179981 73219 180015 82773
rect 181269 64923 181303 74477
rect 184029 66283 184063 75837
rect 191113 74579 191147 84133
rect 192309 66283 192343 84133
rect 201877 77299 201911 86921
rect 217241 84235 217275 95353
rect 219725 93891 219759 103445
rect 224049 95251 224083 99501
rect 225337 95251 225371 99637
rect 235273 96679 235307 99365
rect 236285 96679 236319 106233
rect 258273 99331 258307 106233
rect 277225 104975 277259 114393
rect 354229 113203 354263 114597
rect 261125 95251 261159 104805
rect 275845 95251 275879 104805
rect 277133 95251 277167 104805
rect 282745 95251 282779 104805
rect 283941 95251 283975 104805
rect 300501 103547 300535 109157
rect 315865 104907 315899 109089
rect 299213 102255 299247 103513
rect 315773 87023 315807 96917
rect 317245 96679 317279 109701
rect 318349 104907 318383 109361
rect 329573 96679 329607 106233
rect 341901 103547 341935 113033
rect 344477 93891 344511 103445
rect 354413 96679 354447 109701
rect 355609 103547 355643 113101
rect 194885 66283 194919 77197
rect 203073 71111 203107 80665
rect 235273 77299 235307 80053
rect 232237 75939 232271 77265
rect 236285 75939 236319 86921
rect 258273 77299 258307 86921
rect 260941 75939 260975 85493
rect 262321 77299 262355 86921
rect 282745 75939 282779 77333
rect 283941 75939 283975 85493
rect 289277 75939 289311 85493
rect 355701 84235 355735 93789
rect 361221 85527 361255 93789
rect 318257 75939 318291 77537
rect 217149 66283 217183 75769
rect 341993 73287 342027 74613
rect 343281 74579 343315 84133
rect 219725 66283 219759 70465
rect 344569 67643 344603 79305
rect 345581 74579 345615 84133
rect 361313 79339 361347 84133
rect 355977 67371 356011 75837
rect 362325 67643 362359 84133
rect 177037 57919 177071 63461
rect 179981 53839 180015 63461
rect 181085 53839 181119 58633
rect 171425 38675 171459 48229
rect 183937 45611 183971 55165
rect 200405 48331 200439 61421
rect 201877 53975 201911 61421
rect 203073 55267 203107 64821
rect 230765 56627 230799 65909
rect 179981 35955 180015 45509
rect 171333 19363 171367 28917
rect 181085 26299 181119 44081
rect 182189 27659 182223 41429
rect 189549 27659 189583 40681
rect 201877 27659 201911 45509
rect 212457 37315 212491 48229
rect 228189 46903 228223 55165
rect 262505 48331 262539 57885
rect 275753 53839 275787 63461
rect 277133 48331 277167 63461
rect 283941 56695 283975 66181
rect 285321 56627 285355 66181
rect 286609 56627 286643 66181
rect 289369 56627 289403 66181
rect 329573 56627 329607 66181
rect 283941 46971 283975 56525
rect 318349 46971 318383 56525
rect 344477 55267 344511 64821
rect 219817 35955 219851 42449
rect 232053 37315 232087 46869
rect 258273 31739 258307 38573
rect 273085 37179 273119 45509
rect 275845 33235 275879 38573
rect 317153 37315 317187 46869
rect 329389 37315 329423 42109
rect 344569 41123 344603 51765
rect 345673 46971 345707 59993
rect 354321 48399 354355 57885
rect 355609 48331 355643 64821
rect 362325 48331 362359 57885
rect 354321 41123 354355 48229
rect 200405 26299 200439 27625
rect 178141 16643 178175 26197
rect 179981 16643 180015 26197
rect 182373 17799 182407 17969
rect 192125 9707 192159 19261
rect 194885 16643 194919 26197
rect 212273 19295 212307 27557
rect 236377 19363 236411 28917
rect 212273 9707 212307 12529
rect 214297 9707 214331 19261
rect 261125 18003 261159 27557
rect 268761 18003 268795 27557
rect 275937 18003 275971 27557
rect 228131 17901 228281 17935
rect 277133 9707 277167 27557
rect 317153 19363 317187 28849
rect 328101 27659 328135 31773
rect 329481 19363 329515 28917
rect 343373 28475 343407 37281
rect 344661 29019 344695 38573
rect 361313 29019 361347 31773
rect 362417 29019 362451 31841
rect 283941 8347 283975 9741
rect 289277 8075 289311 13073
rect 291853 9707 291887 19261
rect 328193 9707 328227 19261
rect 341901 13787 341935 18377
rect 343281 13719 343315 27557
rect 344569 13651 344603 27557
rect 345673 18003 345707 27557
rect 329481 9707 329515 12461
rect 352941 11747 352975 19261
rect 354321 18003 354355 27557
rect 355517 18003 355551 27557
rect 361221 18003 361255 27557
rect 362509 9707 362543 19261
rect 287621 4165 288023 4199
rect 234755 3961 234847 3995
rect 225245 3791 225279 3893
rect 225153 3519 225187 3757
rect 225061 3383 225095 3485
rect 226349 3383 226383 3893
rect 234813 3723 234847 3961
rect 238769 3859 238803 4029
rect 273085 3859 273119 4029
rect 286091 4029 286241 4063
rect 273177 3655 273211 3825
rect 274189 3655 274223 3757
rect 67925 3043 67959 3281
rect 69581 3281 69799 3315
rect 69581 3043 69615 3281
rect 69765 3247 69799 3281
rect 64889 2839 64923 2941
rect 69673 2839 69707 3213
rect 74549 3043 74583 3281
rect 77769 3111 77803 3281
rect 78965 3111 78999 3281
rect 77769 3077 78045 3111
rect 69765 2771 69799 3009
rect 79425 2975 79459 3145
rect 79333 2839 79367 2941
rect 79517 2771 79551 3145
rect 81357 2771 81391 3281
rect 82553 3281 82829 3315
rect 82553 3179 82587 3281
rect 224969 3247 225003 3349
rect 228741 3247 228775 3417
rect 274373 3315 274407 3825
rect 224969 3213 225061 3247
rect 275753 3179 275787 3485
rect 277961 3111 277995 3961
rect 278145 3927 278179 4029
rect 287621 3995 287655 4165
rect 287989 4131 288023 4165
rect 287563 3961 287655 3995
rect 287713 3723 287747 3961
rect 287897 3723 287931 4097
rect 278053 3519 278087 3689
rect 297281 3247 297315 3417
rect 301605 3247 301639 3417
rect 277961 3077 278329 3111
rect 84117 2771 84151 3009
rect 86049 2975 86083 3077
rect 280353 3043 280387 3213
rect 95525 2839 95559 3009
rect 277869 2975 277903 3009
rect 278053 3009 278237 3043
rect 297281 3213 297465 3247
rect 278053 2975 278087 3009
rect 277869 2941 278087 2975
rect 297189 2975 297223 3213
rect 306297 2975 306331 3213
rect 313565 3111 313599 3281
rect 308321 2975 308355 3077
rect 364993 3043 365027 3417
rect 121503 2873 121653 2907
<< viali >>
rect 291393 700417 291427 700451
rect 269405 700009 269439 700043
rect 269405 699669 269439 699703
rect 291393 698173 291427 698207
rect 269221 695453 269255 695487
rect 267565 688721 267599 688755
rect 267565 685933 267599 685967
rect 287161 695453 287195 695487
rect 289921 695453 289955 695487
rect 289921 688585 289955 688619
rect 291393 695453 291427 695487
rect 291393 688585 291427 688619
rect 287161 688313 287195 688347
rect 269221 685933 269255 685967
rect 252385 685797 252419 685831
rect 267565 684437 267599 684471
rect 267565 682941 267599 682975
rect 269221 684437 269255 684471
rect 252385 676209 252419 676243
rect 269221 676209 269255 676243
rect 299857 684437 299891 684471
rect 287161 676141 287195 676175
rect 267381 674781 267415 674815
rect 252385 666485 252419 666519
rect 287161 666553 287195 666587
rect 559297 684437 559331 684471
rect 299857 666553 299891 666587
rect 494069 676141 494103 676175
rect 494069 666553 494103 666587
rect 559297 666553 559331 666587
rect 267381 665261 267415 665295
rect 276121 666485 276155 666519
rect 267565 665125 267599 665159
rect 267565 659549 267599 659583
rect 269405 663697 269439 663731
rect 252385 656897 252419 656931
rect 267473 650165 267507 650199
rect 252385 647173 252419 647207
rect 276121 656897 276155 656931
rect 289829 666485 289863 666519
rect 289829 656897 289863 656931
rect 269405 649893 269439 649927
rect 267473 645881 267507 645915
rect 289829 647173 289863 647207
rect 252385 637585 252419 637619
rect 289829 637585 289863 637619
rect 291301 637517 291335 637551
rect 267473 630853 267507 630887
rect 291301 627929 291335 627963
rect 267473 626637 267507 626671
rect 289921 627861 289955 627895
rect 289921 618273 289955 618307
rect 291301 618205 291335 618239
rect 291301 608617 291335 608651
rect 287161 608549 287195 608583
rect 299673 608549 299707 608583
rect 287161 598961 287195 598995
rect 291301 607121 291335 607155
rect 269129 598893 269163 598927
rect 267289 592093 267323 592127
rect 267289 589373 267323 589407
rect 276213 598893 276247 598927
rect 299673 601681 299707 601715
rect 559113 608549 559147 608583
rect 559113 601681 559147 601715
rect 291301 597533 291335 597567
rect 299765 598893 299799 598927
rect 276213 591957 276247 591991
rect 269129 589305 269163 589339
rect 299765 589305 299799 589339
rect 559297 598893 559331 598927
rect 559297 589305 559331 589339
rect 276213 589237 276247 589271
rect 269221 587809 269255 587843
rect 269221 582369 269255 582403
rect 276213 582233 276247 582267
rect 291393 579581 291427 579615
rect 291393 569925 291427 569959
rect 494161 569857 494195 569891
rect 494161 563057 494195 563091
rect 559021 560201 559055 560235
rect 559021 550613 559055 550647
rect 287161 534089 287195 534123
rect 287161 531301 287195 531335
rect 276213 521645 276247 521679
rect 276489 521645 276523 521679
rect 287069 521645 287103 521679
rect 287345 521645 287379 521679
rect 171885 519741 171919 519775
rect 17325 519673 17359 519707
rect 17141 519605 17175 519639
rect 17233 519537 17267 519571
rect 17233 519197 17267 519231
rect 17141 519061 17175 519095
rect 26801 519673 26835 519707
rect 22753 519537 22787 519571
rect 22753 519197 22787 519231
rect 17325 518925 17359 518959
rect 36645 519673 36679 519707
rect 26893 519605 26927 519639
rect 26893 519061 26927 519095
rect 36461 519605 36495 519639
rect 36553 519537 36587 519571
rect 36553 519197 36587 519231
rect 36461 519061 36495 519095
rect 26801 518925 26835 518959
rect 46121 519673 46155 519707
rect 42073 519537 42107 519571
rect 42073 519197 42107 519231
rect 36645 518925 36679 518959
rect 55965 519673 55999 519707
rect 46213 519605 46247 519639
rect 46213 519061 46247 519095
rect 55781 519605 55815 519639
rect 55873 519537 55907 519571
rect 55873 519197 55907 519231
rect 55781 519061 55815 519095
rect 46121 518925 46155 518959
rect 65441 519673 65475 519707
rect 61393 519537 61427 519571
rect 61393 519197 61427 519231
rect 55965 518925 55999 518959
rect 75285 519673 75319 519707
rect 65533 519605 65567 519639
rect 65533 519061 65567 519095
rect 75101 519605 75135 519639
rect 75193 519537 75227 519571
rect 75193 519197 75227 519231
rect 75101 519061 75135 519095
rect 65441 518925 65475 518959
rect 84761 519673 84795 519707
rect 80713 519537 80747 519571
rect 80713 519197 80747 519231
rect 75285 518925 75319 518959
rect 94605 519673 94639 519707
rect 84853 519605 84887 519639
rect 84853 519061 84887 519095
rect 94421 519605 94455 519639
rect 94513 519537 94547 519571
rect 94513 519197 94547 519231
rect 94421 519061 94455 519095
rect 84761 518925 84795 518959
rect 104081 519673 104115 519707
rect 100033 519537 100067 519571
rect 100033 519197 100067 519231
rect 94605 518925 94639 518959
rect 113925 519673 113959 519707
rect 104173 519605 104207 519639
rect 104173 519061 104207 519095
rect 113741 519605 113775 519639
rect 113833 519537 113867 519571
rect 113833 519197 113867 519231
rect 113741 519061 113775 519095
rect 104081 518925 104115 518959
rect 123401 519673 123435 519707
rect 119353 519537 119387 519571
rect 119353 519197 119387 519231
rect 113925 518925 113959 518959
rect 133245 519673 133279 519707
rect 123493 519605 123527 519639
rect 123493 519061 123527 519095
rect 133061 519605 133095 519639
rect 133153 519537 133187 519571
rect 133153 519197 133187 519231
rect 133061 519061 133095 519095
rect 123401 518925 123435 518959
rect 142721 519673 142755 519707
rect 138673 519537 138707 519571
rect 138673 519197 138707 519231
rect 133245 518925 133279 518959
rect 152565 519673 152599 519707
rect 142813 519605 142847 519639
rect 142813 519061 142847 519095
rect 152381 519605 152415 519639
rect 152473 519537 152507 519571
rect 152473 519197 152507 519231
rect 152381 519061 152415 519095
rect 142721 518925 142755 518959
rect 162041 519673 162075 519707
rect 157993 519537 158027 519571
rect 157993 519197 158027 519231
rect 152565 518925 152599 518959
rect 171701 519673 171735 519707
rect 162133 519605 162167 519639
rect 162133 519061 162167 519095
rect 171793 519605 171827 519639
rect 171793 519197 171827 519231
rect 171701 519061 171735 519095
rect 162041 518925 162075 518959
rect 181545 519741 181579 519775
rect 181361 519673 181395 519707
rect 171885 518925 171919 518959
rect 179429 519537 179463 519571
rect 181453 519605 181487 519639
rect 181453 519197 181487 519231
rect 181361 519061 181395 519095
rect 209973 519741 210007 519775
rect 181545 518925 181579 518959
rect 188353 519673 188387 519707
rect 200681 519673 200715 519707
rect 191113 519605 191147 519639
rect 190009 519537 190043 519571
rect 190009 519197 190043 519231
rect 195989 519537 196023 519571
rect 195989 519197 196023 519231
rect 191113 519061 191147 519095
rect 188353 518925 188387 518959
rect 209881 519673 209915 519707
rect 200773 519605 200807 519639
rect 209789 519605 209823 519639
rect 209789 519197 209823 519231
rect 200773 519061 200807 519095
rect 209789 519061 209823 519095
rect 200681 518925 200715 518959
rect 209789 518925 209823 518959
rect 219173 519741 219207 519775
rect 219265 519673 219299 519707
rect 219357 519605 219391 519639
rect 219357 519197 219391 519231
rect 305377 519605 305411 519639
rect 316877 519605 316911 519639
rect 325893 519469 325927 519503
rect 325801 519401 325835 519435
rect 305377 519197 305411 519231
rect 316785 519197 316819 519231
rect 316877 519197 316911 519231
rect 325709 519333 325743 519367
rect 325709 519197 325743 519231
rect 306849 519129 306883 519163
rect 307033 519129 307067 519163
rect 219357 519061 219391 519095
rect 307125 519061 307159 519095
rect 316693 519061 316727 519095
rect 316785 519061 316819 519095
rect 325709 519061 325743 519095
rect 219357 518925 219391 518959
rect 306849 518925 306883 518959
rect 316693 518925 316727 518959
rect 325709 518925 325743 518959
rect 335185 519469 335219 519503
rect 335277 519401 335311 519435
rect 349997 519265 350031 519299
rect 335277 519061 335311 519095
rect 345121 519129 345155 519163
rect 349997 519061 350031 519095
rect 351837 519265 351871 519299
rect 335277 518925 335311 518959
rect 345029 518925 345063 518959
rect 355149 519265 355183 519299
rect 355149 518993 355183 519027
rect 351837 518245 351871 518279
rect 179429 518177 179463 518211
rect 339417 218161 339451 218195
rect 329297 218025 329331 218059
rect 275845 217957 275879 217991
rect 275937 217957 275971 217991
rect 283113 217889 283147 217923
rect 281549 217821 281583 217855
rect 170873 217685 170907 217719
rect 168297 217481 168331 217515
rect 170781 217481 170815 217515
rect 170873 217481 170907 217515
rect 170965 217685 170999 217719
rect 167193 217413 167227 217447
rect 168481 217413 168515 217447
rect 180165 217685 180199 217719
rect 167009 217345 167043 217379
rect 167101 217345 167135 217379
rect 167285 217277 167319 217311
rect 212365 217685 212399 217719
rect 281549 217685 281583 217719
rect 281733 217821 281767 217855
rect 181453 217277 181487 217311
rect 181453 216665 181487 216699
rect 180165 212517 180199 212551
rect 281733 217413 281767 217447
rect 281825 217413 281859 217447
rect 281825 217141 281859 217175
rect 282929 217345 282963 217379
rect 282009 217073 282043 217107
rect 282009 216869 282043 216903
rect 321569 217889 321603 217923
rect 292589 217685 292623 217719
rect 292681 217413 292715 217447
rect 295349 217617 295383 217651
rect 291209 217277 291243 217311
rect 283113 216801 283147 216835
rect 289829 216869 289863 216903
rect 282929 216733 282963 216767
rect 320005 217481 320039 217515
rect 321569 217481 321603 217515
rect 323593 217889 323627 217923
rect 329297 217889 329331 217923
rect 332333 218025 332367 218059
rect 332333 217821 332367 217855
rect 332425 217821 332459 217855
rect 323593 217481 323627 217515
rect 331137 217549 331171 217583
rect 319913 217209 319947 217243
rect 320005 217209 320039 217243
rect 295349 217005 295383 217039
rect 302157 217073 302191 217107
rect 291209 216733 291243 216767
rect 291945 216801 291979 216835
rect 289829 216665 289863 216699
rect 212365 212517 212399 212551
rect 216965 215305 216999 215339
rect 299397 216801 299431 216835
rect 302157 216801 302191 216835
rect 307217 217005 307251 217039
rect 319913 217005 319947 217039
rect 311909 216937 311943 216971
rect 308413 216869 308447 216903
rect 308689 216869 308723 216903
rect 307217 216801 307251 216835
rect 311909 216733 311943 216767
rect 299397 216665 299431 216699
rect 335369 217821 335403 217855
rect 337853 217821 337887 217855
rect 335369 217413 335403 217447
rect 336657 217685 336691 217719
rect 337485 217685 337519 217719
rect 336657 217413 336691 217447
rect 332425 217345 332459 217379
rect 340613 218025 340647 218059
rect 340705 217957 340739 217991
rect 340613 217821 340647 217855
rect 339509 217685 339543 217719
rect 339509 217413 339543 217447
rect 340705 217413 340739 217447
rect 339417 217345 339451 217379
rect 350549 217889 350583 217923
rect 350549 217753 350583 217787
rect 340797 217345 340831 217379
rect 369777 217685 369811 217719
rect 340521 217277 340555 217311
rect 369777 216733 369811 216767
rect 331137 216665 331171 216699
rect 291945 215169 291979 215203
rect 216965 212517 216999 212551
rect 211905 212449 211939 212483
rect 211905 202861 211939 202895
rect 217057 211089 217091 211123
rect 262597 211089 262631 211123
rect 258273 207689 258307 207723
rect 219817 205649 219851 205683
rect 219817 202861 219851 202895
rect 328101 211089 328135 211123
rect 262597 205581 262631 205615
rect 315865 205649 315899 205683
rect 258273 202861 258307 202895
rect 343281 211089 343315 211123
rect 328101 205581 328135 205615
rect 329389 209729 329423 209763
rect 315865 202861 315899 202895
rect 217057 201501 217091 201535
rect 343281 205581 343315 205615
rect 344569 211089 344603 211123
rect 344569 205581 344603 205615
rect 192125 201433 192159 201467
rect 171517 195993 171551 196027
rect 171517 193205 171551 193239
rect 282837 201433 282871 201467
rect 329389 201433 329423 201467
rect 362509 201433 362543 201467
rect 192125 193137 192159 193171
rect 277225 200073 277259 200107
rect 262505 191777 262539 191811
rect 179981 188989 180015 189023
rect 182189 186337 182223 186371
rect 262505 186269 262539 186303
rect 282837 193137 282871 193171
rect 315773 196061 315807 196095
rect 315773 191845 315807 191879
rect 328193 193069 328227 193103
rect 277225 183549 277259 183583
rect 315681 191709 315715 191743
rect 182189 182189 182223 182223
rect 362509 191845 362543 191879
rect 328193 186269 328227 186303
rect 329573 191777 329607 191811
rect 315681 182189 315715 182223
rect 192217 182121 192251 182155
rect 179981 179401 180015 179435
rect 182189 181985 182223 182019
rect 176945 179333 176979 179367
rect 176945 173145 176979 173179
rect 181085 179333 181119 179367
rect 182189 176545 182223 176579
rect 224049 182121 224083 182155
rect 192217 176069 192251 176103
rect 217333 180761 217367 180795
rect 277133 182121 277167 182155
rect 224049 172533 224083 172567
rect 262597 182053 262631 182087
rect 262597 172533 262631 172567
rect 275845 180761 275879 180795
rect 217333 171105 217367 171139
rect 225429 172465 225463 172499
rect 181085 169745 181119 169779
rect 182189 171037 182223 171071
rect 177129 168317 177163 168351
rect 182189 161449 182223 161483
rect 211905 171037 211939 171071
rect 177129 158729 177163 158763
rect 181085 161381 181119 161415
rect 203165 161381 203199 161415
rect 182189 161313 182223 161347
rect 182189 156689 182223 156723
rect 192217 156757 192251 156791
rect 192217 153221 192251 153255
rect 181085 151793 181119 151827
rect 177129 149005 177163 149039
rect 177129 139485 177163 139519
rect 178141 149005 178175 149039
rect 211905 154581 211939 154615
rect 212457 164169 212491 164203
rect 229385 172465 229419 172499
rect 277133 172533 277167 172567
rect 285229 182121 285263 182155
rect 275845 171105 275879 171139
rect 229385 164169 229419 164203
rect 236377 171037 236411 171071
rect 225429 162673 225463 162707
rect 229293 162809 229327 162843
rect 212457 154581 212491 154615
rect 217149 161381 217183 161415
rect 217149 151793 217183 151827
rect 225613 158661 225647 158695
rect 225613 150297 225647 150331
rect 228189 157301 228223 157335
rect 203165 144857 203199 144891
rect 211905 144857 211939 144891
rect 181085 142069 181119 142103
rect 178141 139485 178175 139519
rect 179981 140709 180015 140743
rect 177129 139349 177163 139383
rect 177129 129761 177163 129795
rect 178141 139349 178175 139383
rect 181085 132549 181119 132583
rect 182189 142069 182223 142103
rect 179981 131189 180015 131223
rect 181085 132413 181119 132447
rect 178141 129761 178175 129795
rect 171425 125545 171459 125579
rect 171425 115957 171459 115991
rect 173081 125545 173115 125579
rect 194885 140709 194919 140743
rect 211905 135269 211939 135303
rect 212273 140709 212307 140743
rect 203073 133977 203107 134011
rect 194885 131121 194919 131155
rect 201785 133841 201819 133875
rect 182189 124185 182223 124219
rect 203073 132481 203107 132515
rect 354229 191777 354263 191811
rect 354229 183481 354263 183515
rect 329573 181577 329607 181611
rect 354321 182121 354355 182155
rect 355609 182121 355643 182155
rect 355609 176613 355643 176647
rect 362417 182121 362451 182155
rect 354321 176545 354355 176579
rect 362417 171173 362451 171207
rect 362417 171037 362451 171071
rect 285229 166889 285263 166923
rect 318441 169133 318475 169167
rect 318441 164237 318475 164271
rect 344569 167501 344603 167535
rect 236377 160157 236411 160191
rect 258273 164169 258307 164203
rect 355609 167025 355643 167059
rect 355609 164237 355643 164271
rect 344569 162877 344603 162911
rect 258273 157301 258307 157335
rect 261125 162809 261159 162843
rect 229293 153221 229327 153255
rect 261125 153221 261159 153255
rect 286701 162809 286735 162843
rect 317153 162809 317187 162843
rect 317153 157301 317187 157335
rect 318441 162809 318475 162843
rect 318441 157301 318475 157335
rect 341993 162809 342027 162843
rect 286701 153221 286735 153255
rect 291945 154513 291979 154547
rect 230949 153153 230983 153187
rect 354321 162809 354355 162843
rect 345673 161381 345707 161415
rect 341993 153221 342027 153255
rect 343281 158661 343315 158695
rect 291945 144993 291979 145027
rect 299213 147781 299247 147815
rect 299213 144925 299247 144959
rect 300501 147781 300535 147815
rect 300501 144925 300535 144959
rect 317245 147645 317279 147679
rect 230949 144857 230983 144891
rect 258273 144857 258307 144891
rect 228189 139417 228223 139451
rect 236285 142069 236319 142103
rect 212273 131121 212307 131155
rect 201785 124185 201819 124219
rect 211905 125545 211939 125579
rect 181085 122825 181119 122859
rect 200313 124117 200347 124151
rect 182189 122757 182223 122791
rect 181177 122689 181211 122723
rect 180993 121397 181027 121431
rect 181177 121397 181211 121431
rect 173081 115957 173115 115991
rect 178325 120037 178359 120071
rect 182189 117997 182223 118031
rect 192309 122757 192343 122791
rect 180993 111877 181027 111911
rect 184029 115889 184063 115923
rect 178325 110449 178359 110483
rect 181085 111741 181119 111775
rect 171425 106233 171459 106267
rect 171425 96645 171459 96679
rect 173081 106233 173115 106267
rect 200313 115821 200347 115855
rect 203073 124117 203107 124151
rect 231041 124117 231075 124151
rect 229201 122757 229235 122791
rect 211905 115957 211939 115991
rect 212273 121397 212307 121431
rect 203073 114529 203107 114563
rect 192309 110381 192343 110415
rect 194885 114461 194919 114495
rect 184029 108817 184063 108851
rect 194885 104873 194919 104907
rect 201877 114461 201911 114495
rect 229201 117997 229235 118031
rect 231041 114529 231075 114563
rect 232237 122757 232271 122791
rect 328285 147645 328319 147679
rect 328285 144925 328319 144959
rect 317245 143565 317279 143599
rect 329573 144857 329607 144891
rect 258273 137921 258307 137955
rect 261125 143497 261159 143531
rect 261125 133909 261159 133943
rect 275845 143497 275879 143531
rect 285321 143497 285355 143531
rect 285321 137921 285355 137955
rect 286609 143497 286643 143531
rect 286609 137921 286643 137955
rect 289369 143497 289403 143531
rect 318441 143497 318475 143531
rect 289369 137921 289403 137955
rect 315865 142069 315899 142103
rect 275845 133909 275879 133943
rect 277225 133841 277259 133875
rect 236285 120649 236319 120683
rect 258273 125545 258307 125579
rect 235273 118677 235307 118711
rect 341993 142137 342027 142171
rect 341993 140777 342027 140811
rect 354321 157301 354355 157335
rect 355517 162809 355551 162843
rect 362417 161449 362451 161483
rect 355517 153221 355551 153255
rect 361221 160021 361255 160055
rect 345673 151793 345707 151827
rect 361221 150501 361255 150535
rect 362417 156621 362451 156655
rect 362417 144857 362451 144891
rect 343281 140777 343315 140811
rect 361405 142069 361439 142103
rect 329573 135269 329607 135303
rect 341717 139349 341751 139383
rect 318441 133977 318475 134011
rect 315865 132481 315899 132515
rect 318441 133841 318475 133875
rect 277225 124185 277259 124219
rect 299213 128469 299247 128503
rect 299213 124185 299247 124219
rect 300501 128469 300535 128503
rect 361405 132481 361439 132515
rect 345581 132413 345615 132447
rect 341717 129761 341751 129795
rect 343281 131053 343315 131087
rect 318441 125545 318475 125579
rect 328285 128333 328319 128367
rect 300501 124185 300535 124219
rect 328285 124185 328319 124219
rect 329573 125545 329607 125579
rect 258273 118609 258307 118643
rect 261125 124117 261159 124151
rect 235273 115957 235307 115991
rect 291945 124117 291979 124151
rect 277225 118745 277259 118779
rect 261125 114529 261159 114563
rect 273085 115889 273119 115923
rect 232237 113169 232271 113203
rect 212273 113101 212307 113135
rect 219817 113101 219851 113135
rect 217057 111673 217091 111707
rect 201877 104873 201911 104907
rect 211905 106233 211939 106267
rect 181085 102221 181119 102255
rect 182189 104737 182223 104771
rect 173081 96645 173115 96679
rect 177037 102085 177071 102119
rect 179981 102085 180015 102119
rect 177037 92497 177071 92531
rect 178049 95081 178083 95115
rect 277225 114529 277259 114563
rect 282745 115957 282779 115991
rect 282745 114529 282779 114563
rect 318533 124117 318567 124151
rect 291945 114529 291979 114563
rect 315865 118745 315899 118779
rect 315865 114529 315899 114563
rect 354413 128333 354447 128367
rect 354413 124185 354447 124219
rect 355701 128333 355735 128367
rect 355701 124185 355735 124219
rect 345581 122825 345615 122859
rect 343281 121465 343315 121499
rect 329573 115957 329607 115991
rect 362325 121397 362359 121431
rect 362325 115889 362359 115923
rect 318533 114529 318567 114563
rect 354229 114597 354263 114631
rect 273085 106301 273119 106335
rect 277225 114393 277259 114427
rect 219817 103581 219851 103615
rect 236285 106233 236319 106267
rect 217057 102153 217091 102187
rect 219725 103445 219759 103479
rect 211905 100045 211939 100079
rect 182189 99297 182223 99331
rect 217241 95353 217275 95387
rect 194885 95149 194919 95183
rect 179981 92497 180015 92531
rect 182189 93789 182223 93823
rect 178049 91069 178083 91103
rect 171425 86921 171459 86955
rect 171425 77265 171459 77299
rect 173081 86921 173115 86955
rect 194885 85561 194919 85595
rect 201877 86921 201911 86955
rect 182189 84201 182223 84235
rect 191113 84133 191147 84167
rect 179981 82773 180015 82807
rect 173081 77265 173115 77299
rect 178141 81345 178175 81379
rect 171425 67541 171459 67575
rect 171425 57953 171459 57987
rect 173081 67541 173115 67575
rect 184029 75837 184063 75871
rect 179981 73185 180015 73219
rect 181269 74477 181303 74511
rect 191113 74545 191147 74579
rect 192309 84133 192343 84167
rect 184029 66249 184063 66283
rect 225337 99637 225371 99671
rect 224049 99501 224083 99535
rect 224049 95217 224083 95251
rect 235273 99365 235307 99399
rect 235273 96645 235307 96679
rect 258273 106233 258307 106267
rect 354229 113169 354263 113203
rect 355609 113101 355643 113135
rect 341901 113033 341935 113067
rect 317245 109701 317279 109735
rect 277225 104941 277259 104975
rect 300501 109157 300535 109191
rect 258273 99297 258307 99331
rect 261125 104805 261159 104839
rect 236285 96645 236319 96679
rect 225337 95217 225371 95251
rect 261125 95217 261159 95251
rect 275845 104805 275879 104839
rect 275845 95217 275879 95251
rect 277133 104805 277167 104839
rect 277133 95217 277167 95251
rect 282745 104805 282779 104839
rect 282745 95217 282779 95251
rect 283941 104805 283975 104839
rect 315865 109089 315899 109123
rect 315865 104873 315899 104907
rect 299213 103513 299247 103547
rect 300501 103513 300535 103547
rect 299213 102221 299247 102255
rect 283941 95217 283975 95251
rect 315773 96917 315807 96951
rect 219725 93857 219759 93891
rect 318349 109361 318383 109395
rect 318349 104873 318383 104907
rect 329573 106233 329607 106267
rect 317245 96645 317279 96679
rect 341901 103513 341935 103547
rect 354413 109701 354447 109735
rect 329573 96645 329607 96679
rect 344477 103445 344511 103479
rect 355609 103513 355643 103547
rect 354413 96645 354447 96679
rect 344477 93857 344511 93891
rect 315773 86989 315807 87023
rect 355701 93789 355735 93823
rect 217241 84201 217275 84235
rect 236285 86921 236319 86955
rect 201877 77265 201911 77299
rect 203073 80665 203107 80699
rect 192309 66249 192343 66283
rect 194885 77197 194919 77231
rect 235273 80053 235307 80087
rect 232237 77265 232271 77299
rect 235273 77265 235307 77299
rect 232237 75905 232271 75939
rect 258273 86921 258307 86955
rect 262321 86921 262355 86955
rect 258273 77265 258307 77299
rect 260941 85493 260975 85527
rect 236285 75905 236319 75939
rect 283941 85493 283975 85527
rect 262321 77265 262355 77299
rect 282745 77333 282779 77367
rect 260941 75905 260975 75939
rect 282745 75905 282779 75939
rect 283941 75905 283975 75939
rect 289277 85493 289311 85527
rect 361221 93789 361255 93823
rect 361221 85493 361255 85527
rect 355701 84201 355735 84235
rect 343281 84133 343315 84167
rect 289277 75905 289311 75939
rect 318257 77537 318291 77571
rect 318257 75905 318291 75939
rect 203073 71077 203107 71111
rect 217149 75769 217183 75803
rect 194885 66249 194919 66283
rect 341993 74613 342027 74647
rect 345581 84133 345615 84167
rect 343281 74545 343315 74579
rect 344569 79305 344603 79339
rect 341993 73253 342027 73287
rect 217149 66249 217183 66283
rect 219725 70465 219759 70499
rect 361313 84133 361347 84167
rect 361313 79305 361347 79339
rect 362325 84133 362359 84167
rect 345581 74545 345615 74579
rect 355977 75837 356011 75871
rect 344569 67609 344603 67643
rect 362325 67609 362359 67643
rect 355977 67337 356011 67371
rect 219725 66249 219759 66283
rect 283941 66181 283975 66215
rect 181269 64889 181303 64923
rect 230765 65909 230799 65943
rect 178141 63529 178175 63563
rect 203073 64821 203107 64855
rect 173081 57953 173115 57987
rect 177037 63461 177071 63495
rect 177037 57885 177071 57919
rect 179981 63461 180015 63495
rect 200405 61421 200439 61455
rect 179981 53805 180015 53839
rect 181085 58633 181119 58667
rect 181085 53805 181119 53839
rect 183937 55165 183971 55199
rect 171425 48229 171459 48263
rect 201877 61421 201911 61455
rect 275753 63461 275787 63495
rect 230765 56593 230799 56627
rect 262505 57885 262539 57919
rect 203073 55233 203107 55267
rect 201877 53941 201911 53975
rect 228189 55165 228223 55199
rect 200405 48297 200439 48331
rect 183937 45577 183971 45611
rect 212457 48229 212491 48263
rect 171425 38641 171459 38675
rect 179981 45509 180015 45543
rect 201877 45509 201911 45543
rect 179981 35921 180015 35955
rect 181085 44081 181119 44115
rect 171333 28917 171367 28951
rect 182189 41429 182223 41463
rect 182189 27625 182223 27659
rect 189549 40681 189583 40715
rect 275753 53805 275787 53839
rect 277133 63461 277167 63495
rect 262505 48297 262539 48331
rect 283941 56661 283975 56695
rect 285321 66181 285355 66215
rect 285321 56593 285355 56627
rect 286609 66181 286643 66215
rect 286609 56593 286643 56627
rect 289369 66181 289403 66215
rect 289369 56593 289403 56627
rect 329573 66181 329607 66215
rect 329573 56593 329607 56627
rect 344477 64821 344511 64855
rect 277133 48297 277167 48331
rect 283941 56525 283975 56559
rect 283941 46937 283975 46971
rect 318349 56525 318383 56559
rect 355609 64821 355643 64855
rect 344477 55233 344511 55267
rect 345673 59993 345707 60027
rect 318349 46937 318383 46971
rect 344569 51765 344603 51799
rect 228189 46869 228223 46903
rect 232053 46869 232087 46903
rect 212457 37281 212491 37315
rect 219817 42449 219851 42483
rect 317153 46869 317187 46903
rect 273085 45509 273119 45543
rect 232053 37281 232087 37315
rect 258273 38573 258307 38607
rect 219817 35921 219851 35955
rect 273085 37145 273119 37179
rect 275845 38573 275879 38607
rect 317153 37281 317187 37315
rect 329389 42109 329423 42143
rect 354321 57885 354355 57919
rect 354321 48365 354355 48399
rect 355609 48297 355643 48331
rect 362325 57885 362359 57919
rect 362325 48297 362359 48331
rect 345673 46937 345707 46971
rect 354321 48229 354355 48263
rect 344569 41089 344603 41123
rect 354321 41089 354355 41123
rect 344661 38573 344695 38607
rect 329389 37281 329423 37315
rect 343373 37281 343407 37315
rect 275845 33201 275879 33235
rect 258273 31705 258307 31739
rect 328101 31773 328135 31807
rect 189549 27625 189583 27659
rect 200405 27625 200439 27659
rect 201877 27625 201911 27659
rect 236377 28917 236411 28951
rect 181085 26265 181119 26299
rect 200405 26265 200439 26299
rect 212273 27557 212307 27591
rect 171333 19329 171367 19363
rect 178141 26197 178175 26231
rect 178141 16609 178175 16643
rect 179981 26197 180015 26231
rect 194885 26197 194919 26231
rect 192125 19261 192159 19295
rect 182373 17969 182407 18003
rect 182373 17765 182407 17799
rect 179981 16609 180015 16643
rect 317153 28849 317187 28883
rect 236377 19329 236411 19363
rect 261125 27557 261159 27591
rect 212273 19261 212307 19295
rect 214297 19261 214331 19295
rect 194885 16609 194919 16643
rect 192125 9673 192159 9707
rect 212273 12529 212307 12563
rect 212273 9673 212307 9707
rect 261125 17969 261159 18003
rect 268761 27557 268795 27591
rect 268761 17969 268795 18003
rect 275937 27557 275971 27591
rect 275937 17969 275971 18003
rect 277133 27557 277167 27591
rect 228097 17901 228131 17935
rect 228281 17901 228315 17935
rect 214297 9673 214331 9707
rect 328101 27625 328135 27659
rect 329481 28917 329515 28951
rect 317153 19329 317187 19363
rect 362417 31841 362451 31875
rect 344661 28985 344695 29019
rect 361313 31773 361347 31807
rect 361313 28985 361347 29019
rect 362417 28985 362451 29019
rect 343373 28441 343407 28475
rect 329481 19329 329515 19363
rect 343281 27557 343315 27591
rect 291853 19261 291887 19295
rect 289277 13073 289311 13107
rect 277133 9673 277167 9707
rect 283941 9741 283975 9775
rect 283941 8313 283975 8347
rect 291853 9673 291887 9707
rect 328193 19261 328227 19295
rect 341901 18377 341935 18411
rect 341901 13753 341935 13787
rect 343281 13685 343315 13719
rect 344569 27557 344603 27591
rect 345673 27557 345707 27591
rect 354321 27557 354355 27591
rect 345673 17969 345707 18003
rect 352941 19261 352975 19295
rect 344569 13617 344603 13651
rect 328193 9673 328227 9707
rect 329481 12461 329515 12495
rect 354321 17969 354355 18003
rect 355517 27557 355551 27591
rect 355517 17969 355551 18003
rect 361221 27557 361255 27591
rect 361221 17969 361255 18003
rect 362509 19261 362543 19295
rect 352941 11713 352975 11747
rect 329481 9673 329515 9707
rect 362509 9673 362543 9707
rect 289277 8041 289311 8075
rect 238769 4029 238803 4063
rect 234721 3961 234755 3995
rect 225245 3893 225279 3927
rect 225153 3757 225187 3791
rect 225245 3757 225279 3791
rect 226349 3893 226383 3927
rect 225061 3485 225095 3519
rect 225153 3485 225187 3519
rect 224969 3349 225003 3383
rect 225061 3349 225095 3383
rect 238769 3825 238803 3859
rect 273085 4029 273119 4063
rect 278145 4029 278179 4063
rect 286057 4029 286091 4063
rect 286241 4029 286275 4063
rect 277961 3961 277995 3995
rect 273085 3825 273119 3859
rect 273177 3825 273211 3859
rect 234813 3689 234847 3723
rect 274373 3825 274407 3859
rect 273177 3621 273211 3655
rect 274189 3757 274223 3791
rect 274189 3621 274223 3655
rect 226349 3349 226383 3383
rect 228741 3417 228775 3451
rect 67925 3281 67959 3315
rect 67925 3009 67959 3043
rect 69581 3009 69615 3043
rect 69673 3213 69707 3247
rect 69765 3213 69799 3247
rect 74549 3281 74583 3315
rect 64889 2941 64923 2975
rect 64889 2805 64923 2839
rect 77769 3281 77803 3315
rect 78965 3281 78999 3315
rect 81357 3281 81391 3315
rect 78045 3077 78079 3111
rect 78965 3077 78999 3111
rect 79425 3145 79459 3179
rect 69673 2805 69707 2839
rect 69765 3009 69799 3043
rect 74549 3009 74583 3043
rect 79333 2941 79367 2975
rect 79425 2941 79459 2975
rect 79517 3145 79551 3179
rect 79333 2805 79367 2839
rect 69765 2737 69799 2771
rect 79517 2737 79551 2771
rect 82829 3281 82863 3315
rect 274373 3281 274407 3315
rect 275753 3485 275787 3519
rect 225061 3213 225095 3247
rect 228741 3213 228775 3247
rect 82553 3145 82587 3179
rect 275753 3145 275787 3179
rect 287897 4097 287931 4131
rect 287989 4097 288023 4131
rect 287529 3961 287563 3995
rect 287713 3961 287747 3995
rect 278145 3893 278179 3927
rect 278053 3689 278087 3723
rect 287713 3689 287747 3723
rect 287897 3689 287931 3723
rect 278053 3485 278087 3519
rect 297281 3417 297315 3451
rect 301605 3417 301639 3451
rect 364993 3417 365027 3451
rect 313565 3281 313599 3315
rect 280353 3213 280387 3247
rect 86049 3077 86083 3111
rect 278329 3077 278363 3111
rect 81357 2737 81391 2771
rect 84117 3009 84151 3043
rect 86049 2941 86083 2975
rect 95525 3009 95559 3043
rect 277869 3009 277903 3043
rect 278237 3009 278271 3043
rect 280353 3009 280387 3043
rect 297189 3213 297223 3247
rect 297465 3213 297499 3247
rect 301605 3213 301639 3247
rect 306297 3213 306331 3247
rect 297189 2941 297223 2975
rect 306297 2941 306331 2975
rect 308321 3077 308355 3111
rect 313565 3077 313599 3111
rect 364993 3009 365027 3043
rect 308321 2941 308355 2975
rect 121469 2873 121503 2907
rect 121653 2873 121687 2907
rect 95525 2805 95559 2839
rect 84117 2737 84151 2771
<< metal1 >>
rect 137830 700952 137836 701004
rect 137888 700992 137894 701004
rect 280154 700992 280160 701004
rect 137888 700964 280160 700992
rect 137888 700952 137894 700964
rect 280154 700952 280160 700964
rect 280212 700952 280218 701004
rect 262122 700884 262128 700936
rect 262180 700924 262186 700936
rect 413646 700924 413652 700936
rect 262180 700896 413652 700924
rect 262180 700884 262186 700896
rect 413646 700884 413652 700896
rect 413704 700884 413710 700936
rect 105446 700816 105452 700868
rect 105504 700856 105510 700868
rect 283006 700856 283012 700868
rect 105504 700828 283012 700856
rect 105504 700816 105510 700828
rect 283006 700816 283012 700828
rect 283064 700816 283070 700868
rect 89162 700748 89168 700800
rect 89220 700788 89226 700800
rect 287238 700788 287244 700800
rect 89220 700760 287244 700788
rect 89220 700748 89226 700760
rect 287238 700748 287244 700760
rect 287296 700748 287302 700800
rect 255222 700680 255228 700732
rect 255280 700720 255286 700732
rect 462314 700720 462320 700732
rect 255280 700692 462320 700720
rect 255280 700680 255286 700692
rect 462314 700680 462320 700692
rect 462372 700680 462378 700732
rect 72970 700612 72976 700664
rect 73028 700652 73034 700664
rect 284294 700652 284300 700664
rect 73028 700624 284300 700652
rect 73028 700612 73034 700624
rect 284294 700612 284300 700624
rect 284352 700612 284358 700664
rect 256602 700544 256608 700596
rect 256660 700584 256666 700596
rect 478506 700584 478512 700596
rect 256660 700556 478512 700584
rect 256660 700544 256666 700556
rect 478506 700544 478512 700556
rect 478564 700544 478570 700596
rect 40494 700476 40500 700528
rect 40552 700516 40558 700528
rect 288434 700516 288440 700528
rect 40552 700488 288440 700516
rect 40552 700476 40558 700488
rect 288434 700476 288440 700488
rect 288492 700476 288498 700528
rect 24302 700408 24308 700460
rect 24360 700448 24366 700460
rect 291381 700451 291439 700457
rect 291381 700448 291393 700451
rect 24360 700420 291393 700448
rect 24360 700408 24366 700420
rect 291381 700417 291393 700420
rect 291427 700417 291439 700451
rect 291381 700411 291439 700417
rect 249702 700340 249708 700392
rect 249760 700380 249766 700392
rect 527174 700380 527180 700392
rect 249760 700352 527180 700380
rect 249760 700340 249766 700352
rect 527174 700340 527180 700352
rect 527232 700340 527238 700392
rect 8110 700272 8116 700324
rect 8168 700312 8174 700324
rect 289998 700312 290004 700324
rect 8168 700284 290004 700312
rect 8168 700272 8174 700284
rect 289998 700272 290004 700284
rect 290056 700272 290062 700324
rect 335998 700272 336004 700324
rect 336056 700312 336062 700324
rect 429838 700312 429844 700324
rect 336056 700284 429844 700312
rect 336056 700272 336062 700284
rect 429838 700272 429844 700284
rect 429896 700272 429902 700324
rect 260742 700204 260748 700256
rect 260800 700244 260806 700256
rect 397454 700244 397460 700256
rect 260800 700216 397460 700244
rect 260800 700204 260806 700216
rect 397454 700204 397460 700216
rect 397512 700204 397518 700256
rect 154114 700136 154120 700188
rect 154172 700176 154178 700188
rect 281534 700176 281540 700188
rect 154172 700148 281540 700176
rect 154172 700136 154178 700148
rect 281534 700136 281540 700148
rect 281592 700136 281598 700188
rect 170306 700068 170312 700120
rect 170364 700108 170370 700120
rect 277394 700108 277400 700120
rect 170364 700080 277400 700108
rect 170364 700068 170370 700080
rect 277394 700068 277400 700080
rect 277452 700068 277458 700120
rect 279418 700068 279424 700120
rect 279476 700108 279482 700120
rect 364978 700108 364984 700120
rect 279476 700080 364984 700108
rect 279476 700068 279482 700080
rect 364978 700068 364984 700080
rect 365036 700068 365042 700120
rect 267642 700000 267648 700052
rect 267700 700040 267706 700052
rect 269114 700040 269120 700052
rect 267700 700012 269120 700040
rect 267700 700000 267706 700012
rect 269114 700000 269120 700012
rect 269172 700000 269178 700052
rect 269393 700043 269451 700049
rect 269393 700009 269405 700043
rect 269439 700040 269451 700043
rect 348786 700040 348792 700052
rect 269439 700012 348792 700040
rect 269439 700009 269451 700012
rect 269393 700003 269451 700009
rect 348786 700000 348792 700012
rect 348844 700000 348850 700052
rect 202782 699932 202788 699984
rect 202840 699972 202846 699984
rect 274634 699972 274640 699984
rect 202840 699944 274640 699972
rect 202840 699932 202846 699944
rect 274634 699932 274640 699944
rect 274692 699932 274698 699984
rect 264882 699864 264888 699916
rect 264940 699904 264946 699916
rect 332502 699904 332508 699916
rect 264940 699876 332508 699904
rect 264940 699864 264946 699876
rect 332502 699864 332508 699876
rect 332560 699864 332566 699916
rect 218974 699796 218980 699848
rect 219032 699836 219038 699848
rect 276014 699836 276020 699848
rect 219032 699808 276020 699836
rect 219032 699796 219038 699808
rect 276014 699796 276020 699808
rect 276072 699796 276078 699848
rect 235166 699728 235172 699780
rect 235224 699768 235230 699780
rect 273254 699768 273260 699780
rect 235224 699740 273260 699768
rect 235224 699728 235230 699740
rect 273254 699728 273260 699740
rect 273312 699728 273318 699780
rect 267642 699660 267648 699712
rect 267700 699700 267706 699712
rect 269393 699703 269451 699709
rect 269393 699700 269405 699703
rect 267700 699672 269405 699700
rect 267700 699660 267706 699672
rect 269393 699669 269405 699672
rect 269439 699669 269451 699703
rect 269393 699663 269451 699669
rect 271782 699660 271788 699712
rect 271840 699700 271846 699712
rect 283834 699700 283840 699712
rect 271840 699672 283840 699700
rect 271840 699660 271846 699672
rect 283834 699660 283840 699672
rect 283892 699660 283898 699712
rect 291378 698204 291384 698216
rect 291339 698176 291384 698204
rect 291378 698164 291384 698176
rect 291436 698164 291442 698216
rect 245562 696940 245568 696992
rect 245620 696980 245626 696992
rect 579890 696980 579896 696992
rect 245620 696952 579896 696980
rect 245620 696940 245626 696952
rect 579890 696940 579896 696952
rect 579948 696940 579954 696992
rect 269209 695487 269267 695493
rect 269209 695453 269221 695487
rect 269255 695484 269267 695487
rect 269298 695484 269304 695496
rect 269255 695456 269304 695484
rect 269255 695453 269267 695456
rect 269209 695447 269267 695453
rect 269298 695444 269304 695456
rect 269356 695444 269362 695496
rect 287149 695487 287207 695493
rect 287149 695453 287161 695487
rect 287195 695484 287207 695487
rect 287238 695484 287244 695496
rect 287195 695456 287244 695484
rect 287195 695453 287207 695456
rect 287149 695447 287207 695453
rect 287238 695444 287244 695456
rect 287296 695444 287302 695496
rect 289909 695487 289967 695493
rect 289909 695453 289921 695487
rect 289955 695484 289967 695487
rect 289998 695484 290004 695496
rect 289955 695456 290004 695484
rect 289955 695453 289967 695456
rect 289909 695447 289967 695453
rect 289998 695444 290004 695456
rect 290056 695444 290062 695496
rect 291378 695484 291384 695496
rect 291339 695456 291384 695484
rect 291378 695444 291384 695456
rect 291436 695444 291442 695496
rect 267553 688755 267611 688761
rect 267553 688721 267565 688755
rect 267599 688752 267611 688755
rect 267642 688752 267648 688764
rect 267599 688724 267648 688752
rect 267599 688721 267611 688724
rect 267553 688715 267611 688721
rect 267642 688712 267648 688724
rect 267700 688712 267706 688764
rect 252278 688576 252284 688628
rect 252336 688616 252342 688628
rect 252462 688616 252468 688628
rect 252336 688588 252468 688616
rect 252336 688576 252342 688588
rect 252462 688576 252468 688588
rect 252520 688576 252526 688628
rect 289906 688616 289912 688628
rect 289867 688588 289912 688616
rect 289906 688576 289912 688588
rect 289964 688576 289970 688628
rect 291378 688616 291384 688628
rect 291339 688588 291384 688616
rect 291378 688576 291384 688588
rect 291436 688576 291442 688628
rect 299658 688576 299664 688628
rect 299716 688616 299722 688628
rect 300118 688616 300124 688628
rect 299716 688588 300124 688616
rect 299716 688576 299722 688588
rect 300118 688576 300124 688588
rect 300176 688576 300182 688628
rect 559098 688576 559104 688628
rect 559156 688616 559162 688628
rect 559650 688616 559656 688628
rect 559156 688588 559656 688616
rect 559156 688576 559162 688588
rect 559650 688576 559656 688588
rect 559708 688576 559714 688628
rect 287146 688344 287152 688356
rect 287107 688316 287152 688344
rect 287146 688304 287152 688316
rect 287204 688304 287210 688356
rect 267550 685964 267556 685976
rect 267511 685936 267556 685964
rect 267550 685924 267556 685936
rect 267608 685924 267614 685976
rect 269206 685964 269212 685976
rect 269167 685936 269212 685964
rect 269206 685924 269212 685936
rect 269264 685924 269270 685976
rect 299492 685936 301268 685964
rect 246942 685856 246948 685908
rect 247000 685896 247006 685908
rect 299492 685896 299520 685936
rect 247000 685868 299520 685896
rect 301240 685896 301268 685936
rect 552584 685936 559788 685964
rect 552584 685896 552612 685936
rect 301240 685868 552612 685896
rect 559760 685896 559788 685936
rect 580074 685896 580080 685908
rect 559760 685868 580080 685896
rect 247000 685856 247006 685868
rect 580074 685856 580080 685868
rect 580132 685856 580138 685908
rect 252373 685831 252431 685837
rect 252373 685797 252385 685831
rect 252419 685828 252431 685831
rect 252462 685828 252468 685840
rect 252419 685800 252468 685828
rect 252419 685797 252431 685800
rect 252373 685791 252431 685797
rect 252462 685788 252468 685800
rect 252520 685788 252526 685840
rect 267550 684468 267556 684480
rect 267511 684440 267556 684468
rect 267550 684428 267556 684440
rect 267608 684428 267614 684480
rect 269206 684468 269212 684480
rect 269167 684440 269212 684468
rect 269206 684428 269212 684440
rect 269264 684428 269270 684480
rect 299566 684428 299572 684480
rect 299624 684468 299630 684480
rect 299845 684471 299903 684477
rect 299845 684468 299857 684471
rect 299624 684440 299857 684468
rect 299624 684428 299630 684440
rect 299845 684437 299857 684440
rect 299891 684437 299903 684471
rect 299845 684431 299903 684437
rect 559006 684428 559012 684480
rect 559064 684468 559070 684480
rect 559285 684471 559343 684477
rect 559285 684468 559297 684471
rect 559064 684440 559297 684468
rect 559064 684428 559070 684440
rect 559285 684437 559297 684440
rect 559331 684437 559343 684471
rect 559285 684431 559343 684437
rect 276014 683136 276020 683188
rect 276072 683176 276078 683188
rect 276198 683176 276204 683188
rect 276072 683148 276204 683176
rect 276072 683136 276078 683148
rect 276198 683136 276204 683148
rect 276256 683136 276262 683188
rect 267553 682975 267611 682981
rect 267553 682941 267565 682975
rect 267599 682972 267611 682975
rect 267642 682972 267648 682984
rect 267599 682944 267648 682972
rect 267599 682941 267611 682944
rect 267553 682935 267611 682941
rect 267642 682932 267648 682944
rect 267700 682932 267706 682984
rect 3510 681708 3516 681760
rect 3568 681748 3574 681760
rect 292574 681748 292580 681760
rect 3568 681720 292580 681748
rect 3568 681708 3574 681720
rect 292574 681708 292580 681720
rect 292632 681708 292638 681760
rect 291470 679028 291476 679040
rect 291396 679000 291476 679028
rect 291396 678972 291424 679000
rect 291470 678988 291476 679000
rect 291528 678988 291534 679040
rect 291378 678920 291384 678972
rect 291436 678920 291442 678972
rect 252370 676240 252376 676252
rect 252331 676212 252376 676240
rect 252370 676200 252376 676212
rect 252428 676200 252434 676252
rect 269209 676243 269267 676249
rect 269209 676209 269221 676243
rect 269255 676240 269267 676243
rect 269298 676240 269304 676252
rect 269255 676212 269304 676240
rect 269255 676209 269267 676212
rect 269209 676203 269267 676209
rect 269298 676200 269304 676212
rect 269356 676200 269362 676252
rect 287149 676175 287207 676181
rect 287149 676141 287161 676175
rect 287195 676172 287207 676175
rect 287238 676172 287244 676184
rect 287195 676144 287244 676172
rect 287195 676141 287207 676144
rect 287149 676135 287207 676141
rect 287238 676132 287244 676144
rect 287296 676132 287302 676184
rect 494054 676172 494060 676184
rect 494015 676144 494060 676172
rect 494054 676132 494060 676144
rect 494112 676132 494118 676184
rect 267369 674815 267427 674821
rect 267369 674781 267381 674815
rect 267415 674812 267427 674815
rect 267642 674812 267648 674824
rect 267415 674784 267648 674812
rect 267415 674781 267427 674784
rect 267369 674775 267427 674781
rect 267642 674772 267648 674784
rect 267700 674772 267706 674824
rect 242802 673480 242808 673532
rect 242860 673520 242866 673532
rect 580258 673520 580264 673532
rect 242860 673492 580264 673520
rect 242860 673480 242866 673492
rect 580258 673480 580264 673492
rect 580316 673480 580322 673532
rect 269298 669332 269304 669384
rect 269356 669332 269362 669384
rect 252278 669264 252284 669316
rect 252336 669304 252342 669316
rect 252462 669304 252468 669316
rect 252336 669276 252468 669304
rect 252336 669264 252342 669276
rect 252462 669264 252468 669276
rect 252520 669264 252526 669316
rect 269316 669236 269344 669332
rect 276014 669264 276020 669316
rect 276072 669304 276078 669316
rect 276198 669304 276204 669316
rect 276072 669276 276204 669304
rect 276072 669264 276078 669276
rect 276198 669264 276204 669276
rect 276256 669264 276262 669316
rect 269390 669236 269396 669248
rect 269316 669208 269396 669236
rect 269390 669196 269396 669208
rect 269448 669196 269454 669248
rect 3418 667904 3424 667956
rect 3476 667944 3482 667956
rect 296714 667944 296720 667956
rect 3476 667916 296720 667944
rect 3476 667904 3482 667916
rect 296714 667904 296720 667916
rect 296772 667904 296778 667956
rect 287146 666584 287152 666596
rect 287107 666556 287152 666584
rect 287146 666544 287152 666556
rect 287204 666544 287210 666596
rect 299845 666587 299903 666593
rect 299845 666553 299857 666587
rect 299891 666584 299903 666587
rect 299934 666584 299940 666596
rect 299891 666556 299940 666584
rect 299891 666553 299903 666556
rect 299845 666547 299903 666553
rect 299934 666544 299940 666556
rect 299992 666544 299998 666596
rect 494057 666587 494115 666593
rect 494057 666553 494069 666587
rect 494103 666584 494115 666587
rect 494146 666584 494152 666596
rect 494103 666556 494152 666584
rect 494103 666553 494115 666556
rect 494057 666547 494115 666553
rect 494146 666544 494152 666556
rect 494204 666544 494210 666596
rect 559285 666587 559343 666593
rect 559285 666553 559297 666587
rect 559331 666584 559343 666587
rect 559374 666584 559380 666596
rect 559331 666556 559380 666584
rect 559331 666553 559343 666556
rect 559285 666547 559343 666553
rect 559374 666544 559380 666556
rect 559432 666544 559438 666596
rect 252373 666519 252431 666525
rect 252373 666485 252385 666519
rect 252419 666516 252431 666519
rect 252462 666516 252468 666528
rect 252419 666488 252468 666516
rect 252419 666485 252431 666488
rect 252373 666479 252431 666485
rect 252462 666476 252468 666488
rect 252520 666476 252526 666528
rect 276109 666519 276167 666525
rect 276109 666485 276121 666519
rect 276155 666516 276167 666519
rect 276198 666516 276204 666528
rect 276155 666488 276204 666516
rect 276155 666485 276167 666488
rect 276109 666479 276167 666485
rect 276198 666476 276204 666488
rect 276256 666476 276262 666528
rect 289814 666476 289820 666528
rect 289872 666516 289878 666528
rect 289872 666488 289917 666516
rect 289872 666476 289878 666488
rect 267366 665292 267372 665304
rect 267327 665264 267372 665292
rect 267366 665252 267372 665264
rect 267424 665252 267430 665304
rect 267366 665116 267372 665168
rect 267424 665156 267430 665168
rect 267553 665159 267611 665165
rect 267553 665156 267565 665159
rect 267424 665128 267565 665156
rect 267424 665116 267430 665128
rect 267553 665125 267565 665128
rect 267599 665125 267611 665159
rect 267553 665119 267611 665125
rect 269390 663728 269396 663740
rect 269351 663700 269396 663728
rect 269390 663688 269396 663700
rect 269448 663688 269454 663740
rect 267550 659580 267556 659592
rect 267511 659552 267556 659580
rect 267550 659540 267556 659552
rect 267608 659540 267614 659592
rect 252370 656928 252376 656940
rect 252331 656900 252376 656928
rect 252370 656888 252376 656900
rect 252428 656888 252434 656940
rect 276106 656928 276112 656940
rect 276067 656900 276112 656928
rect 276106 656888 276112 656900
rect 276164 656888 276170 656940
rect 289814 656888 289820 656940
rect 289872 656928 289878 656940
rect 289872 656900 289917 656928
rect 289872 656888 289878 656900
rect 494054 654100 494060 654152
rect 494112 654140 494118 654152
rect 494238 654140 494244 654152
rect 494112 654112 494244 654140
rect 494112 654100 494118 654112
rect 494238 654100 494244 654112
rect 494296 654100 494302 654152
rect 3050 652740 3056 652792
rect 3108 652780 3114 652792
rect 295334 652780 295340 652792
rect 3108 652752 295340 652780
rect 3108 652740 3114 652752
rect 295334 652740 295340 652752
rect 295392 652740 295398 652792
rect 267461 650199 267519 650205
rect 267461 650165 267473 650199
rect 267507 650196 267519 650199
rect 267550 650196 267556 650208
rect 267507 650168 267556 650196
rect 267507 650165 267519 650168
rect 267461 650159 267519 650165
rect 267550 650156 267556 650168
rect 267608 650156 267614 650208
rect 240042 650020 240048 650072
rect 240100 650060 240106 650072
rect 579890 650060 579896 650072
rect 240100 650032 579896 650060
rect 240100 650020 240106 650032
rect 579890 650020 579896 650032
rect 579948 650020 579954 650072
rect 252278 649952 252284 650004
rect 252336 649992 252342 650004
rect 252462 649992 252468 650004
rect 252336 649964 252468 649992
rect 252336 649952 252342 649964
rect 252462 649952 252468 649964
rect 252520 649952 252526 650004
rect 269390 649924 269396 649936
rect 269351 649896 269396 649924
rect 269390 649884 269396 649896
rect 269448 649884 269454 649936
rect 287238 649884 287244 649936
rect 287296 649884 287302 649936
rect 287256 649800 287284 649884
rect 287238 649748 287244 649800
rect 287296 649748 287302 649800
rect 299658 647232 299664 647284
rect 299716 647272 299722 647284
rect 299750 647272 299756 647284
rect 299716 647244 299756 647272
rect 299716 647232 299722 647244
rect 299750 647232 299756 647244
rect 299808 647232 299814 647284
rect 559098 647232 559104 647284
rect 559156 647272 559162 647284
rect 559190 647272 559196 647284
rect 559156 647244 559196 647272
rect 559156 647232 559162 647244
rect 559190 647232 559196 647244
rect 559248 647232 559254 647284
rect 252373 647207 252431 647213
rect 252373 647173 252385 647207
rect 252419 647204 252431 647207
rect 252462 647204 252468 647216
rect 252419 647176 252468 647204
rect 252419 647173 252431 647176
rect 252373 647167 252431 647173
rect 252462 647164 252468 647176
rect 252520 647164 252526 647216
rect 289814 647164 289820 647216
rect 289872 647204 289878 647216
rect 289872 647176 289917 647204
rect 289872 647164 289878 647176
rect 267458 645912 267464 645924
rect 267419 645884 267464 645912
rect 267458 645872 267464 645884
rect 267516 645872 267522 645924
rect 276014 644444 276020 644496
rect 276072 644484 276078 644496
rect 276198 644484 276204 644496
rect 276072 644456 276204 644484
rect 276072 644444 276078 644456
rect 276198 644444 276204 644456
rect 276256 644444 276262 644496
rect 269390 640404 269396 640416
rect 269316 640376 269396 640404
rect 269316 640280 269344 640376
rect 269390 640364 269396 640376
rect 269448 640364 269454 640416
rect 299658 640364 299664 640416
rect 299716 640404 299722 640416
rect 299750 640404 299756 640416
rect 299716 640376 299756 640404
rect 299716 640364 299722 640376
rect 299750 640364 299756 640376
rect 299808 640364 299814 640416
rect 559098 640364 559104 640416
rect 559156 640404 559162 640416
rect 559190 640404 559196 640416
rect 559156 640376 559196 640404
rect 559156 640364 559162 640376
rect 559190 640364 559196 640376
rect 559248 640364 559254 640416
rect 269298 640228 269304 640280
rect 269356 640228 269362 640280
rect 241422 638936 241428 638988
rect 241480 638976 241486 638988
rect 580074 638976 580080 638988
rect 241480 638948 580080 638976
rect 241480 638936 241486 638948
rect 580074 638936 580080 638948
rect 580132 638936 580138 638988
rect 252370 637616 252376 637628
rect 252331 637588 252376 637616
rect 252370 637576 252376 637588
rect 252428 637576 252434 637628
rect 289814 637576 289820 637628
rect 289872 637616 289878 637628
rect 289872 637588 289917 637616
rect 289872 637576 289878 637588
rect 291289 637551 291347 637557
rect 291289 637517 291301 637551
rect 291335 637548 291347 637551
rect 291378 637548 291384 637560
rect 291335 637520 291384 637548
rect 291335 637517 291347 637520
rect 291289 637511 291347 637517
rect 291378 637508 291384 637520
rect 291436 637508 291442 637560
rect 494054 634788 494060 634840
rect 494112 634828 494118 634840
rect 494238 634828 494244 634840
rect 494112 634800 494244 634828
rect 494112 634788 494118 634800
rect 494238 634788 494244 634800
rect 494296 634788 494302 634840
rect 267461 630887 267519 630893
rect 267461 630853 267473 630887
rect 267507 630884 267519 630887
rect 267550 630884 267556 630896
rect 267507 630856 267556 630884
rect 267507 630853 267519 630856
rect 267461 630847 267519 630853
rect 267550 630844 267556 630856
rect 267608 630844 267614 630896
rect 287054 630640 287060 630692
rect 287112 630680 287118 630692
rect 287238 630680 287244 630692
rect 287112 630652 287244 630680
rect 287112 630640 287118 630652
rect 287238 630640 287244 630652
rect 287296 630640 287302 630692
rect 299566 630640 299572 630692
rect 299624 630680 299630 630692
rect 299750 630680 299756 630692
rect 299624 630652 299756 630680
rect 299624 630640 299630 630652
rect 299750 630640 299756 630652
rect 299808 630640 299814 630692
rect 559006 630640 559012 630692
rect 559064 630680 559070 630692
rect 559190 630680 559196 630692
rect 559064 630652 559196 630680
rect 559064 630640 559070 630652
rect 559190 630640 559196 630652
rect 559248 630640 559254 630692
rect 291286 627960 291292 627972
rect 291247 627932 291292 627960
rect 291286 627920 291292 627932
rect 291344 627920 291350 627972
rect 289906 627892 289912 627904
rect 289867 627864 289912 627892
rect 289906 627852 289912 627864
rect 289964 627852 289970 627904
rect 267458 626668 267464 626680
rect 267419 626640 267464 626668
rect 267458 626628 267464 626640
rect 267516 626628 267522 626680
rect 238662 626560 238668 626612
rect 238720 626600 238726 626612
rect 580258 626600 580264 626612
rect 238720 626572 580264 626600
rect 238720 626560 238726 626572
rect 580258 626560 580264 626572
rect 580316 626560 580322 626612
rect 3418 623772 3424 623824
rect 3476 623812 3482 623824
rect 298094 623812 298100 623824
rect 3476 623784 298100 623812
rect 3476 623772 3482 623784
rect 298094 623772 298100 623784
rect 298152 623772 298158 623824
rect 267458 623092 267464 623144
rect 267516 623132 267522 623144
rect 267550 623132 267556 623144
rect 267516 623104 267556 623132
rect 267516 623092 267522 623104
rect 267550 623092 267556 623104
rect 267608 623092 267614 623144
rect 289909 618307 289967 618313
rect 289909 618273 289921 618307
rect 289955 618304 289967 618307
rect 289998 618304 290004 618316
rect 289955 618276 290004 618304
rect 289955 618273 289967 618276
rect 289909 618267 289967 618273
rect 289998 618264 290004 618276
rect 290056 618264 290062 618316
rect 291289 618239 291347 618245
rect 291289 618205 291301 618239
rect 291335 618236 291347 618239
rect 291378 618236 291384 618248
rect 291335 618208 291384 618236
rect 291335 618205 291347 618208
rect 291289 618199 291347 618205
rect 291378 618196 291384 618208
rect 291436 618196 291442 618248
rect 257982 617516 257988 617568
rect 258040 617556 258046 617568
rect 335998 617556 336004 617568
rect 258040 617528 336004 617556
rect 258040 617516 258046 617528
rect 335998 617516 336004 617528
rect 336056 617516 336062 617568
rect 494054 615476 494060 615528
rect 494112 615516 494118 615528
rect 494238 615516 494244 615528
rect 494112 615488 494244 615516
rect 494112 615476 494118 615488
rect 494238 615476 494244 615488
rect 494296 615476 494302 615528
rect 269298 611396 269304 611448
rect 269356 611396 269362 611448
rect 269316 611312 269344 611396
rect 276014 611328 276020 611380
rect 276072 611368 276078 611380
rect 276198 611368 276204 611380
rect 276072 611340 276204 611368
rect 276072 611328 276078 611340
rect 276198 611328 276204 611340
rect 276256 611328 276262 611380
rect 287054 611328 287060 611380
rect 287112 611368 287118 611380
rect 287238 611368 287244 611380
rect 287112 611340 287244 611368
rect 287112 611328 287118 611340
rect 287238 611328 287244 611340
rect 287296 611328 287302 611380
rect 289814 611328 289820 611380
rect 289872 611368 289878 611380
rect 289998 611368 290004 611380
rect 289872 611340 290004 611368
rect 289872 611328 289878 611340
rect 289998 611328 290004 611340
rect 290056 611328 290062 611380
rect 299566 611328 299572 611380
rect 299624 611368 299630 611380
rect 299750 611368 299756 611380
rect 299624 611340 299756 611368
rect 299624 611328 299630 611340
rect 299750 611328 299756 611340
rect 299808 611328 299814 611380
rect 559006 611328 559012 611380
rect 559064 611368 559070 611380
rect 559190 611368 559196 611380
rect 559064 611340 559196 611368
rect 559064 611328 559070 611340
rect 559190 611328 559196 611340
rect 559248 611328 559254 611380
rect 269298 611260 269304 611312
rect 269356 611260 269362 611312
rect 3418 609968 3424 610020
rect 3476 610008 3482 610020
rect 302234 610008 302240 610020
rect 3476 609980 302240 610008
rect 3476 609968 3482 609980
rect 302234 609968 302240 609980
rect 302292 609968 302298 610020
rect 291286 608648 291292 608660
rect 291247 608620 291292 608648
rect 291286 608608 291292 608620
rect 291344 608608 291350 608660
rect 287146 608580 287152 608592
rect 287107 608552 287152 608580
rect 287146 608540 287152 608552
rect 287204 608540 287210 608592
rect 299658 608580 299664 608592
rect 299619 608552 299664 608580
rect 299658 608540 299664 608552
rect 299716 608540 299722 608592
rect 559098 608580 559104 608592
rect 559059 608552 559104 608580
rect 559098 608540 559104 608552
rect 559156 608540 559162 608592
rect 291286 607152 291292 607164
rect 291247 607124 291292 607152
rect 291286 607112 291292 607124
rect 291344 607112 291350 607164
rect 234522 603100 234528 603152
rect 234580 603140 234586 603152
rect 579890 603140 579896 603152
rect 234580 603112 579896 603140
rect 234580 603100 234586 603112
rect 579890 603100 579896 603112
rect 579948 603100 579954 603152
rect 276106 601740 276112 601792
rect 276164 601740 276170 601792
rect 269114 601672 269120 601724
rect 269172 601712 269178 601724
rect 269298 601712 269304 601724
rect 269172 601684 269304 601712
rect 269172 601672 269178 601684
rect 269298 601672 269304 601684
rect 269356 601672 269362 601724
rect 276124 601712 276152 601740
rect 276198 601712 276204 601724
rect 276124 601684 276204 601712
rect 276198 601672 276204 601684
rect 276256 601672 276262 601724
rect 299661 601715 299719 601721
rect 299661 601681 299673 601715
rect 299707 601712 299719 601715
rect 299842 601712 299848 601724
rect 299707 601684 299848 601712
rect 299707 601681 299719 601684
rect 299661 601675 299719 601681
rect 299842 601672 299848 601684
rect 299900 601672 299906 601724
rect 559101 601715 559159 601721
rect 559101 601681 559113 601715
rect 559147 601712 559159 601715
rect 559282 601712 559288 601724
rect 559147 601684 559288 601712
rect 559147 601681 559159 601684
rect 559101 601675 559159 601681
rect 559282 601672 559288 601684
rect 559340 601672 559346 601724
rect 287149 598995 287207 599001
rect 287149 598961 287161 598995
rect 287195 598992 287207 598995
rect 287238 598992 287244 599004
rect 287195 598964 287244 598992
rect 287195 598961 287207 598964
rect 287149 598955 287207 598961
rect 287238 598952 287244 598964
rect 287296 598952 287302 599004
rect 269114 598924 269120 598936
rect 269075 598896 269120 598924
rect 269114 598884 269120 598896
rect 269172 598884 269178 598936
rect 276198 598924 276204 598936
rect 276159 598896 276204 598924
rect 276198 598884 276204 598896
rect 276256 598884 276262 598936
rect 299753 598927 299811 598933
rect 299753 598893 299765 598927
rect 299799 598924 299811 598927
rect 299842 598924 299848 598936
rect 299799 598896 299848 598924
rect 299799 598893 299811 598896
rect 299753 598887 299811 598893
rect 299842 598884 299848 598896
rect 299900 598884 299906 598936
rect 559282 598924 559288 598936
rect 559243 598896 559288 598924
rect 559282 598884 559288 598896
rect 559340 598884 559346 598936
rect 291289 597567 291347 597573
rect 291289 597533 291301 597567
rect 291335 597564 291347 597567
rect 291378 597564 291384 597576
rect 291335 597536 291384 597564
rect 291335 597533 291347 597536
rect 291289 597527 291347 597533
rect 291378 597524 291384 597536
rect 291436 597524 291442 597576
rect 494054 596164 494060 596216
rect 494112 596204 494118 596216
rect 494238 596204 494244 596216
rect 494112 596176 494244 596204
rect 494112 596164 494118 596176
rect 494238 596164 494244 596176
rect 494296 596164 494302 596216
rect 3234 594804 3240 594856
rect 3292 594844 3298 594856
rect 299566 594844 299572 594856
rect 3292 594816 299572 594844
rect 3292 594804 3298 594816
rect 299566 594804 299572 594816
rect 299624 594804 299630 594856
rect 267277 592127 267335 592133
rect 267277 592093 267289 592127
rect 267323 592124 267335 592127
rect 267366 592124 267372 592136
rect 267323 592096 267372 592124
rect 267323 592093 267335 592096
rect 267277 592087 267335 592093
rect 267366 592084 267372 592096
rect 267424 592084 267430 592136
rect 235902 592016 235908 592068
rect 235960 592056 235966 592068
rect 580074 592056 580080 592068
rect 235960 592028 580080 592056
rect 235960 592016 235966 592028
rect 580074 592016 580080 592028
rect 580132 592016 580138 592068
rect 276198 591988 276204 592000
rect 276159 591960 276204 591988
rect 276198 591948 276204 591960
rect 276256 591948 276262 592000
rect 267274 589404 267280 589416
rect 267235 589376 267280 589404
rect 267274 589364 267280 589376
rect 267332 589364 267338 589416
rect 269117 589339 269175 589345
rect 269117 589305 269129 589339
rect 269163 589336 269175 589339
rect 269206 589336 269212 589348
rect 269163 589308 269212 589336
rect 269163 589305 269175 589308
rect 269117 589299 269175 589305
rect 269206 589296 269212 589308
rect 269264 589296 269270 589348
rect 299750 589336 299756 589348
rect 299711 589308 299756 589336
rect 299750 589296 299756 589308
rect 299808 589296 299814 589348
rect 559285 589339 559343 589345
rect 559285 589305 559297 589339
rect 559331 589336 559343 589339
rect 559374 589336 559380 589348
rect 559331 589308 559380 589336
rect 559331 589305 559343 589308
rect 559285 589299 559343 589305
rect 559374 589296 559380 589308
rect 559432 589296 559438 589348
rect 276198 589268 276204 589280
rect 276159 589240 276204 589268
rect 276198 589228 276204 589240
rect 276256 589228 276262 589280
rect 493870 589228 493876 589280
rect 493928 589268 493934 589280
rect 494146 589268 494152 589280
rect 493928 589240 494152 589268
rect 493928 589228 493934 589240
rect 494146 589228 494152 589240
rect 494204 589228 494210 589280
rect 269206 587840 269212 587852
rect 269167 587812 269212 587840
rect 269206 587800 269212 587812
rect 269264 587800 269270 587852
rect 559374 582468 559380 582480
rect 559300 582440 559380 582468
rect 267274 582360 267280 582412
rect 267332 582360 267338 582412
rect 269209 582403 269267 582409
rect 269209 582369 269221 582403
rect 269255 582400 269267 582403
rect 269298 582400 269304 582412
rect 269255 582372 269304 582400
rect 269255 582369 269267 582372
rect 269209 582363 269267 582369
rect 269298 582360 269304 582372
rect 269356 582360 269362 582412
rect 299750 582360 299756 582412
rect 299808 582360 299814 582412
rect 267292 582264 267320 582360
rect 267366 582264 267372 582276
rect 267292 582236 267372 582264
rect 267366 582224 267372 582236
rect 267424 582224 267430 582276
rect 276198 582264 276204 582276
rect 276159 582236 276204 582264
rect 276198 582224 276204 582236
rect 276256 582224 276262 582276
rect 299768 582264 299796 582360
rect 559300 582344 559328 582440
rect 559374 582428 559380 582440
rect 559432 582428 559438 582480
rect 559282 582292 559288 582344
rect 559340 582292 559346 582344
rect 299842 582264 299848 582276
rect 299768 582236 299848 582264
rect 299842 582224 299848 582236
rect 299900 582224 299906 582276
rect 233142 579640 233148 579692
rect 233200 579680 233206 579692
rect 580258 579680 580264 579692
rect 233200 579652 580264 579680
rect 233200 579640 233206 579652
rect 580258 579640 580264 579652
rect 580316 579640 580322 579692
rect 291378 579612 291384 579624
rect 291339 579584 291384 579612
rect 291378 579572 291384 579584
rect 291436 579572 291442 579624
rect 276014 572704 276020 572756
rect 276072 572744 276078 572756
rect 276198 572744 276204 572756
rect 276072 572716 276204 572744
rect 276072 572704 276078 572716
rect 276198 572704 276204 572716
rect 276256 572704 276262 572756
rect 287054 572704 287060 572756
rect 287112 572744 287118 572756
rect 287238 572744 287244 572756
rect 287112 572716 287244 572744
rect 287112 572704 287118 572716
rect 287238 572704 287244 572716
rect 287296 572704 287302 572756
rect 289814 572704 289820 572756
rect 289872 572744 289878 572756
rect 289998 572744 290004 572756
rect 289872 572716 290004 572744
rect 289872 572704 289878 572716
rect 289998 572704 290004 572716
rect 290056 572704 290062 572756
rect 299474 572704 299480 572756
rect 299532 572744 299538 572756
rect 299842 572744 299848 572756
rect 299532 572716 299848 572744
rect 299532 572704 299538 572716
rect 299842 572704 299848 572716
rect 299900 572704 299906 572756
rect 291381 569959 291439 569965
rect 291381 569925 291393 569959
rect 291427 569956 291439 569959
rect 291470 569956 291476 569968
rect 291427 569928 291476 569956
rect 291427 569925 291439 569928
rect 291381 569919 291439 569925
rect 291470 569916 291476 569928
rect 291528 569916 291534 569968
rect 494146 569888 494152 569900
rect 494107 569860 494152 569888
rect 494146 569848 494152 569860
rect 494204 569848 494210 569900
rect 269114 568556 269120 568608
rect 269172 568596 269178 568608
rect 269390 568596 269396 568608
rect 269172 568568 269396 568596
rect 269172 568556 269178 568568
rect 269390 568556 269396 568568
rect 269448 568556 269454 568608
rect 3418 567196 3424 567248
rect 3476 567236 3482 567248
rect 303614 567236 303620 567248
rect 3476 567208 303620 567236
rect 3476 567196 3482 567208
rect 303614 567196 303620 567208
rect 303672 567196 303678 567248
rect 269390 563156 269396 563168
rect 269316 563128 269396 563156
rect 269316 563032 269344 563128
rect 269390 563116 269396 563128
rect 269448 563116 269454 563168
rect 291470 563156 291476 563168
rect 291396 563128 291476 563156
rect 291396 563032 291424 563128
rect 291470 563116 291476 563128
rect 291528 563116 291534 563168
rect 559006 563116 559012 563168
rect 559064 563116 559070 563168
rect 494149 563091 494207 563097
rect 494149 563057 494161 563091
rect 494195 563088 494207 563091
rect 494330 563088 494336 563100
rect 494195 563060 494336 563088
rect 494195 563057 494207 563060
rect 494149 563051 494207 563057
rect 494330 563048 494336 563060
rect 494388 563048 494394 563100
rect 559024 563032 559052 563116
rect 269298 562980 269304 563032
rect 269356 562980 269362 563032
rect 291378 562980 291384 563032
rect 291436 562980 291442 563032
rect 559006 562980 559012 563032
rect 559064 562980 559070 563032
rect 267366 562912 267372 562964
rect 267424 562952 267430 562964
rect 267550 562952 267556 562964
rect 267424 562924 267556 562952
rect 267424 562912 267430 562924
rect 267550 562912 267556 562924
rect 267608 562912 267614 562964
rect 559006 560232 559012 560244
rect 558967 560204 559012 560232
rect 559006 560192 559012 560204
rect 559064 560192 559070 560244
rect 229002 556180 229008 556232
rect 229060 556220 229066 556232
rect 579890 556220 579896 556232
rect 229060 556192 579896 556220
rect 229060 556180 229066 556192
rect 579890 556180 579896 556192
rect 579948 556180 579954 556232
rect 289814 553392 289820 553444
rect 289872 553432 289878 553444
rect 289998 553432 290004 553444
rect 289872 553404 290004 553432
rect 289872 553392 289878 553404
rect 289998 553392 290004 553404
rect 290056 553392 290062 553444
rect 291286 553324 291292 553376
rect 291344 553324 291350 553376
rect 299474 553324 299480 553376
rect 299532 553364 299538 553376
rect 299934 553364 299940 553376
rect 299532 553336 299940 553364
rect 299532 553324 299538 553336
rect 299934 553324 299940 553336
rect 299992 553324 299998 553376
rect 291304 553240 291332 553324
rect 291286 553188 291292 553240
rect 291344 553188 291350 553240
rect 3142 552032 3148 552084
rect 3200 552072 3206 552084
rect 306374 552072 306380 552084
rect 3200 552044 306380 552072
rect 3200 552032 3206 552044
rect 306374 552032 306380 552044
rect 306432 552032 306438 552084
rect 276014 550604 276020 550656
rect 276072 550644 276078 550656
rect 276106 550644 276112 550656
rect 276072 550616 276112 550644
rect 276072 550604 276078 550616
rect 276106 550604 276112 550616
rect 276164 550604 276170 550656
rect 287054 550604 287060 550656
rect 287112 550644 287118 550656
rect 287146 550644 287152 550656
rect 287112 550616 287152 550644
rect 287112 550604 287118 550616
rect 287146 550604 287152 550616
rect 287204 550604 287210 550656
rect 494146 550604 494152 550656
rect 494204 550644 494210 550656
rect 494422 550644 494428 550656
rect 494204 550616 494428 550644
rect 494204 550604 494210 550616
rect 494422 550604 494428 550616
rect 494480 550604 494486 550656
rect 559009 550647 559067 550653
rect 559009 550613 559021 550647
rect 559055 550644 559067 550647
rect 559190 550644 559196 550656
rect 559055 550616 559196 550644
rect 559055 550613 559067 550616
rect 559009 550607 559067 550613
rect 559190 550604 559196 550616
rect 559248 550604 559254 550656
rect 269206 548836 269212 548888
rect 269264 548876 269270 548888
rect 269482 548876 269488 548888
rect 269264 548848 269488 548876
rect 269264 548836 269270 548848
rect 269482 548836 269488 548848
rect 269540 548836 269546 548888
rect 292574 548020 292580 548072
rect 292632 548060 292638 548072
rect 293310 548060 293316 548072
rect 292632 548032 293316 548060
rect 292632 548020 292638 548032
rect 293310 548020 293316 548032
rect 293368 548020 293374 548072
rect 231762 545096 231768 545148
rect 231820 545136 231826 545148
rect 580074 545136 580080 545148
rect 231820 545108 580080 545136
rect 231820 545096 231826 545108
rect 580074 545096 580080 545108
rect 580132 545096 580138 545148
rect 299934 543844 299940 543856
rect 299860 543816 299940 543844
rect 299860 543720 299888 543816
rect 299934 543804 299940 543816
rect 299992 543804 299998 543856
rect 494422 543844 494428 543856
rect 494348 543816 494428 543844
rect 494348 543720 494376 543816
rect 494422 543804 494428 543816
rect 494480 543804 494486 543856
rect 299842 543668 299848 543720
rect 299900 543668 299906 543720
rect 494330 543668 494336 543720
rect 494388 543668 494394 543720
rect 559006 543600 559012 543652
rect 559064 543640 559070 543652
rect 559190 543640 559196 543652
rect 559064 543612 559196 543640
rect 559064 543600 559070 543612
rect 559190 543600 559196 543612
rect 559248 543600 559254 543652
rect 287054 540880 287060 540932
rect 287112 540920 287118 540932
rect 287238 540920 287244 540932
rect 287112 540892 287244 540920
rect 287112 540880 287118 540892
rect 287238 540880 287244 540892
rect 287296 540880 287302 540932
rect 276290 539588 276296 539640
rect 276348 539628 276354 539640
rect 276382 539628 276388 539640
rect 276348 539600 276388 539628
rect 276348 539588 276354 539600
rect 276382 539588 276388 539600
rect 276440 539588 276446 539640
rect 3418 538228 3424 538280
rect 3476 538268 3482 538280
rect 304994 538268 305000 538280
rect 3476 538240 305000 538268
rect 3476 538228 3482 538240
rect 304994 538228 305000 538240
rect 305052 538228 305058 538280
rect 251818 534080 251824 534132
rect 251876 534120 251882 534132
rect 252370 534120 252376 534132
rect 251876 534092 252376 534120
rect 251876 534080 251882 534092
rect 252370 534080 252376 534092
rect 252428 534080 252434 534132
rect 287149 534123 287207 534129
rect 287149 534089 287161 534123
rect 287195 534120 287207 534123
rect 287330 534120 287336 534132
rect 287195 534092 287336 534120
rect 287195 534089 287207 534092
rect 287149 534083 287207 534089
rect 287330 534080 287336 534092
rect 287388 534080 287394 534132
rect 227622 532720 227628 532772
rect 227680 532760 227686 532772
rect 580258 532760 580264 532772
rect 227680 532732 580264 532760
rect 227680 532720 227686 532732
rect 580258 532720 580264 532732
rect 580316 532720 580322 532772
rect 267182 531292 267188 531344
rect 267240 531332 267246 531344
rect 267550 531332 267556 531344
rect 267240 531304 267556 531332
rect 267240 531292 267246 531304
rect 267550 531292 267556 531304
rect 267608 531292 267614 531344
rect 269298 531292 269304 531344
rect 269356 531332 269362 531344
rect 269574 531332 269580 531344
rect 269356 531304 269580 531332
rect 269356 531292 269362 531304
rect 269574 531292 269580 531304
rect 269632 531292 269638 531344
rect 276290 531292 276296 531344
rect 276348 531332 276354 531344
rect 276566 531332 276572 531344
rect 276348 531304 276572 531332
rect 276348 531292 276354 531304
rect 276566 531292 276572 531304
rect 276624 531292 276630 531344
rect 287146 531332 287152 531344
rect 287107 531304 287152 531332
rect 287146 531292 287152 531304
rect 287204 531292 287210 531344
rect 291286 531292 291292 531344
rect 291344 531332 291350 531344
rect 291838 531332 291844 531344
rect 291344 531304 291844 531332
rect 291344 531292 291350 531304
rect 291838 531292 291844 531304
rect 291896 531292 291902 531344
rect 293310 531292 293316 531344
rect 293368 531332 293374 531344
rect 293494 531332 293500 531344
rect 293368 531304 293500 531332
rect 293368 531292 293374 531304
rect 293494 531292 293500 531304
rect 293552 531292 293558 531344
rect 299658 531292 299664 531344
rect 299716 531332 299722 531344
rect 299934 531332 299940 531344
rect 299716 531304 299940 531332
rect 299716 531292 299722 531304
rect 299934 531292 299940 531304
rect 299992 531292 299998 531344
rect 494146 531292 494152 531344
rect 494204 531332 494210 531344
rect 494422 531332 494428 531344
rect 494204 531304 494428 531332
rect 494204 531292 494210 531304
rect 494422 531292 494428 531304
rect 494480 531292 494486 531344
rect 230474 526464 230480 526516
rect 230532 526504 230538 526516
rect 231762 526504 231768 526516
rect 230532 526476 231768 526504
rect 230532 526464 230538 526476
rect 231762 526464 231768 526476
rect 231820 526464 231826 526516
rect 231854 526464 231860 526516
rect 231912 526504 231918 526516
rect 233142 526504 233148 526516
rect 231912 526476 233148 526504
rect 231912 526464 231918 526476
rect 233142 526464 233148 526476
rect 233200 526464 233206 526516
rect 233234 526464 233240 526516
rect 233292 526504 233298 526516
rect 234522 526504 234528 526516
rect 233292 526476 234528 526504
rect 233292 526464 233298 526476
rect 234522 526464 234528 526476
rect 234580 526464 234586 526516
rect 234614 526464 234620 526516
rect 234672 526504 234678 526516
rect 235902 526504 235908 526516
rect 234672 526476 235908 526504
rect 234672 526464 234678 526476
rect 235902 526464 235908 526476
rect 235960 526464 235966 526516
rect 237374 526464 237380 526516
rect 237432 526504 237438 526516
rect 238662 526504 238668 526516
rect 237432 526476 238668 526504
rect 237432 526464 237438 526476
rect 238662 526464 238668 526476
rect 238720 526464 238726 526516
rect 276382 526328 276388 526380
rect 276440 526368 276446 526380
rect 276566 526368 276572 526380
rect 276440 526340 276572 526368
rect 276440 526328 276446 526340
rect 276566 526328 276572 526340
rect 276624 526328 276630 526380
rect 263318 523880 263324 523932
rect 263376 523920 263382 523932
rect 279418 523920 279424 523932
rect 263376 523892 279424 523920
rect 263376 523880 263382 523892
rect 279418 523880 279424 523892
rect 279476 523880 279482 523932
rect 268562 523812 268568 523864
rect 268620 523852 268626 523864
rect 299934 523852 299940 523864
rect 268620 523824 299940 523852
rect 268620 523812 268626 523824
rect 299934 523812 299940 523824
rect 299992 523812 299998 523864
rect 253106 523744 253112 523796
rect 253164 523784 253170 523796
rect 494422 523784 494428 523796
rect 253164 523756 494428 523784
rect 253164 523744 253170 523756
rect 494422 523744 494428 523756
rect 494480 523744 494486 523796
rect 248138 523676 248144 523728
rect 248196 523716 248202 523728
rect 559190 523716 559196 523728
rect 248196 523688 559196 523716
rect 248196 523676 248202 523688
rect 559190 523676 559196 523688
rect 559248 523676 559254 523728
rect 219066 522928 219072 522980
rect 219124 522968 219130 522980
rect 371050 522968 371056 522980
rect 219124 522940 371056 522968
rect 219124 522928 219130 522940
rect 371050 522928 371056 522940
rect 371108 522928 371114 522980
rect 213822 522860 213828 522912
rect 213880 522900 213886 522912
rect 370774 522900 370780 522912
rect 213880 522872 370780 522900
rect 213880 522860 213886 522872
rect 370774 522860 370780 522872
rect 370832 522860 370838 522912
rect 189994 522792 190000 522844
rect 190052 522832 190058 522844
rect 376018 522832 376024 522844
rect 190052 522804 376024 522832
rect 190052 522792 190058 522804
rect 376018 522792 376024 522804
rect 376076 522792 376082 522844
rect 2958 522724 2964 522776
rect 3016 522764 3022 522776
rect 309134 522764 309140 522776
rect 3016 522736 309140 522764
rect 3016 522724 3022 522736
rect 309134 522724 309140 522736
rect 309192 522724 309198 522776
rect 4706 522656 4712 522708
rect 4764 522696 4770 522708
rect 312446 522696 312452 522708
rect 4764 522668 312452 522696
rect 4764 522656 4770 522668
rect 312446 522656 312452 522668
rect 312504 522656 312510 522708
rect 3050 522588 3056 522640
rect 3108 522628 3114 522640
rect 310606 522628 310612 522640
rect 3108 522600 310612 522628
rect 3108 522588 3114 522600
rect 310606 522588 310612 522600
rect 310664 522588 310670 522640
rect 3142 522520 3148 522572
rect 3200 522560 3206 522572
rect 317414 522560 317420 522572
rect 3200 522532 317420 522560
rect 3200 522520 3206 522532
rect 317414 522520 317420 522532
rect 317472 522520 317478 522572
rect 3234 522452 3240 522504
rect 3292 522492 3298 522504
rect 319254 522492 319260 522504
rect 3292 522464 319260 522492
rect 3292 522452 3298 522464
rect 319254 522452 319260 522464
rect 319312 522452 319318 522504
rect 5442 522384 5448 522436
rect 5500 522424 5506 522436
rect 323026 522424 323032 522436
rect 5500 522396 323032 522424
rect 5500 522384 5506 522396
rect 323026 522384 323032 522396
rect 323084 522384 323090 522436
rect 325694 522384 325700 522436
rect 325752 522424 325758 522436
rect 335262 522424 335268 522436
rect 325752 522396 335268 522424
rect 325752 522384 325758 522396
rect 335262 522384 335268 522396
rect 335320 522384 335326 522436
rect 6178 522316 6184 522368
rect 6236 522356 6242 522368
rect 327718 522356 327724 522368
rect 6236 522328 327724 522356
rect 6236 522316 6242 522328
rect 327718 522316 327724 522328
rect 327776 522316 327782 522368
rect 4062 522248 4068 522300
rect 4120 522288 4126 522300
rect 326062 522288 326068 522300
rect 4120 522260 326068 522288
rect 4120 522248 4126 522260
rect 326062 522248 326068 522260
rect 326120 522248 326126 522300
rect 19978 522180 19984 522232
rect 20036 522220 20042 522232
rect 343174 522220 343180 522232
rect 20036 522192 343180 522220
rect 20036 522180 20042 522192
rect 343174 522180 343180 522192
rect 343232 522180 343238 522232
rect 345014 522180 345020 522232
rect 345072 522220 345078 522232
rect 354582 522220 354588 522232
rect 345072 522192 354588 522220
rect 345072 522180 345078 522192
rect 354582 522180 354588 522192
rect 354640 522180 354646 522232
rect 10318 522112 10324 522164
rect 10376 522152 10382 522164
rect 332870 522152 332876 522164
rect 10376 522124 332876 522152
rect 10376 522112 10382 522124
rect 332870 522112 332876 522124
rect 332928 522112 332934 522164
rect 13078 522044 13084 522096
rect 13136 522084 13142 522096
rect 338114 522084 338120 522096
rect 13136 522056 338120 522084
rect 13136 522044 13142 522056
rect 338114 522044 338120 522056
rect 338172 522044 338178 522096
rect 5258 521976 5264 522028
rect 5316 522016 5322 522028
rect 331214 522016 331220 522028
rect 5316 521988 331220 522016
rect 5316 521976 5322 521988
rect 331214 521976 331220 521988
rect 331272 521976 331278 522028
rect 21358 521908 21364 521960
rect 21416 521948 21422 521960
rect 348326 521948 348332 521960
rect 21416 521920 348332 521948
rect 21416 521908 21422 521920
rect 348326 521908 348332 521920
rect 348384 521908 348390 521960
rect 3878 521840 3884 521892
rect 3936 521880 3942 521892
rect 334526 521880 334532 521892
rect 3936 521852 334532 521880
rect 3936 521840 3942 521852
rect 334526 521840 334532 521852
rect 334584 521840 334590 521892
rect 3786 521772 3792 521824
rect 3844 521812 3850 521824
rect 336366 521812 336372 521824
rect 3844 521784 336372 521812
rect 3844 521772 3850 521784
rect 336366 521772 336372 521784
rect 336424 521772 336430 521824
rect 5074 521704 5080 521756
rect 5132 521744 5138 521756
rect 346486 521744 346492 521756
rect 5132 521716 346492 521744
rect 5132 521704 5138 521716
rect 346486 521704 346492 521716
rect 346544 521704 346550 521756
rect 186130 521636 186136 521688
rect 186188 521676 186194 521688
rect 276201 521679 276259 521685
rect 276201 521676 276213 521679
rect 186188 521648 276213 521676
rect 186188 521636 186194 521648
rect 276201 521645 276213 521648
rect 276247 521645 276259 521679
rect 276201 521639 276259 521645
rect 276477 521679 276535 521685
rect 276477 521645 276489 521679
rect 276523 521676 276535 521679
rect 287057 521679 287115 521685
rect 287057 521676 287069 521679
rect 276523 521648 287069 521676
rect 276523 521645 276535 521648
rect 276477 521639 276535 521645
rect 287057 521645 287069 521648
rect 287103 521645 287115 521679
rect 287057 521639 287115 521645
rect 287333 521679 287391 521685
rect 287333 521645 287345 521679
rect 287379 521676 287391 521679
rect 580718 521676 580724 521688
rect 287379 521648 580724 521676
rect 287379 521645 287391 521648
rect 287333 521639 287391 521645
rect 580718 521636 580724 521648
rect 580776 521636 580782 521688
rect 311802 521568 311808 521620
rect 311860 521608 311866 521620
rect 311986 521608 311992 521620
rect 311860 521580 311992 521608
rect 311860 521568 311866 521580
rect 311986 521568 311992 521580
rect 312044 521568 312050 521620
rect 224218 520820 224224 520872
rect 224276 520860 224282 520872
rect 369762 520860 369768 520872
rect 224276 520832 369768 520860
rect 224276 520820 224282 520832
rect 369762 520820 369768 520832
rect 369820 520820 369826 520872
rect 220722 520752 220728 520804
rect 220780 520792 220786 520804
rect 370958 520792 370964 520804
rect 220780 520764 370964 520792
rect 220780 520752 220786 520764
rect 370958 520752 370964 520764
rect 371016 520752 371022 520804
rect 217226 520684 217232 520736
rect 217284 520724 217290 520736
rect 370866 520724 370872 520736
rect 217284 520696 370872 520724
rect 217284 520684 217290 520696
rect 370866 520684 370872 520696
rect 370924 520684 370930 520736
rect 212074 520616 212080 520668
rect 212132 520656 212138 520668
rect 370590 520656 370596 520668
rect 212132 520628 370596 520656
rect 212132 520616 212138 520628
rect 370590 520616 370596 520628
rect 370648 520616 370654 520668
rect 208762 520548 208768 520600
rect 208820 520588 208826 520600
rect 369670 520588 369676 520600
rect 208820 520560 369676 520588
rect 208820 520548 208826 520560
rect 369670 520548 369676 520560
rect 369728 520548 369734 520600
rect 206922 520480 206928 520532
rect 206980 520520 206986 520532
rect 369578 520520 369584 520532
rect 206980 520492 369584 520520
rect 206980 520480 206986 520492
rect 369578 520480 369584 520492
rect 369636 520480 369642 520532
rect 203610 520412 203616 520464
rect 203668 520452 203674 520464
rect 369486 520452 369492 520464
rect 203668 520424 369492 520452
rect 203668 520412 203674 520424
rect 369486 520412 369492 520424
rect 369544 520412 369550 520464
rect 188154 520344 188160 520396
rect 188212 520384 188218 520396
rect 580902 520384 580908 520396
rect 188212 520356 580908 520384
rect 188212 520344 188218 520356
rect 580902 520344 580908 520356
rect 580960 520344 580966 520396
rect 183186 520276 183192 520328
rect 183244 520316 183250 520328
rect 580534 520316 580540 520328
rect 183244 520288 580540 520316
rect 183244 520276 183250 520288
rect 580534 520276 580540 520288
rect 580592 520276 580598 520328
rect 171873 519775 171931 519781
rect 171873 519741 171885 519775
rect 171919 519772 171931 519775
rect 181533 519775 181591 519781
rect 181533 519772 181545 519775
rect 171919 519744 181545 519772
rect 171919 519741 171931 519744
rect 171873 519735 171931 519741
rect 181533 519741 181545 519744
rect 181579 519741 181591 519775
rect 181533 519735 181591 519741
rect 209961 519775 210019 519781
rect 209961 519741 209973 519775
rect 210007 519772 210019 519775
rect 219161 519775 219219 519781
rect 219161 519772 219173 519775
rect 210007 519744 219173 519772
rect 210007 519741 210019 519744
rect 209961 519735 210019 519741
rect 219161 519741 219173 519744
rect 219207 519741 219219 519775
rect 219161 519735 219219 519741
rect 17313 519707 17371 519713
rect 17313 519673 17325 519707
rect 17359 519704 17371 519707
rect 26789 519707 26847 519713
rect 26789 519704 26801 519707
rect 17359 519676 26801 519704
rect 17359 519673 17371 519676
rect 17313 519667 17371 519673
rect 26789 519673 26801 519676
rect 26835 519673 26847 519707
rect 26789 519667 26847 519673
rect 36633 519707 36691 519713
rect 36633 519673 36645 519707
rect 36679 519704 36691 519707
rect 46109 519707 46167 519713
rect 46109 519704 46121 519707
rect 36679 519676 46121 519704
rect 36679 519673 36691 519676
rect 36633 519667 36691 519673
rect 46109 519673 46121 519676
rect 46155 519673 46167 519707
rect 46109 519667 46167 519673
rect 55953 519707 56011 519713
rect 55953 519673 55965 519707
rect 55999 519704 56011 519707
rect 65429 519707 65487 519713
rect 65429 519704 65441 519707
rect 55999 519676 65441 519704
rect 55999 519673 56011 519676
rect 55953 519667 56011 519673
rect 65429 519673 65441 519676
rect 65475 519673 65487 519707
rect 65429 519667 65487 519673
rect 75273 519707 75331 519713
rect 75273 519673 75285 519707
rect 75319 519704 75331 519707
rect 84749 519707 84807 519713
rect 84749 519704 84761 519707
rect 75319 519676 84761 519704
rect 75319 519673 75331 519676
rect 75273 519667 75331 519673
rect 84749 519673 84761 519676
rect 84795 519673 84807 519707
rect 84749 519667 84807 519673
rect 94593 519707 94651 519713
rect 94593 519673 94605 519707
rect 94639 519704 94651 519707
rect 104069 519707 104127 519713
rect 104069 519704 104081 519707
rect 94639 519676 104081 519704
rect 94639 519673 94651 519676
rect 94593 519667 94651 519673
rect 104069 519673 104081 519676
rect 104115 519673 104127 519707
rect 104069 519667 104127 519673
rect 113913 519707 113971 519713
rect 113913 519673 113925 519707
rect 113959 519704 113971 519707
rect 123389 519707 123447 519713
rect 123389 519704 123401 519707
rect 113959 519676 123401 519704
rect 113959 519673 113971 519676
rect 113913 519667 113971 519673
rect 123389 519673 123401 519676
rect 123435 519673 123447 519707
rect 123389 519667 123447 519673
rect 133233 519707 133291 519713
rect 133233 519673 133245 519707
rect 133279 519704 133291 519707
rect 142709 519707 142767 519713
rect 142709 519704 142721 519707
rect 133279 519676 142721 519704
rect 133279 519673 133291 519676
rect 133233 519667 133291 519673
rect 142709 519673 142721 519676
rect 142755 519673 142767 519707
rect 142709 519667 142767 519673
rect 152553 519707 152611 519713
rect 152553 519673 152565 519707
rect 152599 519704 152611 519707
rect 162029 519707 162087 519713
rect 162029 519704 162041 519707
rect 152599 519676 162041 519704
rect 152599 519673 152611 519676
rect 152553 519667 152611 519673
rect 162029 519673 162041 519676
rect 162075 519673 162087 519707
rect 162029 519667 162087 519673
rect 171689 519707 171747 519713
rect 171689 519673 171701 519707
rect 171735 519704 171747 519707
rect 181349 519707 181407 519713
rect 181349 519704 181361 519707
rect 171735 519676 181361 519704
rect 171735 519673 171747 519676
rect 171689 519667 171747 519673
rect 181349 519673 181361 519676
rect 181395 519673 181407 519707
rect 181349 519667 181407 519673
rect 188341 519707 188399 519713
rect 188341 519673 188353 519707
rect 188387 519704 188399 519707
rect 200669 519707 200727 519713
rect 200669 519704 200681 519707
rect 188387 519676 200681 519704
rect 188387 519673 188399 519676
rect 188341 519667 188399 519673
rect 200669 519673 200681 519676
rect 200715 519673 200727 519707
rect 200669 519667 200727 519673
rect 209869 519707 209927 519713
rect 209869 519673 209881 519707
rect 209915 519704 209927 519707
rect 219253 519707 219311 519713
rect 219253 519704 219265 519707
rect 209915 519676 219265 519704
rect 209915 519673 209927 519676
rect 209869 519667 209927 519673
rect 219253 519673 219265 519676
rect 219299 519673 219311 519707
rect 219253 519667 219311 519673
rect 17129 519639 17187 519645
rect 17129 519605 17141 519639
rect 17175 519636 17187 519639
rect 26881 519639 26939 519645
rect 26881 519636 26893 519639
rect 17175 519608 26893 519636
rect 17175 519605 17187 519608
rect 17129 519599 17187 519605
rect 26881 519605 26893 519608
rect 26927 519605 26939 519639
rect 26881 519599 26939 519605
rect 36449 519639 36507 519645
rect 36449 519605 36461 519639
rect 36495 519636 36507 519639
rect 46201 519639 46259 519645
rect 46201 519636 46213 519639
rect 36495 519608 46213 519636
rect 36495 519605 36507 519608
rect 36449 519599 36507 519605
rect 46201 519605 46213 519608
rect 46247 519605 46259 519639
rect 46201 519599 46259 519605
rect 55769 519639 55827 519645
rect 55769 519605 55781 519639
rect 55815 519636 55827 519639
rect 65521 519639 65579 519645
rect 65521 519636 65533 519639
rect 55815 519608 65533 519636
rect 55815 519605 55827 519608
rect 55769 519599 55827 519605
rect 65521 519605 65533 519608
rect 65567 519605 65579 519639
rect 65521 519599 65579 519605
rect 75089 519639 75147 519645
rect 75089 519605 75101 519639
rect 75135 519636 75147 519639
rect 84841 519639 84899 519645
rect 84841 519636 84853 519639
rect 75135 519608 84853 519636
rect 75135 519605 75147 519608
rect 75089 519599 75147 519605
rect 84841 519605 84853 519608
rect 84887 519605 84899 519639
rect 84841 519599 84899 519605
rect 94409 519639 94467 519645
rect 94409 519605 94421 519639
rect 94455 519636 94467 519639
rect 104161 519639 104219 519645
rect 104161 519636 104173 519639
rect 94455 519608 104173 519636
rect 94455 519605 94467 519608
rect 94409 519599 94467 519605
rect 104161 519605 104173 519608
rect 104207 519605 104219 519639
rect 104161 519599 104219 519605
rect 113729 519639 113787 519645
rect 113729 519605 113741 519639
rect 113775 519636 113787 519639
rect 123481 519639 123539 519645
rect 123481 519636 123493 519639
rect 113775 519608 123493 519636
rect 113775 519605 113787 519608
rect 113729 519599 113787 519605
rect 123481 519605 123493 519608
rect 123527 519605 123539 519639
rect 123481 519599 123539 519605
rect 133049 519639 133107 519645
rect 133049 519605 133061 519639
rect 133095 519636 133107 519639
rect 142801 519639 142859 519645
rect 142801 519636 142813 519639
rect 133095 519608 142813 519636
rect 133095 519605 133107 519608
rect 133049 519599 133107 519605
rect 142801 519605 142813 519608
rect 142847 519605 142859 519639
rect 142801 519599 142859 519605
rect 152369 519639 152427 519645
rect 152369 519605 152381 519639
rect 152415 519636 152427 519639
rect 162121 519639 162179 519645
rect 162121 519636 162133 519639
rect 152415 519608 162133 519636
rect 152415 519605 152427 519608
rect 152369 519599 152427 519605
rect 162121 519605 162133 519608
rect 162167 519605 162179 519639
rect 162121 519599 162179 519605
rect 171781 519639 171839 519645
rect 171781 519605 171793 519639
rect 171827 519636 171839 519639
rect 181441 519639 181499 519645
rect 181441 519636 181453 519639
rect 171827 519608 181453 519636
rect 171827 519605 171839 519608
rect 171781 519599 171839 519605
rect 181441 519605 181453 519608
rect 181487 519605 181499 519639
rect 181441 519599 181499 519605
rect 191101 519639 191159 519645
rect 191101 519605 191113 519639
rect 191147 519636 191159 519639
rect 200761 519639 200819 519645
rect 200761 519636 200773 519639
rect 191147 519608 200773 519636
rect 191147 519605 191159 519608
rect 191101 519599 191159 519605
rect 200761 519605 200773 519608
rect 200807 519605 200819 519639
rect 200761 519599 200819 519605
rect 209777 519639 209835 519645
rect 209777 519605 209789 519639
rect 209823 519636 209835 519639
rect 219345 519639 219403 519645
rect 219345 519636 219357 519639
rect 209823 519608 219357 519636
rect 209823 519605 209835 519608
rect 209777 519599 209835 519605
rect 219345 519605 219357 519608
rect 219391 519605 219403 519639
rect 219345 519599 219403 519605
rect 305365 519639 305423 519645
rect 305365 519605 305377 519639
rect 305411 519636 305423 519639
rect 316865 519639 316923 519645
rect 316865 519636 316877 519639
rect 305411 519608 316877 519636
rect 305411 519605 305423 519608
rect 305365 519599 305423 519605
rect 316865 519605 316877 519608
rect 316911 519605 316923 519639
rect 316865 519599 316923 519605
rect 17221 519571 17279 519577
rect 17221 519537 17233 519571
rect 17267 519568 17279 519571
rect 22741 519571 22799 519577
rect 22741 519568 22753 519571
rect 17267 519540 22753 519568
rect 17267 519537 17279 519540
rect 17221 519531 17279 519537
rect 22741 519537 22753 519540
rect 22787 519537 22799 519571
rect 22741 519531 22799 519537
rect 36541 519571 36599 519577
rect 36541 519537 36553 519571
rect 36587 519568 36599 519571
rect 42061 519571 42119 519577
rect 42061 519568 42073 519571
rect 36587 519540 42073 519568
rect 36587 519537 36599 519540
rect 36541 519531 36599 519537
rect 42061 519537 42073 519540
rect 42107 519537 42119 519571
rect 42061 519531 42119 519537
rect 55861 519571 55919 519577
rect 55861 519537 55873 519571
rect 55907 519568 55919 519571
rect 61381 519571 61439 519577
rect 61381 519568 61393 519571
rect 55907 519540 61393 519568
rect 55907 519537 55919 519540
rect 55861 519531 55919 519537
rect 61381 519537 61393 519540
rect 61427 519537 61439 519571
rect 61381 519531 61439 519537
rect 75181 519571 75239 519577
rect 75181 519537 75193 519571
rect 75227 519568 75239 519571
rect 80701 519571 80759 519577
rect 80701 519568 80713 519571
rect 75227 519540 80713 519568
rect 75227 519537 75239 519540
rect 75181 519531 75239 519537
rect 80701 519537 80713 519540
rect 80747 519537 80759 519571
rect 80701 519531 80759 519537
rect 94501 519571 94559 519577
rect 94501 519537 94513 519571
rect 94547 519568 94559 519571
rect 100021 519571 100079 519577
rect 100021 519568 100033 519571
rect 94547 519540 100033 519568
rect 94547 519537 94559 519540
rect 94501 519531 94559 519537
rect 100021 519537 100033 519540
rect 100067 519537 100079 519571
rect 100021 519531 100079 519537
rect 113821 519571 113879 519577
rect 113821 519537 113833 519571
rect 113867 519568 113879 519571
rect 119341 519571 119399 519577
rect 119341 519568 119353 519571
rect 113867 519540 119353 519568
rect 113867 519537 113879 519540
rect 113821 519531 113879 519537
rect 119341 519537 119353 519540
rect 119387 519537 119399 519571
rect 119341 519531 119399 519537
rect 133141 519571 133199 519577
rect 133141 519537 133153 519571
rect 133187 519568 133199 519571
rect 138661 519571 138719 519577
rect 138661 519568 138673 519571
rect 133187 519540 138673 519568
rect 133187 519537 133199 519540
rect 133141 519531 133199 519537
rect 138661 519537 138673 519540
rect 138707 519537 138719 519571
rect 138661 519531 138719 519537
rect 152461 519571 152519 519577
rect 152461 519537 152473 519571
rect 152507 519568 152519 519571
rect 157981 519571 158039 519577
rect 157981 519568 157993 519571
rect 152507 519540 157993 519568
rect 152507 519537 152519 519540
rect 152461 519531 152519 519537
rect 157981 519537 157993 519540
rect 158027 519537 158039 519571
rect 179414 519568 179420 519580
rect 179375 519540 179420 519568
rect 157981 519531 158039 519537
rect 179414 519528 179420 519540
rect 179472 519528 179478 519580
rect 189997 519571 190055 519577
rect 189997 519537 190009 519571
rect 190043 519568 190055 519571
rect 195977 519571 196035 519577
rect 195977 519568 195989 519571
rect 190043 519540 195989 519568
rect 190043 519537 190055 519540
rect 189997 519531 190055 519537
rect 195977 519537 195989 519540
rect 196023 519537 196035 519571
rect 195977 519531 196035 519537
rect 215570 519528 215576 519580
rect 215628 519568 215634 519580
rect 370682 519568 370688 519580
rect 215628 519540 370688 519568
rect 215628 519528 215634 519540
rect 370682 519528 370688 519540
rect 370740 519528 370746 519580
rect 6362 519460 6368 519512
rect 6420 519500 6426 519512
rect 314102 519500 314108 519512
rect 6420 519472 314108 519500
rect 6420 519460 6426 519472
rect 314102 519460 314108 519472
rect 314160 519460 314166 519512
rect 325881 519503 325939 519509
rect 325881 519469 325893 519503
rect 325927 519500 325939 519503
rect 335173 519503 335231 519509
rect 335173 519500 335185 519503
rect 325927 519472 335185 519500
rect 325927 519469 325939 519472
rect 325881 519463 325939 519469
rect 335173 519469 335185 519472
rect 335219 519469 335231 519503
rect 335173 519463 335231 519469
rect 5350 519392 5356 519444
rect 5408 519432 5414 519444
rect 320910 519432 320916 519444
rect 5408 519404 320916 519432
rect 5408 519392 5414 519404
rect 320910 519392 320916 519404
rect 320968 519392 320974 519444
rect 325789 519435 325847 519441
rect 325789 519401 325801 519435
rect 325835 519432 325847 519435
rect 335265 519435 335323 519441
rect 335265 519432 335277 519435
rect 325835 519404 335277 519432
rect 325835 519401 325847 519404
rect 325789 519395 325847 519401
rect 335265 519401 335277 519404
rect 335311 519401 335323 519435
rect 335265 519395 335323 519401
rect 3326 519324 3332 519376
rect 3384 519364 3390 519376
rect 324406 519364 324412 519376
rect 3384 519336 324412 519364
rect 3384 519324 3390 519336
rect 324406 519324 324412 519336
rect 324464 519324 324470 519376
rect 325697 519367 325755 519373
rect 325697 519333 325709 519367
rect 325743 519364 325755 519367
rect 339678 519364 339684 519376
rect 325743 519336 339684 519364
rect 325743 519333 325755 519336
rect 325697 519327 325755 519333
rect 339678 519324 339684 519336
rect 339736 519324 339742 519376
rect 3970 519256 3976 519308
rect 4028 519296 4034 519308
rect 329650 519296 329656 519308
rect 4028 519268 329656 519296
rect 4028 519256 4034 519268
rect 329650 519256 329656 519268
rect 329708 519256 329714 519308
rect 345014 519256 345020 519308
rect 345072 519256 345078 519308
rect 349982 519296 349988 519308
rect 349943 519268 349988 519296
rect 349982 519256 349988 519268
rect 350040 519256 350046 519308
rect 351822 519296 351828 519308
rect 351783 519268 351828 519296
rect 351822 519256 351828 519268
rect 351880 519256 351886 519308
rect 355134 519296 355140 519308
rect 355095 519268 355140 519296
rect 355134 519256 355140 519268
rect 355192 519256 355198 519308
rect 360286 519296 360292 519308
rect 355244 519268 360292 519296
rect 3694 519188 3700 519240
rect 3752 519228 3758 519240
rect 17221 519231 17279 519237
rect 17221 519228 17233 519231
rect 3752 519200 17233 519228
rect 3752 519188 3758 519200
rect 17221 519197 17233 519200
rect 17267 519197 17279 519231
rect 17221 519191 17279 519197
rect 22741 519231 22799 519237
rect 22741 519197 22753 519231
rect 22787 519228 22799 519231
rect 36541 519231 36599 519237
rect 36541 519228 36553 519231
rect 22787 519200 36553 519228
rect 22787 519197 22799 519200
rect 22741 519191 22799 519197
rect 36541 519197 36553 519200
rect 36587 519197 36599 519231
rect 36541 519191 36599 519197
rect 42061 519231 42119 519237
rect 42061 519197 42073 519231
rect 42107 519228 42119 519231
rect 55861 519231 55919 519237
rect 55861 519228 55873 519231
rect 42107 519200 55873 519228
rect 42107 519197 42119 519200
rect 42061 519191 42119 519197
rect 55861 519197 55873 519200
rect 55907 519197 55919 519231
rect 55861 519191 55919 519197
rect 61381 519231 61439 519237
rect 61381 519197 61393 519231
rect 61427 519228 61439 519231
rect 75181 519231 75239 519237
rect 75181 519228 75193 519231
rect 61427 519200 75193 519228
rect 61427 519197 61439 519200
rect 61381 519191 61439 519197
rect 75181 519197 75193 519200
rect 75227 519197 75239 519231
rect 75181 519191 75239 519197
rect 80701 519231 80759 519237
rect 80701 519197 80713 519231
rect 80747 519228 80759 519231
rect 94501 519231 94559 519237
rect 94501 519228 94513 519231
rect 80747 519200 94513 519228
rect 80747 519197 80759 519200
rect 80701 519191 80759 519197
rect 94501 519197 94513 519200
rect 94547 519197 94559 519231
rect 94501 519191 94559 519197
rect 100021 519231 100079 519237
rect 100021 519197 100033 519231
rect 100067 519228 100079 519231
rect 113821 519231 113879 519237
rect 113821 519228 113833 519231
rect 100067 519200 113833 519228
rect 100067 519197 100079 519200
rect 100021 519191 100079 519197
rect 113821 519197 113833 519200
rect 113867 519197 113879 519231
rect 113821 519191 113879 519197
rect 119341 519231 119399 519237
rect 119341 519197 119353 519231
rect 119387 519228 119399 519231
rect 133141 519231 133199 519237
rect 133141 519228 133153 519231
rect 119387 519200 133153 519228
rect 119387 519197 119399 519200
rect 119341 519191 119399 519197
rect 133141 519197 133153 519200
rect 133187 519197 133199 519231
rect 133141 519191 133199 519197
rect 138661 519231 138719 519237
rect 138661 519197 138673 519231
rect 138707 519228 138719 519231
rect 152461 519231 152519 519237
rect 152461 519228 152473 519231
rect 138707 519200 152473 519228
rect 138707 519197 138719 519200
rect 138661 519191 138719 519197
rect 152461 519197 152473 519200
rect 152507 519197 152519 519231
rect 152461 519191 152519 519197
rect 157981 519231 158039 519237
rect 157981 519197 157993 519231
rect 158027 519228 158039 519231
rect 171781 519231 171839 519237
rect 171781 519228 171793 519231
rect 158027 519200 171793 519228
rect 158027 519197 158039 519200
rect 157981 519191 158039 519197
rect 171781 519197 171793 519200
rect 171827 519197 171839 519231
rect 171781 519191 171839 519197
rect 181441 519231 181499 519237
rect 181441 519197 181453 519231
rect 181487 519228 181499 519231
rect 189997 519231 190055 519237
rect 189997 519228 190009 519231
rect 181487 519200 190009 519228
rect 181487 519197 181499 519200
rect 181441 519191 181499 519197
rect 189997 519197 190009 519200
rect 190043 519197 190055 519231
rect 189997 519191 190055 519197
rect 195977 519231 196035 519237
rect 195977 519197 195989 519231
rect 196023 519228 196035 519231
rect 209777 519231 209835 519237
rect 209777 519228 209789 519231
rect 196023 519200 209789 519228
rect 196023 519197 196035 519200
rect 195977 519191 196035 519197
rect 209777 519197 209789 519200
rect 209823 519197 209835 519231
rect 209777 519191 209835 519197
rect 219345 519231 219403 519237
rect 219345 519197 219357 519231
rect 219391 519228 219403 519231
rect 305365 519231 305423 519237
rect 305365 519228 305377 519231
rect 219391 519200 305377 519228
rect 219391 519197 219403 519200
rect 219345 519191 219403 519197
rect 305365 519197 305377 519200
rect 305411 519197 305423 519231
rect 316773 519231 316831 519237
rect 316773 519228 316785 519231
rect 305365 519191 305423 519197
rect 306944 519200 316785 519228
rect 5166 519120 5172 519172
rect 5224 519160 5230 519172
rect 306837 519163 306895 519169
rect 306837 519160 306849 519163
rect 5224 519132 306849 519160
rect 5224 519120 5230 519132
rect 306837 519129 306849 519132
rect 306883 519129 306895 519163
rect 306837 519123 306895 519129
rect 4982 519052 4988 519104
rect 5040 519092 5046 519104
rect 17129 519095 17187 519101
rect 17129 519092 17141 519095
rect 5040 519064 17141 519092
rect 5040 519052 5046 519064
rect 17129 519061 17141 519064
rect 17175 519061 17187 519095
rect 17129 519055 17187 519061
rect 26881 519095 26939 519101
rect 26881 519061 26893 519095
rect 26927 519092 26939 519095
rect 36449 519095 36507 519101
rect 36449 519092 36461 519095
rect 26927 519064 36461 519092
rect 26927 519061 26939 519064
rect 26881 519055 26939 519061
rect 36449 519061 36461 519064
rect 36495 519061 36507 519095
rect 36449 519055 36507 519061
rect 46201 519095 46259 519101
rect 46201 519061 46213 519095
rect 46247 519092 46259 519095
rect 55769 519095 55827 519101
rect 55769 519092 55781 519095
rect 46247 519064 55781 519092
rect 46247 519061 46259 519064
rect 46201 519055 46259 519061
rect 55769 519061 55781 519064
rect 55815 519061 55827 519095
rect 55769 519055 55827 519061
rect 65521 519095 65579 519101
rect 65521 519061 65533 519095
rect 65567 519092 65579 519095
rect 75089 519095 75147 519101
rect 75089 519092 75101 519095
rect 65567 519064 75101 519092
rect 65567 519061 65579 519064
rect 65521 519055 65579 519061
rect 75089 519061 75101 519064
rect 75135 519061 75147 519095
rect 75089 519055 75147 519061
rect 84841 519095 84899 519101
rect 84841 519061 84853 519095
rect 84887 519092 84899 519095
rect 94409 519095 94467 519101
rect 94409 519092 94421 519095
rect 84887 519064 94421 519092
rect 84887 519061 84899 519064
rect 84841 519055 84899 519061
rect 94409 519061 94421 519064
rect 94455 519061 94467 519095
rect 94409 519055 94467 519061
rect 104161 519095 104219 519101
rect 104161 519061 104173 519095
rect 104207 519092 104219 519095
rect 113729 519095 113787 519101
rect 113729 519092 113741 519095
rect 104207 519064 113741 519092
rect 104207 519061 104219 519064
rect 104161 519055 104219 519061
rect 113729 519061 113741 519064
rect 113775 519061 113787 519095
rect 113729 519055 113787 519061
rect 123481 519095 123539 519101
rect 123481 519061 123493 519095
rect 123527 519092 123539 519095
rect 133049 519095 133107 519101
rect 133049 519092 133061 519095
rect 123527 519064 133061 519092
rect 123527 519061 123539 519064
rect 123481 519055 123539 519061
rect 133049 519061 133061 519064
rect 133095 519061 133107 519095
rect 133049 519055 133107 519061
rect 142801 519095 142859 519101
rect 142801 519061 142813 519095
rect 142847 519092 142859 519095
rect 152369 519095 152427 519101
rect 152369 519092 152381 519095
rect 142847 519064 152381 519092
rect 142847 519061 142859 519064
rect 142801 519055 142859 519061
rect 152369 519061 152381 519064
rect 152415 519061 152427 519095
rect 152369 519055 152427 519061
rect 162121 519095 162179 519101
rect 162121 519061 162133 519095
rect 162167 519092 162179 519095
rect 171689 519095 171747 519101
rect 171689 519092 171701 519095
rect 162167 519064 171701 519092
rect 162167 519061 162179 519064
rect 162121 519055 162179 519061
rect 171689 519061 171701 519064
rect 171735 519061 171747 519095
rect 171689 519055 171747 519061
rect 181349 519095 181407 519101
rect 181349 519061 181361 519095
rect 181395 519092 181407 519095
rect 191101 519095 191159 519101
rect 191101 519092 191113 519095
rect 181395 519064 191113 519092
rect 181395 519061 181407 519064
rect 181349 519055 181407 519061
rect 191101 519061 191113 519064
rect 191147 519061 191159 519095
rect 191101 519055 191159 519061
rect 200761 519095 200819 519101
rect 200761 519061 200773 519095
rect 200807 519092 200819 519095
rect 209777 519095 209835 519101
rect 209777 519092 209789 519095
rect 200807 519064 209789 519092
rect 200807 519061 200819 519064
rect 200761 519055 200819 519061
rect 209777 519061 209789 519064
rect 209823 519061 209835 519095
rect 209777 519055 209835 519061
rect 219345 519095 219403 519101
rect 219345 519061 219357 519095
rect 219391 519092 219403 519095
rect 306944 519092 306972 519200
rect 316773 519197 316785 519200
rect 316819 519197 316831 519231
rect 316773 519191 316831 519197
rect 316865 519231 316923 519237
rect 316865 519197 316877 519231
rect 316911 519228 316923 519231
rect 325697 519231 325755 519237
rect 325697 519228 325709 519231
rect 316911 519200 325709 519228
rect 316911 519197 316923 519200
rect 316865 519191 316923 519197
rect 325697 519197 325709 519200
rect 325743 519197 325755 519231
rect 325697 519191 325755 519197
rect 307021 519163 307079 519169
rect 307021 519129 307033 519163
rect 307067 519160 307079 519163
rect 345032 519160 345060 519256
rect 307067 519132 345060 519160
rect 345109 519163 345167 519169
rect 307067 519129 307079 519132
rect 307021 519123 307079 519129
rect 345109 519129 345121 519163
rect 345155 519160 345167 519163
rect 355244 519160 355272 519268
rect 360286 519256 360292 519268
rect 360344 519256 360350 519308
rect 345155 519132 355272 519160
rect 345155 519129 345167 519132
rect 345109 519123 345167 519129
rect 219391 519064 306972 519092
rect 307113 519095 307171 519101
rect 219391 519061 219403 519064
rect 219345 519055 219403 519061
rect 307113 519061 307125 519095
rect 307159 519092 307171 519095
rect 316681 519095 316739 519101
rect 316681 519092 316693 519095
rect 307159 519064 316693 519092
rect 307159 519061 307171 519064
rect 307113 519055 307171 519061
rect 316681 519061 316693 519064
rect 316727 519061 316739 519095
rect 316681 519055 316739 519061
rect 316773 519095 316831 519101
rect 316773 519061 316785 519095
rect 316819 519092 316831 519095
rect 325697 519095 325755 519101
rect 325697 519092 325709 519095
rect 316819 519064 325709 519092
rect 316819 519061 316831 519064
rect 316773 519055 316831 519061
rect 325697 519061 325709 519064
rect 325743 519061 325755 519095
rect 325697 519055 325755 519061
rect 335265 519095 335323 519101
rect 335265 519061 335277 519095
rect 335311 519092 335323 519095
rect 349985 519095 350043 519101
rect 349985 519092 349997 519095
rect 335311 519064 349997 519092
rect 335311 519061 335323 519064
rect 335265 519055 335323 519061
rect 349985 519061 349997 519064
rect 350031 519061 350043 519095
rect 349985 519055 350043 519061
rect 3418 518984 3424 519036
rect 3476 519024 3482 519036
rect 355137 519027 355195 519033
rect 355137 519024 355149 519027
rect 3476 518996 306972 519024
rect 3476 518984 3482 518996
rect 4798 518916 4804 518968
rect 4856 518956 4862 518968
rect 17313 518959 17371 518965
rect 17313 518956 17325 518959
rect 4856 518928 17325 518956
rect 4856 518916 4862 518928
rect 17313 518925 17325 518928
rect 17359 518925 17371 518959
rect 17313 518919 17371 518925
rect 26789 518959 26847 518965
rect 26789 518925 26801 518959
rect 26835 518956 26847 518959
rect 36633 518959 36691 518965
rect 36633 518956 36645 518959
rect 26835 518928 36645 518956
rect 26835 518925 26847 518928
rect 26789 518919 26847 518925
rect 36633 518925 36645 518928
rect 36679 518925 36691 518959
rect 36633 518919 36691 518925
rect 46109 518959 46167 518965
rect 46109 518925 46121 518959
rect 46155 518956 46167 518959
rect 55953 518959 56011 518965
rect 55953 518956 55965 518959
rect 46155 518928 55965 518956
rect 46155 518925 46167 518928
rect 46109 518919 46167 518925
rect 55953 518925 55965 518928
rect 55999 518925 56011 518959
rect 55953 518919 56011 518925
rect 65429 518959 65487 518965
rect 65429 518925 65441 518959
rect 65475 518956 65487 518959
rect 75273 518959 75331 518965
rect 75273 518956 75285 518959
rect 65475 518928 75285 518956
rect 65475 518925 65487 518928
rect 65429 518919 65487 518925
rect 75273 518925 75285 518928
rect 75319 518925 75331 518959
rect 75273 518919 75331 518925
rect 84749 518959 84807 518965
rect 84749 518925 84761 518959
rect 84795 518956 84807 518959
rect 94593 518959 94651 518965
rect 94593 518956 94605 518959
rect 84795 518928 94605 518956
rect 84795 518925 84807 518928
rect 84749 518919 84807 518925
rect 94593 518925 94605 518928
rect 94639 518925 94651 518959
rect 94593 518919 94651 518925
rect 104069 518959 104127 518965
rect 104069 518925 104081 518959
rect 104115 518956 104127 518959
rect 113913 518959 113971 518965
rect 113913 518956 113925 518959
rect 104115 518928 113925 518956
rect 104115 518925 104127 518928
rect 104069 518919 104127 518925
rect 113913 518925 113925 518928
rect 113959 518925 113971 518959
rect 113913 518919 113971 518925
rect 123389 518959 123447 518965
rect 123389 518925 123401 518959
rect 123435 518956 123447 518959
rect 133233 518959 133291 518965
rect 133233 518956 133245 518959
rect 123435 518928 133245 518956
rect 123435 518925 123447 518928
rect 123389 518919 123447 518925
rect 133233 518925 133245 518928
rect 133279 518925 133291 518959
rect 133233 518919 133291 518925
rect 142709 518959 142767 518965
rect 142709 518925 142721 518959
rect 142755 518956 142767 518959
rect 152553 518959 152611 518965
rect 152553 518956 152565 518959
rect 142755 518928 152565 518956
rect 142755 518925 142767 518928
rect 142709 518919 142767 518925
rect 152553 518925 152565 518928
rect 152599 518925 152611 518959
rect 152553 518919 152611 518925
rect 162029 518959 162087 518965
rect 162029 518925 162041 518959
rect 162075 518956 162087 518959
rect 171873 518959 171931 518965
rect 171873 518956 171885 518959
rect 162075 518928 171885 518956
rect 162075 518925 162087 518928
rect 162029 518919 162087 518925
rect 171873 518925 171885 518928
rect 171919 518925 171931 518959
rect 171873 518919 171931 518925
rect 181533 518959 181591 518965
rect 181533 518925 181545 518959
rect 181579 518956 181591 518959
rect 188341 518959 188399 518965
rect 188341 518956 188353 518959
rect 181579 518928 188353 518956
rect 181579 518925 181591 518928
rect 181533 518919 181591 518925
rect 188341 518925 188353 518928
rect 188387 518925 188399 518959
rect 188341 518919 188399 518925
rect 200669 518959 200727 518965
rect 200669 518925 200681 518959
rect 200715 518956 200727 518959
rect 209777 518959 209835 518965
rect 209777 518956 209789 518959
rect 200715 518928 209789 518956
rect 200715 518925 200727 518928
rect 200669 518919 200727 518925
rect 209777 518925 209789 518928
rect 209823 518925 209835 518959
rect 209777 518919 209835 518925
rect 219345 518959 219403 518965
rect 219345 518925 219357 518959
rect 219391 518956 219403 518959
rect 306837 518959 306895 518965
rect 306837 518956 306849 518959
rect 219391 518928 306849 518956
rect 219391 518925 219403 518928
rect 219345 518919 219403 518925
rect 306837 518925 306849 518928
rect 306883 518925 306895 518959
rect 306837 518919 306895 518925
rect 306944 518888 306972 518996
rect 311912 518996 355149 519024
rect 311912 518956 311940 518996
rect 355137 518993 355149 518996
rect 355183 518993 355195 519027
rect 355137 518987 355195 518993
rect 307128 518928 311940 518956
rect 316681 518959 316739 518965
rect 307128 518888 307156 518928
rect 316681 518925 316693 518959
rect 316727 518956 316739 518959
rect 325697 518959 325755 518965
rect 325697 518956 325709 518959
rect 316727 518928 325709 518956
rect 316727 518925 316739 518928
rect 316681 518919 316739 518925
rect 325697 518925 325709 518928
rect 325743 518925 325755 518959
rect 325697 518919 325755 518925
rect 335265 518959 335323 518965
rect 335265 518925 335277 518959
rect 335311 518956 335323 518959
rect 345017 518959 345075 518965
rect 345017 518956 345029 518959
rect 335311 518928 345029 518956
rect 335311 518925 335323 518928
rect 335265 518919 335323 518925
rect 345017 518925 345029 518928
rect 345063 518925 345075 518959
rect 345017 518919 345075 518925
rect 306944 518860 307156 518888
rect 370314 518644 370320 518696
rect 370372 518684 370378 518696
rect 375282 518684 375288 518696
rect 370372 518656 375288 518684
rect 370372 518644 370378 518656
rect 375282 518644 375288 518656
rect 375340 518644 375346 518696
rect 3510 518236 3516 518288
rect 3568 518276 3574 518288
rect 351825 518279 351883 518285
rect 351825 518276 351837 518279
rect 3568 518248 351837 518276
rect 3568 518236 3574 518248
rect 351825 518245 351837 518248
rect 351871 518245 351883 518279
rect 351825 518239 351883 518245
rect 179417 518211 179475 518217
rect 179417 518177 179429 518211
rect 179463 518208 179475 518211
rect 580350 518208 580356 518220
rect 179463 518180 580356 518208
rect 179463 518177 179475 518180
rect 179417 518171 179475 518177
rect 580350 518168 580356 518180
rect 580408 518168 580414 518220
rect 50982 517828 50988 517880
rect 51040 517868 51046 517880
rect 57882 517868 57888 517880
rect 51040 517840 57888 517868
rect 51040 517828 51046 517840
rect 57882 517828 57888 517840
rect 57940 517828 57946 517880
rect 70302 517828 70308 517880
rect 70360 517868 70366 517880
rect 77202 517868 77208 517880
rect 70360 517840 77208 517868
rect 70360 517828 70366 517840
rect 77202 517828 77208 517840
rect 77260 517828 77266 517880
rect 89622 517828 89628 517880
rect 89680 517868 89686 517880
rect 96522 517868 96528 517880
rect 89680 517840 96528 517868
rect 89680 517828 89686 517840
rect 96522 517828 96528 517840
rect 96580 517828 96586 517880
rect 108942 517828 108948 517880
rect 109000 517868 109006 517880
rect 115842 517868 115848 517880
rect 109000 517840 115848 517868
rect 109000 517828 109006 517840
rect 115842 517828 115848 517840
rect 115900 517828 115906 517880
rect 128262 517828 128268 517880
rect 128320 517868 128326 517880
rect 135162 517868 135168 517880
rect 128320 517840 135168 517868
rect 128320 517828 128326 517840
rect 135162 517828 135168 517840
rect 135220 517828 135226 517880
rect 147582 517828 147588 517880
rect 147640 517868 147646 517880
rect 154482 517868 154488 517880
rect 147640 517840 154488 517868
rect 147640 517828 147646 517840
rect 154482 517828 154488 517840
rect 154540 517828 154546 517880
rect 27614 517556 27620 517608
rect 27672 517596 27678 517608
rect 37182 517596 37188 517608
rect 27672 517568 37188 517596
rect 27672 517556 27678 517568
rect 37182 517556 37188 517568
rect 37240 517556 37246 517608
rect 369762 510552 369768 510604
rect 369820 510592 369826 510604
rect 579982 510592 579988 510604
rect 369820 510564 579988 510592
rect 369820 510552 369826 510564
rect 579982 510552 579988 510564
rect 580040 510552 580046 510604
rect 579706 510212 579712 510264
rect 579764 510252 579770 510264
rect 579982 510252 579988 510264
rect 579764 510224 579988 510252
rect 579764 510212 579770 510224
rect 579982 510212 579988 510224
rect 580040 510212 580046 510264
rect 371142 499468 371148 499520
rect 371200 499508 371206 499520
rect 579890 499508 579896 499520
rect 371200 499480 579896 499508
rect 371200 499468 371206 499480
rect 579890 499468 579896 499480
rect 579948 499468 579954 499520
rect 2774 495524 2780 495576
rect 2832 495564 2838 495576
rect 4706 495564 4712 495576
rect 2832 495536 4712 495564
rect 2832 495524 2838 495536
rect 4706 495524 4712 495536
rect 4764 495524 4770 495576
rect 398742 486004 398748 486056
rect 398800 486044 398806 486056
rect 405642 486044 405648 486056
rect 398800 486016 405648 486044
rect 398800 486004 398806 486016
rect 405642 486004 405648 486016
rect 405700 486004 405706 486056
rect 371050 463632 371056 463684
rect 371108 463672 371114 463684
rect 579890 463672 579896 463684
rect 371108 463644 579896 463672
rect 371108 463632 371114 463644
rect 579890 463632 579896 463644
rect 579948 463632 579954 463684
rect 370958 452548 370964 452600
rect 371016 452588 371022 452600
rect 579890 452588 579896 452600
rect 371016 452560 579896 452588
rect 371016 452548 371022 452560
rect 579890 452548 579896 452560
rect 579948 452548 579954 452600
rect 3050 452412 3056 452464
rect 3108 452452 3114 452464
rect 6362 452452 6368 452464
rect 3108 452424 6368 452452
rect 3108 452412 3114 452424
rect 6362 452412 6368 452424
rect 6420 452412 6426 452464
rect 370866 440172 370872 440224
rect 370924 440212 370930 440224
rect 579890 440212 579896 440224
rect 370924 440184 579896 440212
rect 370924 440172 370930 440184
rect 579890 440172 579896 440184
rect 579948 440172 579954 440224
rect 3142 424056 3148 424108
rect 3200 424096 3206 424108
rect 6270 424096 6276 424108
rect 3200 424068 6276 424096
rect 3200 424056 3206 424068
rect 6270 424056 6276 424068
rect 6328 424056 6334 424108
rect 370774 416712 370780 416764
rect 370832 416752 370838 416764
rect 579890 416752 579896 416764
rect 370832 416724 579896 416752
rect 370832 416712 370838 416724
rect 579890 416712 579896 416724
rect 579948 416712 579954 416764
rect 370682 405628 370688 405680
rect 370740 405668 370746 405680
rect 579890 405668 579896 405680
rect 370740 405640 579896 405668
rect 370740 405628 370746 405640
rect 579890 405628 579896 405640
rect 579948 405628 579954 405680
rect 370590 393252 370596 393304
rect 370648 393292 370654 393304
rect 579890 393292 579896 393304
rect 370648 393264 579896 393292
rect 370648 393252 370654 393264
rect 579890 393252 579896 393264
rect 579948 393252 579954 393304
rect 2774 380604 2780 380656
rect 2832 380644 2838 380656
rect 5442 380644 5448 380656
rect 2832 380616 5448 380644
rect 2832 380604 2838 380616
rect 5442 380604 5448 380616
rect 5500 380604 5506 380656
rect 369670 369792 369676 369844
rect 369728 369832 369734 369844
rect 579890 369832 579896 369844
rect 369728 369804 579896 369832
rect 369728 369792 369734 369804
rect 579890 369792 579896 369804
rect 579948 369792 579954 369844
rect 2774 366936 2780 366988
rect 2832 366976 2838 366988
rect 5350 366976 5356 366988
rect 2832 366948 5356 366976
rect 2832 366936 2838 366948
rect 5350 366936 5356 366948
rect 5408 366936 5414 366988
rect 369578 346332 369584 346384
rect 369636 346372 369642 346384
rect 580074 346372 580080 346384
rect 369636 346344 580080 346372
rect 369636 346332 369642 346344
rect 580074 346332 580080 346344
rect 580132 346332 580138 346384
rect 3142 324164 3148 324216
rect 3200 324204 3206 324216
rect 6178 324204 6184 324216
rect 3200 324176 6184 324204
rect 3200 324164 3206 324176
rect 6178 324164 6184 324176
rect 6236 324164 6242 324216
rect 369670 322872 369676 322924
rect 369728 322912 369734 322924
rect 580074 322912 580080 322924
rect 369728 322884 580080 322912
rect 369728 322872 369734 322884
rect 580074 322872 580080 322884
rect 580132 322872 580138 322924
rect 3326 280100 3332 280152
rect 3384 280140 3390 280152
rect 10318 280140 10324 280152
rect 3384 280112 10324 280140
rect 3384 280100 3390 280112
rect 10318 280100 10324 280112
rect 10376 280100 10382 280152
rect 2774 266024 2780 266076
rect 2832 266064 2838 266076
rect 5258 266064 5264 266076
rect 2832 266036 5264 266064
rect 2832 266024 2838 266036
rect 5258 266024 5264 266036
rect 5316 266024 5322 266076
rect 3326 237328 3332 237380
rect 3384 237368 3390 237380
rect 13078 237368 13084 237380
rect 3384 237340 13084 237368
rect 3384 237328 3390 237340
rect 13078 237328 13084 237340
rect 13136 237328 13142 237380
rect 315758 219376 315764 219428
rect 315816 219416 315822 219428
rect 315942 219416 315948 219428
rect 315816 219388 315948 219416
rect 315816 219376 315822 219388
rect 315942 219376 315948 219388
rect 316000 219376 316006 219428
rect 334618 218152 334624 218204
rect 334676 218192 334682 218204
rect 339405 218195 339463 218201
rect 339405 218192 339417 218195
rect 334676 218164 339417 218192
rect 334676 218152 334682 218164
rect 339405 218161 339417 218164
rect 339451 218161 339463 218195
rect 339405 218155 339463 218161
rect 223758 218084 223764 218136
rect 223816 218124 223822 218136
rect 223942 218124 223948 218136
rect 223816 218096 223948 218124
rect 223816 218084 223822 218096
rect 223942 218084 223948 218096
rect 224000 218084 224006 218136
rect 340138 218124 340144 218136
rect 331416 218096 340144 218124
rect 329285 218059 329343 218065
rect 223960 218028 224724 218056
rect 88978 217948 88984 218000
rect 89036 217988 89042 218000
rect 197078 217988 197084 218000
rect 89036 217960 197084 217988
rect 89036 217948 89042 217960
rect 197078 217948 197084 217960
rect 197136 217948 197142 218000
rect 218698 217948 218704 218000
rect 218756 217988 218762 218000
rect 223960 217988 223988 218028
rect 218756 217960 223988 217988
rect 218756 217948 218762 217960
rect 224034 217948 224040 218000
rect 224092 217988 224098 218000
rect 224586 217988 224592 218000
rect 224092 217960 224592 217988
rect 224092 217948 224098 217960
rect 224586 217948 224592 217960
rect 224644 217948 224650 218000
rect 224696 217988 224724 218028
rect 329285 218025 329297 218059
rect 329331 218056 329343 218059
rect 330478 218056 330484 218068
rect 329331 218028 330484 218056
rect 329331 218025 329343 218028
rect 329285 218019 329343 218025
rect 330478 218016 330484 218028
rect 330536 218016 330542 218068
rect 331416 218056 331444 218096
rect 340138 218084 340144 218096
rect 340196 218084 340202 218136
rect 331232 218028 331444 218056
rect 332321 218059 332379 218065
rect 244458 217988 244464 218000
rect 224696 217960 244464 217988
rect 244458 217948 244464 217960
rect 244516 217948 244522 218000
rect 266906 217948 266912 218000
rect 266964 217988 266970 218000
rect 275833 217991 275891 217997
rect 275833 217988 275845 217991
rect 266964 217960 275845 217988
rect 266964 217948 266970 217960
rect 275833 217957 275845 217960
rect 275879 217957 275891 217991
rect 275833 217951 275891 217957
rect 275925 217991 275983 217997
rect 275925 217957 275937 217991
rect 275971 217988 275983 217991
rect 279418 217988 279424 218000
rect 275971 217960 279424 217988
rect 275971 217957 275983 217960
rect 275925 217951 275983 217957
rect 279418 217948 279424 217960
rect 279476 217948 279482 218000
rect 281994 217948 282000 218000
rect 282052 217988 282058 218000
rect 308398 217988 308404 218000
rect 282052 217960 308404 217988
rect 282052 217948 282058 217960
rect 308398 217948 308404 217960
rect 308456 217948 308462 218000
rect 315850 217948 315856 218000
rect 315908 217988 315914 218000
rect 331232 217988 331260 218028
rect 332321 218025 332333 218059
rect 332367 218056 332379 218059
rect 334618 218056 334624 218068
rect 332367 218028 334624 218056
rect 332367 218025 332379 218028
rect 332321 218019 332379 218025
rect 334618 218016 334624 218028
rect 334676 218016 334682 218068
rect 340601 218059 340659 218065
rect 340601 218025 340613 218059
rect 340647 218056 340659 218059
rect 340647 218028 340828 218056
rect 340647 218025 340659 218028
rect 340601 218019 340659 218025
rect 340693 217991 340751 217997
rect 340693 217988 340705 217991
rect 315908 217960 331260 217988
rect 331324 217960 340705 217988
rect 315908 217948 315914 217960
rect 86218 217880 86224 217932
rect 86276 217920 86282 217932
rect 194686 217920 194692 217932
rect 86276 217892 194692 217920
rect 86276 217880 86282 217892
rect 194686 217880 194692 217892
rect 194744 217880 194750 217932
rect 196618 217880 196624 217932
rect 196676 217920 196682 217932
rect 212994 217920 213000 217932
rect 196676 217892 213000 217920
rect 196676 217880 196682 217892
rect 212994 217880 213000 217892
rect 213052 217880 213058 217932
rect 215202 217880 215208 217932
rect 215260 217920 215266 217932
rect 243630 217920 243636 217932
rect 215260 217892 243636 217920
rect 215260 217880 215266 217892
rect 243630 217880 243636 217892
rect 243688 217880 243694 217932
rect 271782 217880 271788 217932
rect 271840 217920 271846 217932
rect 283101 217923 283159 217929
rect 283101 217920 283113 217923
rect 271840 217892 283113 217920
rect 271840 217880 271846 217892
rect 283101 217889 283113 217892
rect 283147 217889 283159 217923
rect 283101 217883 283159 217889
rect 283190 217880 283196 217932
rect 283248 217920 283254 217932
rect 284110 217920 284116 217932
rect 283248 217892 284116 217920
rect 283248 217880 283254 217892
rect 284110 217880 284116 217892
rect 284168 217880 284174 217932
rect 284478 217880 284484 217932
rect 284536 217920 284542 217932
rect 285490 217920 285496 217932
rect 284536 217892 285496 217920
rect 284536 217880 284542 217892
rect 285490 217880 285496 217892
rect 285548 217880 285554 217932
rect 286502 217880 286508 217932
rect 286560 217920 286566 217932
rect 286962 217920 286968 217932
rect 286560 217892 286968 217920
rect 286560 217880 286566 217892
rect 286962 217880 286968 217892
rect 287020 217880 287026 217932
rect 287698 217880 287704 217932
rect 287756 217920 287762 217932
rect 288342 217920 288348 217932
rect 287756 217892 288348 217920
rect 287756 217880 287762 217892
rect 288342 217880 288348 217892
rect 288400 217880 288406 217932
rect 289354 217880 289360 217932
rect 289412 217920 289418 217932
rect 289722 217920 289728 217932
rect 289412 217892 289728 217920
rect 289412 217880 289418 217892
rect 289722 217880 289728 217892
rect 289780 217880 289786 217932
rect 290550 217880 290556 217932
rect 290608 217920 290614 217932
rect 291010 217920 291016 217932
rect 290608 217892 291016 217920
rect 290608 217880 290614 217892
rect 291010 217880 291016 217892
rect 291068 217880 291074 217932
rect 291378 217880 291384 217932
rect 291436 217920 291442 217932
rect 292482 217920 292488 217932
rect 291436 217892 292488 217920
rect 291436 217880 291442 217892
rect 292482 217880 292488 217892
rect 292540 217880 292546 217932
rect 293862 217880 293868 217932
rect 293920 217920 293926 217932
rect 319438 217920 319444 217932
rect 293920 217892 319444 217920
rect 293920 217880 293926 217892
rect 319438 217880 319444 217892
rect 319496 217880 319502 217932
rect 320818 217880 320824 217932
rect 320876 217920 320882 217932
rect 321557 217923 321615 217929
rect 321557 217920 321569 217923
rect 320876 217892 321569 217920
rect 320876 217880 320882 217892
rect 321557 217889 321569 217892
rect 321603 217889 321615 217923
rect 321557 217883 321615 217889
rect 321646 217880 321652 217932
rect 321704 217920 321710 217932
rect 322658 217920 322664 217932
rect 321704 217892 322664 217920
rect 321704 217880 321710 217892
rect 322658 217880 322664 217892
rect 322716 217880 322722 217932
rect 323581 217923 323639 217929
rect 323581 217889 323593 217923
rect 323627 217920 323639 217923
rect 329285 217923 329343 217929
rect 329285 217920 329297 217923
rect 323627 217892 329297 217920
rect 323627 217889 323639 217892
rect 323581 217883 323639 217889
rect 329285 217889 329297 217892
rect 329331 217889 329343 217923
rect 329285 217883 329343 217889
rect 329374 217880 329380 217932
rect 329432 217920 329438 217932
rect 331324 217920 331352 217960
rect 340693 217957 340705 217960
rect 340739 217957 340751 217991
rect 340800 217988 340828 218028
rect 340800 217960 349200 217988
rect 340693 217951 340751 217957
rect 329432 217892 331352 217920
rect 329432 217880 329438 217892
rect 77938 217812 77944 217864
rect 77996 217852 78002 217864
rect 187326 217852 187332 217864
rect 77996 217824 187332 217852
rect 77996 217812 78002 217824
rect 187326 217812 187332 217824
rect 187384 217812 187390 217864
rect 212350 217812 212356 217864
rect 212408 217852 212414 217864
rect 240778 217852 240784 217864
rect 212408 217824 240784 217852
rect 212408 217812 212414 217824
rect 240778 217812 240784 217824
rect 240836 217812 240842 217864
rect 281537 217855 281595 217861
rect 281537 217852 281549 217855
rect 275940 217824 281549 217852
rect 275940 217796 275968 217824
rect 281537 217821 281549 217824
rect 281583 217821 281595 217855
rect 281537 217815 281595 217821
rect 281721 217855 281779 217861
rect 281721 217821 281733 217855
rect 281767 217852 281779 217855
rect 298738 217852 298744 217864
rect 281767 217824 298744 217852
rect 281767 217821 281779 217824
rect 281721 217815 281779 217821
rect 298738 217812 298744 217824
rect 298796 217812 298802 217864
rect 301222 217812 301228 217864
rect 301280 217852 301286 217864
rect 332321 217855 332379 217861
rect 332321 217852 332333 217855
rect 301280 217824 332333 217852
rect 301280 217812 301286 217824
rect 332321 217821 332333 217824
rect 332367 217821 332379 217855
rect 332321 217815 332379 217821
rect 332413 217855 332471 217861
rect 332413 217821 332425 217855
rect 332459 217852 332471 217855
rect 335357 217855 335415 217861
rect 335357 217852 335369 217855
rect 332459 217824 335369 217852
rect 332459 217821 332471 217824
rect 332413 217815 332471 217821
rect 335357 217821 335369 217824
rect 335403 217821 335415 217855
rect 335357 217815 335415 217821
rect 335446 217812 335452 217864
rect 335504 217852 335510 217864
rect 336642 217852 336648 217864
rect 335504 217824 336648 217852
rect 335504 217812 335510 217824
rect 336642 217812 336648 217824
rect 336700 217812 336706 217864
rect 336734 217812 336740 217864
rect 336792 217852 336798 217864
rect 337746 217852 337752 217864
rect 336792 217824 337752 217852
rect 336792 217812 336798 217824
rect 337746 217812 337752 217824
rect 337804 217812 337810 217864
rect 337841 217855 337899 217861
rect 337841 217821 337853 217855
rect 337887 217852 337899 217855
rect 340601 217855 340659 217861
rect 340601 217852 340613 217855
rect 337887 217824 340613 217852
rect 337887 217821 337899 217824
rect 337841 217815 337899 217821
rect 340601 217821 340613 217824
rect 340647 217821 340659 217855
rect 340601 217815 340659 217821
rect 340782 217812 340788 217864
rect 340840 217852 340846 217864
rect 345566 217852 345572 217864
rect 340840 217824 345572 217852
rect 340840 217812 340846 217824
rect 345566 217812 345572 217824
rect 345624 217812 345630 217864
rect 345658 217812 345664 217864
rect 345716 217852 345722 217864
rect 346302 217852 346308 217864
rect 345716 217824 346308 217852
rect 345716 217812 345722 217824
rect 346302 217812 346308 217824
rect 346360 217812 346366 217864
rect 346486 217812 346492 217864
rect 346544 217852 346550 217864
rect 347498 217852 347504 217864
rect 346544 217824 347504 217852
rect 346544 217812 346550 217824
rect 347498 217812 347504 217824
rect 347556 217812 347562 217864
rect 348142 217812 348148 217864
rect 348200 217852 348206 217864
rect 349062 217852 349068 217864
rect 348200 217824 349068 217852
rect 348200 217812 348206 217824
rect 349062 217812 349068 217824
rect 349120 217812 349126 217864
rect 349172 217852 349200 217960
rect 349338 217948 349344 218000
rect 349396 217988 349402 218000
rect 350442 217988 350448 218000
rect 349396 217960 350448 217988
rect 349396 217948 349402 217960
rect 350442 217948 350448 217960
rect 350500 217948 350506 218000
rect 358722 217948 358728 218000
rect 358780 217988 358786 218000
rect 469858 217988 469864 218000
rect 358780 217960 469864 217988
rect 358780 217948 358786 217960
rect 469858 217948 469864 217960
rect 469916 217948 469922 218000
rect 350537 217923 350595 217929
rect 350537 217889 350549 217923
rect 350583 217920 350595 217923
rect 358078 217920 358084 217932
rect 350583 217892 358084 217920
rect 350583 217889 350595 217892
rect 350537 217883 350595 217889
rect 358078 217880 358084 217892
rect 358136 217880 358142 217932
rect 366082 217880 366088 217932
rect 366140 217920 366146 217932
rect 478138 217920 478144 217932
rect 366140 217892 478144 217920
rect 366140 217880 366146 217892
rect 478138 217880 478144 217892
rect 478196 217880 478202 217932
rect 352558 217852 352564 217864
rect 349172 217824 352564 217852
rect 352558 217812 352564 217824
rect 352616 217812 352622 217864
rect 355042 217812 355048 217864
rect 355100 217852 355106 217864
rect 355594 217852 355600 217864
rect 355100 217824 355600 217852
rect 355100 217812 355106 217824
rect 355594 217812 355600 217824
rect 355652 217812 355658 217864
rect 362034 217812 362040 217864
rect 362092 217852 362098 217864
rect 362586 217852 362592 217864
rect 362092 217824 362592 217852
rect 362092 217812 362098 217824
rect 362586 217812 362592 217824
rect 362644 217812 362650 217864
rect 363690 217812 363696 217864
rect 363748 217852 363754 217864
rect 475378 217852 475384 217864
rect 363748 217824 475384 217852
rect 363748 217812 363754 217824
rect 475378 217812 475384 217824
rect 475436 217812 475442 217864
rect 75178 217744 75184 217796
rect 75236 217784 75242 217796
rect 185670 217784 185676 217796
rect 75236 217756 185676 217784
rect 75236 217744 75242 217756
rect 185670 217744 185676 217756
rect 185728 217744 185734 217796
rect 191190 217744 191196 217796
rect 191248 217784 191254 217796
rect 195882 217784 195888 217796
rect 191248 217756 195888 217784
rect 191248 217744 191254 217756
rect 195882 217744 195888 217756
rect 195940 217744 195946 217796
rect 209038 217744 209044 217796
rect 209096 217784 209102 217796
rect 239582 217784 239588 217796
rect 209096 217756 239588 217784
rect 209096 217744 209102 217756
rect 239582 217744 239588 217756
rect 239640 217744 239646 217796
rect 275922 217744 275928 217796
rect 275980 217744 275986 217796
rect 278314 217744 278320 217796
rect 278372 217784 278378 217796
rect 304258 217784 304264 217796
rect 278372 217756 304264 217784
rect 278372 217744 278378 217756
rect 304258 217744 304264 217756
rect 304316 217744 304322 217796
rect 318334 217744 318340 217796
rect 318392 217784 318398 217796
rect 350537 217787 350595 217793
rect 350537 217784 350549 217787
rect 318392 217756 350549 217784
rect 318392 217744 318398 217756
rect 350537 217753 350549 217756
rect 350583 217753 350595 217787
rect 350537 217747 350595 217753
rect 350626 217744 350632 217796
rect 350684 217784 350690 217796
rect 351822 217784 351828 217796
rect 350684 217756 351828 217784
rect 350684 217744 350690 217756
rect 351822 217744 351828 217756
rect 351880 217744 351886 217796
rect 354674 217744 354680 217796
rect 354732 217784 354738 217796
rect 355870 217784 355876 217796
rect 354732 217756 355876 217784
rect 354732 217744 354738 217756
rect 355870 217744 355876 217756
rect 355928 217744 355934 217796
rect 356698 217744 356704 217796
rect 356756 217784 356762 217796
rect 357342 217784 357348 217796
rect 356756 217756 357348 217784
rect 356756 217744 356762 217756
rect 357342 217744 357348 217756
rect 357400 217744 357406 217796
rect 357894 217744 357900 217796
rect 357952 217784 357958 217796
rect 358722 217784 358728 217796
rect 357952 217756 358728 217784
rect 357952 217744 357958 217756
rect 358722 217744 358728 217756
rect 358780 217744 358786 217796
rect 361574 217744 361580 217796
rect 361632 217784 361638 217796
rect 362770 217784 362776 217796
rect 361632 217756 362776 217784
rect 361632 217744 361638 217756
rect 362770 217744 362776 217756
rect 362828 217744 362834 217796
rect 364886 217744 364892 217796
rect 364944 217784 364950 217796
rect 365622 217784 365628 217796
rect 364944 217756 365628 217784
rect 364944 217744 364950 217756
rect 365622 217744 365628 217756
rect 365680 217744 365686 217796
rect 365714 217744 365720 217796
rect 365772 217784 365778 217796
rect 366818 217784 366824 217796
rect 365772 217756 366824 217784
rect 365772 217744 365778 217756
rect 366818 217744 366824 217756
rect 366876 217744 366882 217796
rect 367278 217744 367284 217796
rect 367336 217784 367342 217796
rect 368382 217784 368388 217796
rect 367336 217756 368388 217784
rect 367336 217744 367342 217756
rect 368382 217744 368388 217756
rect 368440 217744 368446 217796
rect 368566 217744 368572 217796
rect 368624 217784 368630 217796
rect 480898 217784 480904 217796
rect 368624 217756 480904 217784
rect 368624 217744 368630 217756
rect 480898 217744 480904 217756
rect 480956 217744 480962 217796
rect 71038 217676 71044 217728
rect 71096 217716 71102 217728
rect 170861 217719 170919 217725
rect 170861 217716 170873 217719
rect 71096 217688 170873 217716
rect 71096 217676 71102 217688
rect 170861 217685 170873 217688
rect 170907 217685 170919 217719
rect 170861 217679 170919 217685
rect 170953 217719 171011 217725
rect 170953 217685 170965 217719
rect 170999 217716 171011 217719
rect 175458 217716 175464 217728
rect 170999 217688 175464 217716
rect 170999 217685 171011 217688
rect 170953 217679 171011 217685
rect 175458 217676 175464 217688
rect 175516 217676 175522 217728
rect 180153 217719 180211 217725
rect 180153 217685 180165 217719
rect 180199 217716 180211 217719
rect 210142 217716 210148 217728
rect 180199 217688 210148 217716
rect 180199 217685 180211 217688
rect 180153 217679 180211 217685
rect 210142 217676 210148 217688
rect 210200 217676 210206 217728
rect 212353 217719 212411 217725
rect 212353 217685 212365 217719
rect 212399 217716 212411 217719
rect 242802 217716 242808 217728
rect 212399 217688 242808 217716
rect 212399 217685 212411 217688
rect 212353 217679 212411 217685
rect 242802 217676 242808 217688
rect 242860 217676 242866 217728
rect 256602 217676 256608 217728
rect 256660 217716 256666 217728
rect 257890 217716 257896 217728
rect 256660 217688 257896 217716
rect 256660 217676 256666 217688
rect 257890 217676 257896 217688
rect 257948 217676 257954 217728
rect 262858 217676 262864 217728
rect 262916 217716 262922 217728
rect 263502 217716 263508 217728
rect 262916 217688 263508 217716
rect 262916 217676 262922 217688
rect 263502 217676 263508 217688
rect 263560 217676 263566 217728
rect 264882 217676 264888 217728
rect 264940 217716 264946 217728
rect 265618 217716 265624 217728
rect 264940 217688 265624 217716
rect 264940 217676 264946 217688
rect 265618 217676 265624 217688
rect 265676 217676 265682 217728
rect 267734 217676 267740 217728
rect 267792 217716 267798 217728
rect 268930 217716 268936 217728
rect 267792 217688 268936 217716
rect 267792 217676 267798 217688
rect 268930 217676 268936 217688
rect 268988 217676 268994 217728
rect 270586 217676 270592 217728
rect 270644 217716 270650 217728
rect 271782 217716 271788 217728
rect 270644 217688 271788 217716
rect 270644 217676 270650 217688
rect 271782 217676 271788 217688
rect 271840 217676 271846 217728
rect 277946 217676 277952 217728
rect 278004 217716 278010 217728
rect 278682 217716 278688 217728
rect 278004 217688 278688 217716
rect 278004 217676 278010 217688
rect 278682 217676 278688 217688
rect 278740 217676 278746 217728
rect 279142 217676 279148 217728
rect 279200 217716 279206 217728
rect 280062 217716 280068 217728
rect 279200 217688 280068 217716
rect 279200 217676 279206 217688
rect 280062 217676 280068 217688
rect 280120 217676 280126 217728
rect 280338 217676 280344 217728
rect 280396 217716 280402 217728
rect 281442 217716 281448 217728
rect 280396 217688 281448 217716
rect 280396 217676 280402 217688
rect 281442 217676 281448 217688
rect 281500 217676 281506 217728
rect 281537 217719 281595 217725
rect 281537 217685 281549 217719
rect 281583 217716 281595 217719
rect 292577 217719 292635 217725
rect 292577 217716 292589 217719
rect 281583 217688 292589 217716
rect 281583 217685 281595 217688
rect 281537 217679 281595 217685
rect 292577 217685 292589 217688
rect 292623 217685 292635 217719
rect 292577 217679 292635 217685
rect 292666 217676 292672 217728
rect 292724 217716 292730 217728
rect 293862 217716 293868 217728
rect 292724 217688 293868 217716
rect 292724 217676 292730 217688
rect 293862 217676 293868 217688
rect 293920 217676 293926 217728
rect 295886 217676 295892 217728
rect 295944 217716 295950 217728
rect 296530 217716 296536 217728
rect 295944 217688 296536 217716
rect 295944 217676 295950 217688
rect 296530 217676 296536 217688
rect 296588 217676 296594 217728
rect 296714 217676 296720 217728
rect 296772 217716 296778 217728
rect 298002 217716 298008 217728
rect 296772 217688 298008 217716
rect 296772 217676 296778 217688
rect 298002 217676 298008 217688
rect 298060 217676 298066 217728
rect 300394 217676 300400 217728
rect 300452 217716 300458 217728
rect 300762 217716 300768 217728
rect 300452 217688 300768 217716
rect 300452 217676 300458 217688
rect 300762 217676 300768 217688
rect 300820 217676 300826 217728
rect 301590 217676 301596 217728
rect 301648 217716 301654 217728
rect 302142 217716 302148 217728
rect 301648 217688 302148 217716
rect 301648 217676 301654 217688
rect 302142 217676 302148 217688
rect 302200 217676 302206 217728
rect 303614 217676 303620 217728
rect 303672 217716 303678 217728
rect 331306 217716 331312 217728
rect 303672 217688 331312 217716
rect 303672 217676 303678 217688
rect 331306 217676 331312 217688
rect 331364 217676 331370 217728
rect 331398 217676 331404 217728
rect 331456 217716 331462 217728
rect 332410 217716 332416 217728
rect 331456 217688 332416 217716
rect 331456 217676 331462 217688
rect 332410 217676 332416 217688
rect 332468 217676 332474 217728
rect 333422 217676 333428 217728
rect 333480 217716 333486 217728
rect 333790 217716 333796 217728
rect 333480 217688 333796 217716
rect 333480 217676 333486 217688
rect 333790 217676 333796 217688
rect 333848 217676 333854 217728
rect 334710 217676 334716 217728
rect 334768 217716 334774 217728
rect 335262 217716 335268 217728
rect 334768 217688 335268 217716
rect 334768 217676 334774 217688
rect 335262 217676 335268 217688
rect 335320 217676 335326 217728
rect 335906 217676 335912 217728
rect 335964 217716 335970 217728
rect 336550 217716 336556 217728
rect 335964 217688 336556 217716
rect 335964 217676 335970 217688
rect 336550 217676 336556 217688
rect 336608 217676 336614 217728
rect 336645 217719 336703 217725
rect 336645 217685 336657 217719
rect 336691 217716 336703 217719
rect 337473 217719 337531 217725
rect 337473 217716 337485 217719
rect 336691 217688 337485 217716
rect 336691 217685 336703 217688
rect 336645 217679 336703 217685
rect 337473 217685 337485 217688
rect 337519 217685 337531 217719
rect 337473 217679 337531 217685
rect 337562 217676 337568 217728
rect 337620 217716 337626 217728
rect 337930 217716 337936 217728
rect 337620 217688 337936 217716
rect 337620 217676 337626 217688
rect 337930 217676 337936 217688
rect 337988 217676 337994 217728
rect 338298 217676 338304 217728
rect 338356 217716 338362 217728
rect 339402 217716 339408 217728
rect 338356 217688 339408 217716
rect 338356 217676 338362 217688
rect 339402 217676 339408 217688
rect 339460 217676 339466 217728
rect 339497 217719 339555 217725
rect 339497 217685 339509 217719
rect 339543 217716 339555 217719
rect 341058 217716 341064 217728
rect 339543 217688 341064 217716
rect 339543 217685 339555 217688
rect 339497 217679 339555 217685
rect 341058 217676 341064 217688
rect 341116 217676 341122 217728
rect 341150 217676 341156 217728
rect 341208 217716 341214 217728
rect 342070 217716 342076 217728
rect 341208 217688 342076 217716
rect 341208 217676 341214 217688
rect 342070 217676 342076 217688
rect 342128 217676 342134 217728
rect 342438 217676 342444 217728
rect 342496 217716 342502 217728
rect 343450 217716 343456 217728
rect 342496 217688 343456 217716
rect 342496 217676 342502 217688
rect 343450 217676 343456 217688
rect 343508 217676 343514 217728
rect 345290 217676 345296 217728
rect 345348 217716 345354 217728
rect 346118 217716 346124 217728
rect 345348 217688 346124 217716
rect 345348 217676 345354 217688
rect 346118 217676 346124 217688
rect 346176 217676 346182 217728
rect 347406 217676 347412 217728
rect 347464 217716 347470 217728
rect 347682 217716 347688 217728
rect 347464 217688 347688 217716
rect 347464 217676 347470 217688
rect 347682 217676 347688 217688
rect 347740 217676 347746 217728
rect 348510 217676 348516 217728
rect 348568 217716 348574 217728
rect 348970 217716 348976 217728
rect 348568 217688 348976 217716
rect 348568 217676 348574 217688
rect 348970 217676 348976 217688
rect 349028 217676 349034 217728
rect 349798 217676 349804 217728
rect 349856 217716 349862 217728
rect 350350 217716 350356 217728
rect 349856 217688 350356 217716
rect 349856 217676 349862 217688
rect 350350 217676 350356 217688
rect 350408 217676 350414 217728
rect 350994 217676 351000 217728
rect 351052 217716 351058 217728
rect 351638 217716 351644 217728
rect 351052 217688 351644 217716
rect 351052 217676 351058 217688
rect 351638 217676 351644 217688
rect 351696 217676 351702 217728
rect 352190 217676 352196 217728
rect 352248 217716 352254 217728
rect 353110 217716 353116 217728
rect 352248 217688 353116 217716
rect 352248 217676 352254 217688
rect 353110 217676 353116 217688
rect 353168 217676 353174 217728
rect 353478 217676 353484 217728
rect 353536 217716 353542 217728
rect 354490 217716 354496 217728
rect 353536 217688 354496 217716
rect 353536 217676 353542 217688
rect 354490 217676 354496 217688
rect 354548 217676 354554 217728
rect 355502 217676 355508 217728
rect 355560 217716 355566 217728
rect 355962 217716 355968 217728
rect 355560 217688 355968 217716
rect 355560 217676 355566 217688
rect 355962 217676 355968 217688
rect 356020 217676 356026 217728
rect 356330 217676 356336 217728
rect 356388 217716 356394 217728
rect 357158 217716 357164 217728
rect 356388 217688 357164 217716
rect 356388 217676 356394 217688
rect 357158 217676 357164 217688
rect 357216 217676 357222 217728
rect 357526 217676 357532 217728
rect 357584 217716 357590 217728
rect 358538 217716 358544 217728
rect 357584 217688 358544 217716
rect 357584 217676 357590 217688
rect 358538 217676 358544 217688
rect 358596 217676 358602 217728
rect 359182 217676 359188 217728
rect 359240 217716 359246 217728
rect 360010 217716 360016 217728
rect 359240 217688 360016 217716
rect 359240 217676 359246 217688
rect 360010 217676 360016 217688
rect 360068 217676 360074 217728
rect 360378 217676 360384 217728
rect 360436 217716 360442 217728
rect 361482 217716 361488 217728
rect 360436 217688 361488 217716
rect 360436 217676 360442 217688
rect 361482 217676 361488 217688
rect 361540 217676 361546 217728
rect 362402 217676 362408 217728
rect 362460 217716 362466 217728
rect 362862 217716 362868 217728
rect 362460 217688 362868 217716
rect 362460 217676 362466 217688
rect 362862 217676 362868 217688
rect 362920 217676 362926 217728
rect 363230 217676 363236 217728
rect 363288 217716 363294 217728
rect 364150 217716 364156 217728
rect 363288 217688 364156 217716
rect 363288 217676 363294 217688
rect 364150 217676 364156 217688
rect 364208 217676 364214 217728
rect 364426 217676 364432 217728
rect 364484 217716 364490 217728
rect 365438 217716 365444 217728
rect 364484 217688 365444 217716
rect 364484 217676 364490 217688
rect 365438 217676 365444 217688
rect 365496 217676 365502 217728
rect 366542 217676 366548 217728
rect 366600 217716 366606 217728
rect 367002 217716 367008 217728
rect 366600 217688 367008 217716
rect 366600 217676 366606 217688
rect 367002 217676 367008 217688
rect 367060 217676 367066 217728
rect 367738 217676 367744 217728
rect 367796 217716 367802 217728
rect 368290 217716 368296 217728
rect 367796 217688 368296 217716
rect 367796 217676 367802 217688
rect 368290 217676 368296 217688
rect 368348 217676 368354 217728
rect 368934 217676 368940 217728
rect 368992 217716 368998 217728
rect 369670 217716 369676 217728
rect 368992 217688 369676 217716
rect 368992 217676 368998 217688
rect 369670 217676 369676 217688
rect 369728 217676 369734 217728
rect 369765 217719 369823 217725
rect 369765 217685 369777 217719
rect 369811 217716 369823 217719
rect 473998 217716 474004 217728
rect 369811 217688 474004 217716
rect 369811 217685 369823 217688
rect 369765 217679 369823 217685
rect 473998 217676 474004 217688
rect 474056 217676 474062 217728
rect 42058 217608 42064 217660
rect 42116 217648 42122 217660
rect 183646 217648 183652 217660
rect 42116 217620 183652 217648
rect 42116 217608 42122 217620
rect 183646 217608 183652 217620
rect 183704 217608 183710 217660
rect 188338 217608 188344 217660
rect 188396 217648 188402 217660
rect 193398 217648 193404 217660
rect 188396 217620 193404 217648
rect 188396 217608 188402 217620
rect 193398 217608 193404 217620
rect 193456 217608 193462 217660
rect 195422 217608 195428 217660
rect 195480 217648 195486 217660
rect 209314 217648 209320 217660
rect 195480 217620 209320 217648
rect 195480 217608 195486 217620
rect 209314 217608 209320 217620
rect 209372 217608 209378 217660
rect 212258 217608 212264 217660
rect 212316 217648 212322 217660
rect 242434 217648 242440 217660
rect 212316 217620 242440 217648
rect 212316 217608 212322 217620
rect 242434 217608 242440 217620
rect 242492 217608 242498 217660
rect 247770 217608 247776 217660
rect 247828 217648 247834 217660
rect 250622 217648 250628 217660
rect 247828 217620 250628 217648
rect 247828 217608 247834 217620
rect 250622 217608 250628 217620
rect 250680 217608 250686 217660
rect 255222 217608 255228 217660
rect 255280 217648 255286 217660
rect 257522 217648 257528 217660
rect 255280 217620 257528 217648
rect 255280 217608 255286 217620
rect 257522 217608 257528 217620
rect 257580 217608 257586 217660
rect 260742 217608 260748 217660
rect 260800 217648 260806 217660
rect 261570 217648 261576 217660
rect 260800 217620 261576 217648
rect 260800 217608 260806 217620
rect 261570 217608 261576 217620
rect 261628 217608 261634 217660
rect 264422 217608 264428 217660
rect 264480 217648 264486 217660
rect 272518 217648 272524 217660
rect 264480 217620 272524 217648
rect 264480 217608 264486 217620
rect 272518 217608 272524 217620
rect 272576 217608 272582 217660
rect 279602 217608 279608 217660
rect 279660 217648 279666 217660
rect 295337 217651 295395 217657
rect 295337 217648 295349 217651
rect 279660 217620 295349 217648
rect 279660 217608 279666 217620
rect 295337 217617 295349 217620
rect 295383 217617 295395 217651
rect 295337 217611 295395 217617
rect 295518 217608 295524 217660
rect 295576 217648 295582 217660
rect 296622 217648 296628 217660
rect 295576 217620 296628 217648
rect 295576 217608 295582 217620
rect 296622 217608 296628 217620
rect 296680 217608 296686 217660
rect 299566 217608 299572 217660
rect 299624 217648 299630 217660
rect 300578 217648 300584 217660
rect 299624 217620 300584 217648
rect 299624 217608 299630 217620
rect 300578 217608 300584 217620
rect 300636 217608 300642 217660
rect 302878 217648 302884 217660
rect 300688 217620 302884 217648
rect 35158 217540 35164 217592
rect 35216 217580 35222 217592
rect 181162 217580 181168 217592
rect 35216 217552 181168 217580
rect 35216 217540 35222 217552
rect 181162 217540 181168 217552
rect 181220 217540 181226 217592
rect 181346 217540 181352 217592
rect 181404 217580 181410 217592
rect 181898 217580 181904 217592
rect 181404 217552 181904 217580
rect 181404 217540 181410 217552
rect 181898 217540 181904 217552
rect 181956 217540 181962 217592
rect 195238 217540 195244 217592
rect 195296 217580 195302 217592
rect 206922 217580 206928 217592
rect 195296 217552 206928 217580
rect 195296 217540 195302 217552
rect 206922 217540 206928 217552
rect 206980 217540 206986 217592
rect 208302 217540 208308 217592
rect 208360 217580 208366 217592
rect 241146 217580 241152 217592
rect 208360 217552 241152 217580
rect 208360 217540 208366 217552
rect 241146 217540 241152 217552
rect 241204 217540 241210 217592
rect 245562 217540 245568 217592
rect 245620 217580 245626 217592
rect 253842 217580 253848 217592
rect 245620 217552 253848 217580
rect 245620 217540 245626 217552
rect 253842 217540 253848 217552
rect 253900 217540 253906 217592
rect 277118 217540 277124 217592
rect 277176 217580 277182 217592
rect 300688 217580 300716 217620
rect 302878 217608 302884 217620
rect 302936 217608 302942 217660
rect 319530 217608 319536 217660
rect 319588 217648 319594 217660
rect 434714 217648 434720 217660
rect 319588 217620 434720 217648
rect 319588 217608 319594 217620
rect 434714 217608 434720 217620
rect 434772 217608 434778 217660
rect 277176 217552 300716 217580
rect 277176 217540 277182 217552
rect 322382 217540 322388 217592
rect 322440 217580 322446 217592
rect 322842 217580 322848 217592
rect 322440 217552 322848 217580
rect 322440 217540 322446 217552
rect 322842 217540 322848 217552
rect 322900 217540 322906 217592
rect 324866 217540 324872 217592
rect 324924 217580 324930 217592
rect 325602 217580 325608 217592
rect 324924 217552 325608 217580
rect 324924 217540 324930 217552
rect 325602 217540 325608 217552
rect 325660 217540 325666 217592
rect 326062 217540 326068 217592
rect 326120 217580 326126 217592
rect 326982 217580 326988 217592
rect 326120 217552 326988 217580
rect 326120 217540 326126 217552
rect 326982 217540 326988 217552
rect 327040 217540 327046 217592
rect 327350 217540 327356 217592
rect 327408 217580 327414 217592
rect 328362 217580 328368 217592
rect 327408 217552 328368 217580
rect 327408 217540 327414 217552
rect 328362 217540 328368 217552
rect 328420 217540 328426 217592
rect 328546 217540 328552 217592
rect 328604 217580 328610 217592
rect 329650 217580 329656 217592
rect 328604 217552 329656 217580
rect 328604 217540 328610 217552
rect 329650 217540 329656 217552
rect 329708 217540 329714 217592
rect 330202 217540 330208 217592
rect 330260 217580 330266 217592
rect 331030 217580 331036 217592
rect 330260 217552 331036 217580
rect 330260 217540 330266 217552
rect 331030 217540 331036 217552
rect 331088 217540 331094 217592
rect 331125 217583 331183 217589
rect 331125 217549 331137 217583
rect 331171 217580 331183 217583
rect 442994 217580 443000 217592
rect 331171 217552 443000 217580
rect 331171 217549 331183 217552
rect 331125 217543 331183 217549
rect 442994 217540 443000 217552
rect 443052 217540 443058 217592
rect 32398 217472 32404 217524
rect 32456 217512 32462 217524
rect 168285 217515 168343 217521
rect 168285 217512 168297 217515
rect 32456 217484 168297 217512
rect 32456 217472 32462 217484
rect 168285 217481 168297 217484
rect 168331 217481 168343 217515
rect 170769 217515 170827 217521
rect 170769 217512 170781 217515
rect 168285 217475 168343 217481
rect 168392 217484 170781 217512
rect 31018 217404 31024 217456
rect 31076 217444 31082 217456
rect 167181 217447 167239 217453
rect 31076 217416 167132 217444
rect 31076 217404 31082 217416
rect 24118 217336 24124 217388
rect 24176 217376 24182 217388
rect 167104 217385 167132 217416
rect 167181 217413 167193 217447
rect 167227 217444 167239 217447
rect 168392 217444 168420 217484
rect 170769 217481 170781 217484
rect 170815 217481 170827 217515
rect 170769 217475 170827 217481
rect 170861 217515 170919 217521
rect 170861 217481 170873 217515
rect 170907 217512 170919 217515
rect 183186 217512 183192 217524
rect 170907 217484 183192 217512
rect 170907 217481 170919 217484
rect 170861 217475 170919 217481
rect 183186 217472 183192 217484
rect 183244 217472 183250 217524
rect 186958 217472 186964 217524
rect 187016 217512 187022 217524
rect 191006 217512 191012 217524
rect 187016 217484 191012 217512
rect 187016 217472 187022 217484
rect 191006 217472 191012 217484
rect 191064 217472 191070 217524
rect 195330 217472 195336 217524
rect 195388 217512 195394 217524
rect 204438 217512 204444 217524
rect 195388 217484 204444 217512
rect 195388 217472 195394 217484
rect 204438 217472 204444 217484
rect 204496 217472 204502 217524
rect 204898 217472 204904 217524
rect 204956 217512 204962 217524
rect 237558 217512 237564 217524
rect 204956 217484 237564 217512
rect 204956 217472 204962 217484
rect 237558 217472 237564 217484
rect 237616 217472 237622 217524
rect 238018 217472 238024 217524
rect 238076 217512 238082 217524
rect 245654 217512 245660 217524
rect 238076 217484 245660 217512
rect 238076 217472 238082 217484
rect 245654 217472 245660 217484
rect 245712 217472 245718 217524
rect 248322 217472 248328 217524
rect 248380 217512 248386 217524
rect 255038 217512 255044 217524
rect 248380 217484 255044 217512
rect 248380 217472 248386 217484
rect 255038 217472 255044 217484
rect 255096 217472 255102 217524
rect 281626 217472 281632 217524
rect 281684 217512 281690 217524
rect 309778 217512 309784 217524
rect 281684 217484 309784 217512
rect 281684 217472 281690 217484
rect 309778 217472 309784 217484
rect 309836 217472 309842 217524
rect 317138 217472 317144 217524
rect 317196 217512 317202 217524
rect 319993 217515 320051 217521
rect 319993 217512 320005 217515
rect 317196 217484 320005 217512
rect 317196 217472 317202 217484
rect 319993 217481 320005 217484
rect 320039 217481 320051 217515
rect 319993 217475 320051 217481
rect 321557 217515 321615 217521
rect 321557 217481 321569 217515
rect 321603 217512 321615 217515
rect 323581 217515 323639 217521
rect 323581 217512 323593 217515
rect 321603 217484 323593 217512
rect 321603 217481 321615 217484
rect 321557 217475 321615 217481
rect 323581 217481 323593 217484
rect 323627 217481 323639 217515
rect 323581 217475 323639 217481
rect 323670 217472 323676 217524
rect 323728 217512 323734 217524
rect 324222 217512 324228 217524
rect 323728 217484 324228 217512
rect 323728 217472 323734 217484
rect 324222 217472 324228 217484
rect 324280 217472 324286 217524
rect 324498 217472 324504 217524
rect 324556 217512 324562 217524
rect 449894 217512 449900 217524
rect 324556 217484 449900 217512
rect 324556 217472 324562 217484
rect 449894 217472 449900 217484
rect 449952 217472 449958 217524
rect 167227 217416 168420 217444
rect 168469 217447 168527 217453
rect 167227 217413 167239 217416
rect 167181 217407 167239 217413
rect 168469 217413 168481 217447
rect 168515 217444 168527 217447
rect 178770 217444 178776 217456
rect 168515 217416 178776 217444
rect 168515 217413 168527 217416
rect 168469 217407 168527 217413
rect 178770 217404 178776 217416
rect 178828 217404 178834 217456
rect 203518 217404 203524 217456
rect 203576 217444 203582 217456
rect 238294 217444 238300 217456
rect 203576 217416 238300 217444
rect 203576 217404 203582 217416
rect 238294 217404 238300 217416
rect 238352 217404 238358 217456
rect 238662 217404 238668 217456
rect 238720 217444 238726 217456
rect 251818 217444 251824 217456
rect 238720 217416 251824 217444
rect 238720 217404 238726 217416
rect 251818 217404 251824 217416
rect 251876 217404 251882 217456
rect 260006 217404 260012 217456
rect 260064 217444 260070 217456
rect 261478 217444 261484 217456
rect 260064 217416 261484 217444
rect 260064 217404 260070 217416
rect 261478 217404 261484 217416
rect 261536 217404 261542 217456
rect 269390 217404 269396 217456
rect 269448 217444 269454 217456
rect 270218 217444 270224 217456
rect 269448 217416 270224 217444
rect 269448 217404 269454 217416
rect 270218 217404 270224 217416
rect 270276 217404 270282 217456
rect 273806 217404 273812 217456
rect 273864 217444 273870 217456
rect 281721 217447 281779 217453
rect 281721 217444 281733 217447
rect 273864 217416 281733 217444
rect 273864 217404 273870 217416
rect 281721 217413 281733 217416
rect 281767 217413 281779 217447
rect 281721 217407 281779 217413
rect 281813 217447 281871 217453
rect 281813 217413 281825 217447
rect 281859 217444 281871 217447
rect 292669 217447 292727 217453
rect 281859 217416 292620 217444
rect 281859 217413 281871 217416
rect 281813 217407 281871 217413
rect 166997 217379 167055 217385
rect 166997 217376 167009 217379
rect 24176 217348 167009 217376
rect 24176 217336 24182 217348
rect 166997 217345 167009 217348
rect 167043 217345 167055 217379
rect 166997 217339 167055 217345
rect 167089 217379 167147 217385
rect 167089 217345 167101 217379
rect 167135 217345 167147 217379
rect 175090 217376 175096 217388
rect 167089 217339 167147 217345
rect 167196 217348 175096 217376
rect 17218 217268 17224 217320
rect 17276 217308 17282 217320
rect 167196 217308 167224 217348
rect 175090 217336 175096 217348
rect 175148 217336 175154 217388
rect 204162 217336 204168 217388
rect 204220 217376 204226 217388
rect 239950 217376 239956 217388
rect 204220 217348 239956 217376
rect 204220 217336 204226 217348
rect 239950 217336 239956 217348
rect 240008 217336 240014 217388
rect 240778 217336 240784 217388
rect 240836 217376 240842 217388
rect 249886 217376 249892 217388
rect 240836 217348 249892 217376
rect 240836 217336 240842 217348
rect 249886 217336 249892 217348
rect 249944 217336 249950 217388
rect 264054 217336 264060 217388
rect 264112 217376 264118 217388
rect 266998 217376 267004 217388
rect 264112 217348 267004 217376
rect 264112 217336 264118 217348
rect 266998 217336 267004 217348
rect 267056 217336 267062 217388
rect 276290 217336 276296 217388
rect 276348 217376 276354 217388
rect 277302 217376 277308 217388
rect 276348 217348 277308 217376
rect 276348 217336 276354 217348
rect 277302 217336 277308 217348
rect 277360 217336 277366 217388
rect 277486 217336 277492 217388
rect 277544 217376 277550 217388
rect 282917 217379 282975 217385
rect 282917 217376 282929 217379
rect 277544 217348 282929 217376
rect 277544 217336 277550 217348
rect 282917 217345 282929 217348
rect 282963 217345 282975 217379
rect 292592 217376 292620 217416
rect 292669 217413 292681 217447
rect 292715 217444 292727 217447
rect 301498 217444 301504 217456
rect 292715 217416 301504 217444
rect 292715 217413 292727 217416
rect 292669 217407 292727 217413
rect 301498 217404 301504 217416
rect 301556 217404 301562 217456
rect 306098 217404 306104 217456
rect 306156 217444 306162 217456
rect 322198 217444 322204 217456
rect 306156 217416 322204 217444
rect 306156 217404 306162 217416
rect 322198 217404 322204 217416
rect 322256 217404 322262 217456
rect 323210 217404 323216 217456
rect 323268 217444 323274 217456
rect 323268 217416 332548 217444
rect 323268 217404 323274 217416
rect 302970 217376 302976 217388
rect 292592 217348 302976 217376
rect 282917 217339 282975 217345
rect 302970 217336 302976 217348
rect 303028 217336 303034 217388
rect 310974 217336 310980 217388
rect 311032 217376 311038 217388
rect 311032 217348 312676 217376
rect 311032 217336 311038 217348
rect 17276 217280 167224 217308
rect 167273 217311 167331 217317
rect 17276 217268 17282 217280
rect 167273 217277 167285 217311
rect 167319 217308 167331 217311
rect 178310 217308 178316 217320
rect 167319 217280 178316 217308
rect 167319 217277 167331 217280
rect 167273 217271 167331 217277
rect 178310 217268 178316 217280
rect 178368 217268 178374 217320
rect 181441 217311 181499 217317
rect 181441 217277 181453 217311
rect 181487 217308 181499 217311
rect 192202 217308 192208 217320
rect 181487 217280 192208 217308
rect 181487 217277 181499 217280
rect 181441 217271 181499 217277
rect 192202 217268 192208 217280
rect 192260 217268 192266 217320
rect 192478 217268 192484 217320
rect 192536 217308 192542 217320
rect 199562 217308 199568 217320
rect 192536 217280 199568 217308
rect 192536 217268 192542 217280
rect 199562 217268 199568 217280
rect 199620 217268 199626 217320
rect 201402 217268 201408 217320
rect 201460 217308 201466 217320
rect 238754 217308 238760 217320
rect 201460 217280 238760 217308
rect 201460 217268 201466 217280
rect 238754 217268 238760 217280
rect 238812 217268 238818 217320
rect 241422 217268 241428 217320
rect 241480 217308 241486 217320
rect 252646 217308 252652 217320
rect 241480 217280 252652 217308
rect 241480 217268 241486 217280
rect 252646 217268 252652 217280
rect 252704 217268 252710 217320
rect 265250 217268 265256 217320
rect 265308 217308 265314 217320
rect 276658 217308 276664 217320
rect 265308 217280 276664 217308
rect 265308 217268 265314 217280
rect 276658 217268 276664 217280
rect 276716 217268 276722 217320
rect 280798 217268 280804 217320
rect 280856 217308 280862 217320
rect 280856 217280 287744 217308
rect 280856 217268 280862 217280
rect 84838 217200 84844 217252
rect 84896 217240 84902 217252
rect 189718 217240 189724 217252
rect 84896 217212 189724 217240
rect 84896 217200 84902 217212
rect 189718 217200 189724 217212
rect 189776 217200 189782 217252
rect 192570 217200 192576 217252
rect 192628 217240 192634 217252
rect 198366 217240 198372 217252
rect 192628 217212 198372 217240
rect 192628 217200 192634 217212
rect 198366 217200 198372 217212
rect 198424 217200 198430 217252
rect 219342 217200 219348 217252
rect 219400 217240 219406 217252
rect 245286 217240 245292 217252
rect 219400 217212 245292 217240
rect 219400 217200 219406 217212
rect 245286 217200 245292 217212
rect 245344 217200 245350 217252
rect 278774 217200 278780 217252
rect 278832 217240 278838 217252
rect 283650 217240 283656 217252
rect 278832 217212 283656 217240
rect 278832 217200 278838 217212
rect 283650 217200 283656 217212
rect 283708 217200 283714 217252
rect 285674 217200 285680 217252
rect 285732 217240 285738 217252
rect 286870 217240 286876 217252
rect 285732 217212 286876 217240
rect 285732 217200 285738 217212
rect 286870 217200 286876 217212
rect 286928 217200 286934 217252
rect 287716 217240 287744 217280
rect 288526 217268 288532 217320
rect 288584 217308 288590 217320
rect 289630 217308 289636 217320
rect 288584 217280 289636 217308
rect 288584 217268 288590 217280
rect 289630 217268 289636 217280
rect 289688 217268 289694 217320
rect 290182 217268 290188 217320
rect 290240 217308 290246 217320
rect 291102 217308 291108 217320
rect 290240 217280 291108 217308
rect 290240 217268 290246 217280
rect 291102 217268 291108 217280
rect 291160 217268 291166 217320
rect 291197 217311 291255 217317
rect 291197 217277 291209 217311
rect 291243 217308 291255 217311
rect 312538 217308 312544 217320
rect 291243 217280 312544 217308
rect 291243 217277 291255 217280
rect 291197 217271 291255 217277
rect 312538 217268 312544 217280
rect 312596 217268 312602 217320
rect 312648 217308 312676 217348
rect 313458 217336 313464 217388
rect 313516 217376 313522 217388
rect 327718 217376 327724 217388
rect 313516 217348 327724 217376
rect 313516 217336 313522 217348
rect 327718 217336 327724 217348
rect 327776 217336 327782 217388
rect 328178 217336 328184 217388
rect 328236 217376 328242 217388
rect 332413 217379 332471 217385
rect 332413 217376 332425 217379
rect 328236 217348 332425 217376
rect 328236 217336 328242 217348
rect 332413 217345 332425 217348
rect 332459 217345 332471 217379
rect 332520 217376 332548 217416
rect 332594 217404 332600 217456
rect 332652 217444 332658 217456
rect 333698 217444 333704 217456
rect 332652 217416 333704 217444
rect 332652 217404 332658 217416
rect 333698 217404 333704 217416
rect 333756 217404 333762 217456
rect 335357 217447 335415 217453
rect 335357 217413 335369 217447
rect 335403 217444 335415 217447
rect 336645 217447 336703 217453
rect 336645 217444 336657 217447
rect 335403 217416 336657 217444
rect 335403 217413 335415 217416
rect 335357 217407 335415 217413
rect 336645 217413 336657 217416
rect 336691 217413 336703 217447
rect 336645 217407 336703 217413
rect 337102 217404 337108 217456
rect 337160 217444 337166 217456
rect 338022 217444 338028 217456
rect 337160 217416 338028 217444
rect 337160 217404 337166 217416
rect 338022 217404 338028 217416
rect 338080 217404 338086 217456
rect 339497 217447 339555 217453
rect 339497 217444 339509 217447
rect 338132 217416 339509 217444
rect 338132 217376 338160 217416
rect 339497 217413 339509 217416
rect 339543 217413 339555 217447
rect 339497 217407 339555 217413
rect 339954 217404 339960 217456
rect 340012 217444 340018 217456
rect 340598 217444 340604 217456
rect 340012 217416 340604 217444
rect 340012 217404 340018 217416
rect 340598 217404 340604 217416
rect 340656 217404 340662 217456
rect 340693 217447 340751 217453
rect 340693 217413 340705 217447
rect 340739 217444 340751 217447
rect 456794 217444 456800 217456
rect 340739 217416 456800 217444
rect 340739 217413 340751 217416
rect 340693 217407 340751 217413
rect 456794 217404 456800 217416
rect 456852 217404 456858 217456
rect 332520 217348 338160 217376
rect 332413 217339 332471 217345
rect 338758 217336 338764 217388
rect 338816 217376 338822 217388
rect 339310 217376 339316 217388
rect 338816 217348 339316 217376
rect 338816 217336 338822 217348
rect 339310 217336 339316 217348
rect 339368 217336 339374 217388
rect 339405 217379 339463 217385
rect 339405 217345 339417 217379
rect 339451 217376 339463 217379
rect 340785 217379 340843 217385
rect 339451 217348 340644 217376
rect 339451 217345 339463 217348
rect 339405 217339 339463 217345
rect 326338 217308 326344 217320
rect 312648 217280 326344 217308
rect 326338 217268 326344 217280
rect 326396 217268 326402 217320
rect 326890 217268 326896 217320
rect 326948 217308 326954 217320
rect 340509 217311 340567 217317
rect 340509 217308 340521 217311
rect 326948 217280 340521 217308
rect 326948 217268 326954 217280
rect 340509 217277 340521 217280
rect 340555 217277 340567 217311
rect 340616 217308 340644 217348
rect 340785 217345 340797 217379
rect 340831 217376 340843 217379
rect 463694 217376 463700 217388
rect 340831 217348 463700 217376
rect 340831 217345 340843 217348
rect 340785 217339 340843 217345
rect 463694 217336 463700 217348
rect 463752 217336 463758 217388
rect 477494 217308 477500 217320
rect 340616 217280 477500 217308
rect 340509 217271 340567 217277
rect 477494 217268 477500 217280
rect 477552 217268 477558 217320
rect 305730 217240 305736 217252
rect 287716 217212 305736 217240
rect 305730 217200 305736 217212
rect 305788 217200 305794 217252
rect 313826 217200 313832 217252
rect 313884 217240 313890 217252
rect 314562 217240 314568 217252
rect 313884 217212 314568 217240
rect 313884 217200 313890 217212
rect 314562 217200 314568 217212
rect 314620 217200 314626 217252
rect 319901 217243 319959 217249
rect 319901 217240 319913 217243
rect 314672 217212 319913 217240
rect 95878 217132 95884 217184
rect 95936 217172 95942 217184
rect 200758 217172 200764 217184
rect 95936 217144 200764 217172
rect 95936 217132 95942 217144
rect 200758 217132 200764 217144
rect 200816 217132 200822 217184
rect 226242 217132 226248 217184
rect 226300 217172 226306 217184
rect 247310 217172 247316 217184
rect 226300 217144 247316 217172
rect 226300 217132 226306 217144
rect 247310 217132 247316 217144
rect 247368 217132 247374 217184
rect 275094 217132 275100 217184
rect 275152 217172 275158 217184
rect 281813 217175 281871 217181
rect 281813 217172 281825 217175
rect 275152 217144 281825 217172
rect 275152 217132 275158 217144
rect 281813 217141 281825 217144
rect 281859 217141 281871 217175
rect 281813 217135 281871 217141
rect 281920 217144 296392 217172
rect 104802 217064 104808 217116
rect 104860 217104 104866 217116
rect 205634 217104 205640 217116
rect 104860 217076 205640 217104
rect 104860 217064 104866 217076
rect 205634 217064 205640 217076
rect 205692 217064 205698 217116
rect 227622 217064 227628 217116
rect 227680 217104 227686 217116
rect 247678 217104 247684 217116
rect 227680 217076 247684 217104
rect 227680 217064 227686 217076
rect 247678 217064 247684 217076
rect 247736 217064 247742 217116
rect 261202 217064 261208 217116
rect 261260 217104 261266 217116
rect 261260 217076 263548 217104
rect 261260 217064 261266 217076
rect 102778 216996 102784 217048
rect 102836 217036 102842 217048
rect 203242 217036 203248 217048
rect 102836 217008 203248 217036
rect 102836 216996 102842 217008
rect 203242 216996 203248 217008
rect 203300 216996 203306 217048
rect 230382 216996 230388 217048
rect 230440 217036 230446 217048
rect 248966 217036 248972 217048
rect 230440 217008 248972 217036
rect 230440 216996 230446 217008
rect 248966 216996 248972 217008
rect 249024 216996 249030 217048
rect 249334 216996 249340 217048
rect 249392 217036 249398 217048
rect 253014 217036 253020 217048
rect 249392 217008 253020 217036
rect 249392 216996 249398 217008
rect 253014 216996 253020 217008
rect 253072 216996 253078 217048
rect 262398 216996 262404 217048
rect 262456 217036 262462 217048
rect 263410 217036 263416 217048
rect 262456 217008 263416 217036
rect 262456 216996 262462 217008
rect 263410 216996 263416 217008
rect 263468 216996 263474 217048
rect 263520 217036 263548 217076
rect 274634 217064 274640 217116
rect 274692 217104 274698 217116
rect 281920 217104 281948 217144
rect 274692 217076 281948 217104
rect 281997 217107 282055 217113
rect 274692 217064 274698 217076
rect 281997 217073 282009 217107
rect 282043 217104 282055 217107
rect 282043 217076 292988 217104
rect 282043 217073 282055 217076
rect 281997 217067 282055 217073
rect 265250 217036 265256 217048
rect 263520 217008 265256 217036
rect 265250 216996 265256 217008
rect 265308 216996 265314 217048
rect 266538 216996 266544 217048
rect 266596 217036 266602 217048
rect 267642 217036 267648 217048
rect 266596 217008 267648 217036
rect 266596 216996 266602 217008
rect 267642 216996 267648 217008
rect 267700 216996 267706 217048
rect 272242 216996 272248 217048
rect 272300 217036 272306 217048
rect 272300 217008 286548 217036
rect 272300 216996 272306 217008
rect 111702 216928 111708 216980
rect 111760 216968 111766 216980
rect 208118 216968 208124 216980
rect 111760 216940 208124 216968
rect 111760 216928 111766 216940
rect 208118 216928 208124 216940
rect 208176 216928 208182 216980
rect 229738 216928 229744 216980
rect 229796 216968 229802 216980
rect 246482 216968 246488 216980
rect 229796 216940 246488 216968
rect 229796 216928 229802 216940
rect 246482 216928 246488 216940
rect 246540 216928 246546 216980
rect 252462 216928 252468 216980
rect 252520 216968 252526 216980
rect 256326 216968 256332 216980
rect 252520 216940 256332 216968
rect 252520 216928 252526 216940
rect 256326 216928 256332 216940
rect 256384 216928 256390 216980
rect 270954 216928 270960 216980
rect 271012 216968 271018 216980
rect 283558 216968 283564 216980
rect 271012 216940 283564 216968
rect 271012 216928 271018 216940
rect 283558 216928 283564 216940
rect 283616 216928 283622 216980
rect 286520 216968 286548 217008
rect 287330 216996 287336 217048
rect 287388 217036 287394 217048
rect 288250 217036 288256 217048
rect 287388 217008 288256 217036
rect 287388 216996 287394 217008
rect 288250 216996 288256 217008
rect 288308 216996 288314 217048
rect 290458 216968 290464 216980
rect 286520 216940 290464 216968
rect 290458 216928 290464 216940
rect 290516 216928 290522 216980
rect 292960 216968 292988 217076
rect 293034 217064 293040 217116
rect 293092 217104 293098 217116
rect 293770 217104 293776 217116
rect 293092 217076 293776 217104
rect 293092 217064 293098 217076
rect 293770 217064 293776 217076
rect 293828 217064 293834 217116
rect 296364 217104 296392 217144
rect 297082 217132 297088 217184
rect 297140 217172 297146 217184
rect 297818 217172 297824 217184
rect 297140 217144 297824 217172
rect 297140 217132 297146 217144
rect 297818 217132 297824 217144
rect 297876 217132 297882 217184
rect 300118 217172 300124 217184
rect 297928 217144 300124 217172
rect 297928 217104 297956 217144
rect 300118 217132 300124 217144
rect 300176 217132 300182 217184
rect 310054 217132 310060 217184
rect 310112 217172 310118 217184
rect 314672 217172 314700 217212
rect 319901 217209 319913 217212
rect 319947 217209 319959 217243
rect 319901 217203 319959 217209
rect 319993 217243 320051 217249
rect 319993 217209 320005 217243
rect 320039 217240 320051 217243
rect 427814 217240 427820 217252
rect 320039 217212 427820 217240
rect 320039 217209 320051 217212
rect 319993 217203 320051 217209
rect 427814 217200 427820 217212
rect 427872 217200 427878 217252
rect 310112 217144 314700 217172
rect 310112 217132 310118 217144
rect 314838 217132 314844 217184
rect 314896 217172 314902 217184
rect 420914 217172 420920 217184
rect 314896 217144 420920 217172
rect 314896 217132 314902 217144
rect 420914 217132 420920 217144
rect 420972 217132 420978 217184
rect 296364 217076 297956 217104
rect 298370 217064 298376 217116
rect 298428 217104 298434 217116
rect 299290 217104 299296 217116
rect 298428 217076 299296 217104
rect 298428 217064 298434 217076
rect 299290 217064 299296 217076
rect 299348 217064 299354 217116
rect 302145 217107 302203 217113
rect 302145 217073 302157 217107
rect 302191 217104 302203 217107
rect 316678 217104 316684 217116
rect 302191 217076 316684 217104
rect 302191 217073 302203 217076
rect 302145 217067 302203 217073
rect 316678 217064 316684 217076
rect 316736 217064 316742 217116
rect 414014 217104 414020 217116
rect 317432 217076 414020 217104
rect 294230 216996 294236 217048
rect 294288 217036 294294 217048
rect 295242 217036 295248 217048
rect 294288 217008 295248 217036
rect 294288 216996 294294 217008
rect 295242 216996 295248 217008
rect 295300 216996 295306 217048
rect 295337 217039 295395 217045
rect 295337 217005 295349 217039
rect 295383 217036 295395 217039
rect 295383 217008 297496 217036
rect 295383 217005 295395 217008
rect 295337 216999 295395 217005
rect 297358 216968 297364 216980
rect 292960 216940 297364 216968
rect 297358 216928 297364 216940
rect 297416 216928 297422 216980
rect 297468 216968 297496 217008
rect 302418 216996 302424 217048
rect 302476 217036 302482 217048
rect 307205 217039 307263 217045
rect 307205 217036 307217 217039
rect 302476 217008 307217 217036
rect 302476 216996 302482 217008
rect 307205 217005 307217 217008
rect 307251 217005 307263 217039
rect 307205 216999 307263 217005
rect 307294 216996 307300 217048
rect 307352 217036 307358 217048
rect 307352 217008 312032 217036
rect 307352 216996 307358 217008
rect 305638 216968 305644 216980
rect 297468 216940 305644 216968
rect 305638 216928 305644 216940
rect 305696 216928 305702 216980
rect 308582 216928 308588 216980
rect 308640 216968 308646 216980
rect 311897 216971 311955 216977
rect 311897 216968 311909 216971
rect 308640 216940 311909 216968
rect 308640 216928 308646 216940
rect 311897 216937 311909 216940
rect 311943 216937 311955 216971
rect 312004 216968 312032 217008
rect 312170 216996 312176 217048
rect 312228 217036 312234 217048
rect 317432 217036 317460 217076
rect 414014 217064 414020 217076
rect 414072 217064 414078 217116
rect 312228 217008 317460 217036
rect 312228 216996 312234 217008
rect 318150 216996 318156 217048
rect 318208 217036 318214 217048
rect 318518 217036 318524 217048
rect 318208 217008 318524 217036
rect 318208 216996 318214 217008
rect 318518 216996 318524 217008
rect 318576 216996 318582 217048
rect 319901 217039 319959 217045
rect 319901 217005 319913 217039
rect 319947 217036 319959 217039
rect 407114 217036 407120 217048
rect 319947 217008 407120 217036
rect 319947 217005 319959 217008
rect 319901 216999 319959 217005
rect 407114 216996 407120 217008
rect 407172 216996 407178 217048
rect 400214 216968 400220 216980
rect 312004 216940 400220 216968
rect 311897 216931 311955 216937
rect 400214 216928 400220 216940
rect 400272 216928 400278 216980
rect 118602 216860 118608 216912
rect 118660 216900 118666 216912
rect 210602 216900 210608 216912
rect 118660 216872 210608 216900
rect 118660 216860 118666 216872
rect 210602 216860 210608 216872
rect 210660 216860 210666 216912
rect 237282 216860 237288 216912
rect 237340 216900 237346 216912
rect 251358 216900 251364 216912
rect 237340 216872 251364 216900
rect 237340 216860 237346 216872
rect 251358 216860 251364 216872
rect 251416 216860 251422 216912
rect 251910 216860 251916 216912
rect 251968 216900 251974 216912
rect 255498 216900 255504 216912
rect 251968 216872 255504 216900
rect 251968 216860 251974 216872
rect 255498 216860 255504 216872
rect 255556 216860 255562 216912
rect 263686 216860 263692 216912
rect 263744 216900 263750 216912
rect 269758 216900 269764 216912
rect 263744 216872 269764 216900
rect 263744 216860 263750 216872
rect 269758 216860 269764 216872
rect 269816 216860 269822 216912
rect 273438 216860 273444 216912
rect 273496 216900 273502 216912
rect 281997 216903 282055 216909
rect 281997 216900 282009 216903
rect 273496 216872 282009 216900
rect 273496 216860 273502 216872
rect 281997 216869 282009 216872
rect 282043 216869 282055 216903
rect 281997 216863 282055 216869
rect 282822 216860 282828 216912
rect 282880 216900 282886 216912
rect 289817 216903 289875 216909
rect 289817 216900 289829 216903
rect 282880 216872 289829 216900
rect 282880 216860 282886 216872
rect 289817 216869 289829 216872
rect 289863 216869 289875 216903
rect 289817 216863 289875 216869
rect 304902 216860 304908 216912
rect 304960 216900 304966 216912
rect 308401 216903 308459 216909
rect 308401 216900 308413 216903
rect 304960 216872 308413 216900
rect 304960 216860 304966 216872
rect 308401 216869 308413 216872
rect 308447 216869 308459 216903
rect 308401 216863 308459 216869
rect 308677 216903 308735 216909
rect 308677 216869 308689 216903
rect 308723 216900 308735 216903
rect 391934 216900 391940 216912
rect 308723 216872 391940 216900
rect 308723 216869 308735 216872
rect 308677 216863 308735 216869
rect 391934 216860 391940 216872
rect 391992 216860 391998 216912
rect 122742 216792 122748 216844
rect 122800 216832 122806 216844
rect 211522 216832 211528 216844
rect 122800 216804 211528 216832
rect 122800 216792 122806 216804
rect 211522 216792 211528 216804
rect 211580 216792 211586 216844
rect 232498 216792 232504 216844
rect 232556 216832 232562 216844
rect 241974 216832 241980 216844
rect 232556 216804 241980 216832
rect 232556 216792 232562 216804
rect 241974 216792 241980 216804
rect 242032 216792 242038 216844
rect 243538 216792 243544 216844
rect 243596 216832 243602 216844
rect 246942 216832 246948 216844
rect 243596 216804 246948 216832
rect 243596 216792 243602 216804
rect 246942 216792 246948 216804
rect 247000 216792 247006 216844
rect 250898 216792 250904 216844
rect 250956 216832 250962 216844
rect 254210 216832 254216 216844
rect 250956 216804 254216 216832
rect 250956 216792 250962 216804
rect 254210 216792 254216 216804
rect 254268 216792 254274 216844
rect 254578 216792 254584 216844
rect 254636 216832 254642 216844
rect 256694 216832 256700 216844
rect 254636 216804 256700 216832
rect 254636 216792 254642 216804
rect 256694 216792 256700 216804
rect 256752 216792 256758 216844
rect 271414 216792 271420 216844
rect 271472 216832 271478 216844
rect 273898 216832 273904 216844
rect 271472 216804 273904 216832
rect 271472 216792 271478 216804
rect 273898 216792 273904 216804
rect 273956 216792 273962 216844
rect 283101 216835 283159 216841
rect 283101 216801 283113 216835
rect 283147 216832 283159 216835
rect 291933 216835 291991 216841
rect 291933 216832 291945 216835
rect 283147 216804 291945 216832
rect 283147 216801 283159 216804
rect 283101 216795 283159 216801
rect 291933 216801 291945 216804
rect 291979 216801 291991 216835
rect 291933 216795 291991 216801
rect 299385 216835 299443 216841
rect 299385 216801 299397 216835
rect 299431 216832 299443 216835
rect 302145 216835 302203 216841
rect 302145 216832 302157 216835
rect 299431 216804 302157 216832
rect 299431 216801 299443 216804
rect 299385 216795 299443 216801
rect 302145 216801 302157 216804
rect 302191 216801 302203 216835
rect 302145 216795 302203 216801
rect 307205 216835 307263 216841
rect 307205 216801 307217 216835
rect 307251 216832 307263 216835
rect 385034 216832 385040 216844
rect 307251 216804 385040 216832
rect 307251 216801 307263 216804
rect 307205 216795 307263 216801
rect 385034 216792 385040 216804
rect 385092 216792 385098 216844
rect 97258 216724 97264 216776
rect 97316 216764 97322 216776
rect 186130 216764 186136 216776
rect 97316 216736 186136 216764
rect 97316 216724 97322 216736
rect 186130 216724 186136 216736
rect 186188 216724 186194 216776
rect 244918 216724 244924 216776
rect 244976 216764 244982 216776
rect 248138 216764 248144 216776
rect 244976 216736 248144 216764
rect 244976 216724 244982 216736
rect 248138 216724 248144 216736
rect 248196 216724 248202 216776
rect 250806 216724 250812 216776
rect 250864 216764 250870 216776
rect 252186 216764 252192 216776
rect 250864 216736 252192 216764
rect 250864 216724 250870 216736
rect 252186 216724 252192 216736
rect 252244 216724 252250 216776
rect 282917 216767 282975 216773
rect 282917 216733 282929 216767
rect 282963 216764 282975 216767
rect 291197 216767 291255 216773
rect 291197 216764 291209 216767
rect 282963 216736 291209 216764
rect 282963 216733 282975 216736
rect 282917 216727 282975 216733
rect 291197 216733 291209 216736
rect 291243 216733 291255 216767
rect 291197 216727 291255 216733
rect 291838 216724 291844 216776
rect 291896 216764 291902 216776
rect 292390 216764 292396 216776
rect 291896 216736 292396 216764
rect 291896 216724 291902 216736
rect 292390 216724 292396 216736
rect 292448 216724 292454 216776
rect 302786 216724 302792 216776
rect 302844 216764 302850 216776
rect 303522 216764 303528 216776
rect 302844 216736 303528 216764
rect 302844 216724 302850 216736
rect 303522 216724 303528 216736
rect 303580 216724 303586 216776
rect 304074 216724 304080 216776
rect 304132 216764 304138 216776
rect 304902 216764 304908 216776
rect 304132 216736 304908 216764
rect 304132 216724 304138 216736
rect 304902 216724 304908 216736
rect 304960 216724 304966 216776
rect 305270 216724 305276 216776
rect 305328 216764 305334 216776
rect 306190 216764 306196 216776
rect 305328 216736 306196 216764
rect 305328 216724 305334 216736
rect 306190 216724 306196 216736
rect 306248 216724 306254 216776
rect 306466 216724 306472 216776
rect 306524 216764 306530 216776
rect 307570 216764 307576 216776
rect 306524 216736 307576 216764
rect 306524 216724 306530 216736
rect 307570 216724 307576 216736
rect 307628 216724 307634 216776
rect 307754 216724 307760 216776
rect 307812 216764 307818 216776
rect 308858 216764 308864 216776
rect 307812 216736 308864 216764
rect 307812 216724 307818 216736
rect 308858 216724 308864 216736
rect 308916 216724 308922 216776
rect 311434 216724 311440 216776
rect 311492 216764 311498 216776
rect 311802 216764 311808 216776
rect 311492 216736 311808 216764
rect 311492 216724 311498 216736
rect 311802 216724 311808 216736
rect 311860 216724 311866 216776
rect 311897 216767 311955 216773
rect 311897 216733 311909 216767
rect 311943 216764 311955 216767
rect 311943 216736 321508 216764
rect 311943 216733 311955 216736
rect 311897 216727 311955 216733
rect 106918 216656 106924 216708
rect 106976 216696 106982 216708
rect 181441 216699 181499 216705
rect 181441 216696 181453 216699
rect 106976 216668 181453 216696
rect 106976 216656 106982 216668
rect 181441 216665 181453 216668
rect 181487 216665 181499 216699
rect 181441 216659 181499 216665
rect 185578 216656 185584 216708
rect 185636 216696 185642 216708
rect 188522 216696 188528 216708
rect 185636 216668 188528 216696
rect 185636 216656 185642 216668
rect 188522 216656 188528 216668
rect 188580 216656 188586 216708
rect 211798 216656 211804 216708
rect 211856 216696 211862 216708
rect 212258 216696 212264 216708
rect 211856 216668 212264 216696
rect 211856 216656 211862 216668
rect 212258 216656 212264 216668
rect 212316 216656 212322 216708
rect 239398 216656 239404 216708
rect 239456 216696 239462 216708
rect 244826 216696 244832 216708
rect 239456 216668 244832 216696
rect 239456 216656 239462 216668
rect 244826 216656 244832 216668
rect 244884 216656 244890 216708
rect 245010 216656 245016 216708
rect 245068 216696 245074 216708
rect 246114 216696 246120 216708
rect 245068 216668 246120 216696
rect 245068 216656 245074 216668
rect 246114 216656 246120 216668
rect 246172 216656 246178 216708
rect 247678 216656 247684 216708
rect 247736 216696 247742 216708
rect 248506 216696 248512 216708
rect 247736 216668 248512 216696
rect 247736 216656 247742 216668
rect 248506 216656 248512 216668
rect 248564 216656 248570 216708
rect 249150 216656 249156 216708
rect 249208 216696 249214 216708
rect 249794 216696 249800 216708
rect 249208 216668 249800 216696
rect 249208 216656 249214 216668
rect 249794 216656 249800 216668
rect 249852 216656 249858 216708
rect 251818 216656 251824 216708
rect 251876 216696 251882 216708
rect 253474 216696 253480 216708
rect 251876 216668 253480 216696
rect 251876 216656 251882 216668
rect 253474 216656 253480 216668
rect 253532 216656 253538 216708
rect 289817 216699 289875 216705
rect 289817 216665 289829 216699
rect 289863 216696 289875 216699
rect 299385 216699 299443 216705
rect 299385 216696 299397 216699
rect 289863 216668 299397 216696
rect 289863 216665 289875 216668
rect 289817 216659 289875 216665
rect 299385 216665 299397 216668
rect 299431 216665 299443 216699
rect 299385 216659 299443 216665
rect 306926 216656 306932 216708
rect 306984 216696 306990 216708
rect 307662 216696 307668 216708
rect 306984 216668 307668 216696
rect 306984 216656 306990 216668
rect 307662 216656 307668 216668
rect 307720 216656 307726 216708
rect 308122 216656 308128 216708
rect 308180 216696 308186 216708
rect 308950 216696 308956 216708
rect 308180 216668 308956 216696
rect 308180 216656 308186 216668
rect 308950 216656 308956 216668
rect 309008 216656 309014 216708
rect 309318 216656 309324 216708
rect 309376 216696 309382 216708
rect 310330 216696 310336 216708
rect 309376 216668 310336 216696
rect 309376 216656 309382 216668
rect 310330 216656 310336 216668
rect 310388 216656 310394 216708
rect 310606 216656 310612 216708
rect 310664 216696 310670 216708
rect 311618 216696 311624 216708
rect 310664 216668 311624 216696
rect 310664 216656 310670 216668
rect 311618 216656 311624 216668
rect 311676 216656 311682 216708
rect 312630 216656 312636 216708
rect 312688 216696 312694 216708
rect 313182 216696 313188 216708
rect 312688 216668 313188 216696
rect 312688 216656 312694 216668
rect 313182 216656 313188 216668
rect 313240 216656 313246 216708
rect 315114 216656 315120 216708
rect 315172 216696 315178 216708
rect 315942 216696 315948 216708
rect 315172 216668 315948 216696
rect 315172 216656 315178 216668
rect 315942 216656 315948 216668
rect 316000 216656 316006 216708
rect 316310 216656 316316 216708
rect 316368 216696 316374 216708
rect 317322 216696 317328 216708
rect 316368 216668 317328 216696
rect 316368 216656 316374 216668
rect 317322 216656 317328 216668
rect 317380 216656 317386 216708
rect 317506 216656 317512 216708
rect 317564 216696 317570 216708
rect 318610 216696 318616 216708
rect 317564 216668 318616 216696
rect 317564 216656 317570 216668
rect 318610 216656 318616 216668
rect 318668 216656 318674 216708
rect 319162 216656 319168 216708
rect 319220 216696 319226 216708
rect 319990 216696 319996 216708
rect 319220 216668 319996 216696
rect 319220 216656 319226 216668
rect 319990 216656 319996 216668
rect 320048 216656 320054 216708
rect 320358 216656 320364 216708
rect 320416 216696 320422 216708
rect 321370 216696 321376 216708
rect 320416 216668 321376 216696
rect 320416 216656 320422 216668
rect 321370 216656 321376 216668
rect 321428 216656 321434 216708
rect 321480 216696 321508 216736
rect 322014 216724 322020 216776
rect 322072 216764 322078 216776
rect 322072 216736 330524 216764
rect 322072 216724 322078 216736
rect 323578 216696 323584 216708
rect 321480 216668 323584 216696
rect 323578 216656 323584 216668
rect 323636 216656 323642 216708
rect 325694 216656 325700 216708
rect 325752 216696 325758 216708
rect 330496 216696 330524 216736
rect 330570 216724 330576 216776
rect 330628 216764 330634 216776
rect 337378 216764 337384 216776
rect 330628 216736 337384 216764
rect 330628 216724 330634 216736
rect 337378 216724 337384 216736
rect 337436 216724 337442 216776
rect 339586 216724 339592 216776
rect 339644 216764 339650 216776
rect 340782 216764 340788 216776
rect 339644 216736 340788 216764
rect 339644 216724 339650 216736
rect 340782 216724 340788 216736
rect 340840 216724 340846 216776
rect 341058 216724 341064 216776
rect 341116 216764 341122 216776
rect 341518 216764 341524 216776
rect 341116 216736 341524 216764
rect 341116 216724 341122 216736
rect 341518 216724 341524 216736
rect 341576 216724 341582 216776
rect 343634 216724 343640 216776
rect 343692 216764 343698 216776
rect 344738 216764 344744 216776
rect 343692 216736 344744 216764
rect 343692 216724 343698 216736
rect 344738 216724 344744 216736
rect 344796 216724 344802 216776
rect 361206 216724 361212 216776
rect 361264 216764 361270 216776
rect 369765 216767 369823 216773
rect 369765 216764 369777 216767
rect 361264 216736 369777 216764
rect 361264 216724 361270 216736
rect 369765 216733 369777 216736
rect 369811 216733 369823 216767
rect 369765 216727 369823 216733
rect 331125 216699 331183 216705
rect 331125 216696 331137 216699
rect 325752 216668 330432 216696
rect 330496 216668 331137 216696
rect 325752 216656 325758 216668
rect 330404 216560 330432 216668
rect 331125 216665 331137 216668
rect 331171 216665 331183 216699
rect 345658 216696 345664 216708
rect 331125 216659 331183 216665
rect 331232 216668 345664 216696
rect 331232 216560 331260 216668
rect 345658 216656 345664 216668
rect 345716 216656 345722 216708
rect 330404 216532 331260 216560
rect 194686 216316 194692 216368
rect 194744 216356 194750 216368
rect 195514 216356 195520 216368
rect 194744 216328 195520 216356
rect 194744 216316 194750 216328
rect 195514 216316 195520 216328
rect 195572 216316 195578 216368
rect 219802 215704 219808 215756
rect 219860 215744 219866 215756
rect 220354 215744 220360 215756
rect 219860 215716 220360 215744
rect 219860 215704 219866 215716
rect 220354 215704 220360 215716
rect 220412 215704 220418 215756
rect 216858 215568 216864 215620
rect 216916 215608 216922 215620
rect 217502 215608 217508 215620
rect 216916 215580 217508 215608
rect 216916 215568 216922 215580
rect 217502 215568 217508 215580
rect 217560 215568 217566 215620
rect 173986 215296 173992 215348
rect 174044 215336 174050 215348
rect 174630 215336 174636 215348
rect 174044 215308 174636 215336
rect 174044 215296 174050 215308
rect 174630 215296 174636 215308
rect 174688 215296 174694 215348
rect 209866 215296 209872 215348
rect 209924 215336 209930 215348
rect 210786 215336 210792 215348
rect 209924 215308 210792 215336
rect 209924 215296 209930 215308
rect 210786 215296 210792 215308
rect 210844 215296 210850 215348
rect 216953 215339 217011 215345
rect 216953 215305 216965 215339
rect 216999 215336 217011 215339
rect 217134 215336 217140 215348
rect 216999 215308 217140 215336
rect 216999 215305 217011 215308
rect 216953 215299 217011 215305
rect 217134 215296 217140 215308
rect 217192 215296 217198 215348
rect 291930 215200 291936 215212
rect 291891 215172 291936 215200
rect 291930 215160 291936 215172
rect 291988 215160 291994 215212
rect 205726 214548 205732 214600
rect 205784 214588 205790 214600
rect 206186 214588 206192 214600
rect 205784 214560 206192 214588
rect 205784 214548 205790 214560
rect 206186 214548 206192 214560
rect 206244 214548 206250 214600
rect 208486 214548 208492 214600
rect 208544 214588 208550 214600
rect 208670 214588 208676 214600
rect 208544 214560 208676 214588
rect 208544 214548 208550 214560
rect 208670 214548 208676 214560
rect 208728 214548 208734 214600
rect 212810 214548 212816 214600
rect 212868 214588 212874 214600
rect 213546 214588 213552 214600
rect 212868 214560 213552 214588
rect 212868 214548 212874 214560
rect 213546 214548 213552 214560
rect 213604 214548 213610 214600
rect 214006 214548 214012 214600
rect 214064 214588 214070 214600
rect 214742 214588 214748 214600
rect 214064 214560 214748 214588
rect 214064 214548 214070 214560
rect 214742 214548 214748 214560
rect 214800 214548 214806 214600
rect 333330 214548 333336 214600
rect 333388 214588 333394 214600
rect 333882 214588 333888 214600
rect 333388 214560 333888 214588
rect 333388 214548 333394 214560
rect 333882 214548 333888 214560
rect 333940 214548 333946 214600
rect 179414 213800 179420 213852
rect 179472 213840 179478 213852
rect 179966 213840 179972 213852
rect 179472 213812 179972 213840
rect 179472 213800 179478 213812
rect 179966 213800 179972 213812
rect 180024 213800 180030 213852
rect 193858 212848 193864 212900
rect 193916 212888 193922 212900
rect 202046 212888 202052 212900
rect 193916 212860 202052 212888
rect 193916 212848 193922 212860
rect 202046 212848 202052 212860
rect 202104 212848 202110 212900
rect 171410 212508 171416 212560
rect 171468 212548 171474 212560
rect 171778 212548 171784 212560
rect 171468 212520 171784 212548
rect 171468 212508 171474 212520
rect 171778 212508 171784 212520
rect 171836 212508 171842 212560
rect 173250 212508 173256 212560
rect 173308 212548 173314 212560
rect 173802 212548 173808 212560
rect 173308 212520 173808 212548
rect 173308 212508 173314 212520
rect 173802 212508 173808 212520
rect 173860 212508 173866 212560
rect 177298 212508 177304 212560
rect 177356 212548 177362 212560
rect 177942 212548 177948 212560
rect 177356 212520 177948 212548
rect 177356 212508 177362 212520
rect 177942 212508 177948 212520
rect 178000 212508 178006 212560
rect 178862 212508 178868 212560
rect 178920 212548 178926 212560
rect 179138 212548 179144 212560
rect 178920 212520 179144 212548
rect 178920 212508 178926 212520
rect 179138 212508 179144 212520
rect 179196 212508 179202 212560
rect 180150 212548 180156 212560
rect 180111 212520 180156 212548
rect 180150 212508 180156 212520
rect 180208 212508 180214 212560
rect 184014 212508 184020 212560
rect 184072 212548 184078 212560
rect 184474 212548 184480 212560
rect 184072 212520 184480 212548
rect 184072 212508 184078 212520
rect 184474 212508 184480 212520
rect 184532 212508 184538 212560
rect 189350 212508 189356 212560
rect 189408 212548 189414 212560
rect 190178 212548 190184 212560
rect 189408 212520 190184 212548
rect 189408 212508 189414 212520
rect 190178 212508 190184 212520
rect 190236 212508 190242 212560
rect 192386 212508 192392 212560
rect 192444 212548 192450 212560
rect 192662 212548 192668 212560
rect 192444 212520 192668 212548
rect 192444 212508 192450 212520
rect 192662 212508 192668 212520
rect 192720 212508 192726 212560
rect 200850 212508 200856 212560
rect 200908 212548 200914 212560
rect 201218 212548 201224 212560
rect 200908 212520 201224 212548
rect 200908 212508 200914 212520
rect 201218 212508 201224 212520
rect 201276 212508 201282 212560
rect 201862 212508 201868 212560
rect 201920 212548 201926 212560
rect 202414 212548 202420 212560
rect 201920 212520 202420 212548
rect 201920 212508 201926 212520
rect 202414 212508 202420 212520
rect 202472 212508 202478 212560
rect 203426 212508 203432 212560
rect 203484 212548 203490 212560
rect 203610 212548 203616 212560
rect 203484 212520 203616 212548
rect 203484 212508 203490 212520
rect 203610 212508 203616 212520
rect 203668 212508 203674 212560
rect 212350 212548 212356 212560
rect 212311 212520 212356 212548
rect 212350 212508 212356 212520
rect 212408 212508 212414 212560
rect 216950 212548 216956 212560
rect 216911 212520 216956 212548
rect 216950 212508 216956 212520
rect 217008 212508 217014 212560
rect 236270 212508 236276 212560
rect 236328 212548 236334 212560
rect 236730 212548 236736 212560
rect 236328 212520 236736 212548
rect 236328 212508 236334 212520
rect 236730 212508 236736 212520
rect 236788 212508 236794 212560
rect 283742 212508 283748 212560
rect 283800 212548 283806 212560
rect 284018 212548 284024 212560
rect 283800 212520 284024 212548
rect 283800 212508 283806 212520
rect 284018 212508 284024 212520
rect 284076 212508 284082 212560
rect 284846 212508 284852 212560
rect 284904 212548 284910 212560
rect 285306 212548 285312 212560
rect 284904 212520 285312 212548
rect 284904 212508 284910 212520
rect 285306 212508 285312 212520
rect 285364 212508 285370 212560
rect 286134 212508 286140 212560
rect 286192 212548 286198 212560
rect 286594 212548 286600 212560
rect 286192 212520 286600 212548
rect 286192 212508 286198 212520
rect 286594 212508 286600 212520
rect 286652 212508 286658 212560
rect 288986 212508 288992 212560
rect 289044 212548 289050 212560
rect 289354 212548 289360 212560
rect 289044 212520 289360 212548
rect 289044 212508 289050 212520
rect 289354 212508 289360 212520
rect 289412 212508 289418 212560
rect 294690 212508 294696 212560
rect 294748 212548 294754 212560
rect 295058 212548 295064 212560
rect 294748 212520 295064 212548
rect 294748 212508 294754 212520
rect 295058 212508 295064 212520
rect 295116 212508 295122 212560
rect 299934 212508 299940 212560
rect 299992 212548 299998 212560
rect 300486 212548 300492 212560
rect 299992 212520 300492 212548
rect 299992 212508 299998 212520
rect 300486 212508 300492 212520
rect 300544 212508 300550 212560
rect 360746 212508 360752 212560
rect 360804 212548 360810 212560
rect 361298 212548 361304 212560
rect 360804 212520 361304 212548
rect 360804 212508 360810 212520
rect 361298 212508 361304 212520
rect 361356 212508 361362 212560
rect 211890 212480 211896 212492
rect 211851 212452 211896 212480
rect 211890 212440 211896 212452
rect 211948 212440 211954 212492
rect 261938 211896 261944 211948
rect 261996 211936 262002 211948
rect 266538 211936 266544 211948
rect 261996 211908 266544 211936
rect 261996 211896 262002 211908
rect 266538 211896 266544 211908
rect 266596 211896 266602 211948
rect 260374 211216 260380 211268
rect 260432 211256 260438 211268
rect 262582 211256 262588 211268
rect 260432 211228 262588 211256
rect 260432 211216 260438 211228
rect 262582 211216 262588 211228
rect 262640 211216 262646 211268
rect 259546 211148 259552 211200
rect 259604 211188 259610 211200
rect 261110 211188 261116 211200
rect 259604 211160 261116 211188
rect 259604 211148 259610 211160
rect 261110 211148 261116 211160
rect 261168 211148 261174 211200
rect 217042 211120 217048 211132
rect 217003 211092 217048 211120
rect 217042 211080 217048 211092
rect 217100 211080 217106 211132
rect 262582 211120 262588 211132
rect 262543 211092 262588 211120
rect 262582 211080 262588 211092
rect 262640 211080 262646 211132
rect 266538 211080 266544 211132
rect 266596 211120 266602 211132
rect 266722 211120 266728 211132
rect 266596 211092 266728 211120
rect 266596 211080 266602 211092
rect 266722 211080 266728 211092
rect 266780 211080 266786 211132
rect 283834 211080 283840 211132
rect 283892 211120 283898 211132
rect 284018 211120 284024 211132
rect 283892 211092 284024 211120
rect 283892 211080 283898 211092
rect 284018 211080 284024 211092
rect 284076 211080 284082 211132
rect 328086 211120 328092 211132
rect 328047 211092 328092 211120
rect 328086 211080 328092 211092
rect 328144 211080 328150 211132
rect 341794 211080 341800 211132
rect 341852 211120 341858 211132
rect 341978 211120 341984 211132
rect 341852 211092 341984 211120
rect 341852 211080 341858 211092
rect 341978 211080 341984 211092
rect 342036 211080 342042 211132
rect 343266 211120 343272 211132
rect 343227 211092 343272 211120
rect 343266 211080 343272 211092
rect 343324 211080 343330 211132
rect 344554 211120 344560 211132
rect 344515 211092 344560 211120
rect 344554 211080 344560 211092
rect 344612 211080 344618 211132
rect 354122 211080 354128 211132
rect 354180 211120 354186 211132
rect 354214 211120 354220 211132
rect 354180 211092 354220 211120
rect 354180 211080 354186 211092
rect 354214 211080 354220 211092
rect 354272 211080 354278 211132
rect 355410 211080 355416 211132
rect 355468 211120 355474 211132
rect 355594 211120 355600 211132
rect 355468 211092 355600 211120
rect 355468 211080 355474 211092
rect 355594 211080 355600 211092
rect 355652 211080 355658 211132
rect 194686 210876 194692 210928
rect 194744 210916 194750 210928
rect 195146 210916 195152 210928
rect 194744 210888 195152 210916
rect 194744 210876 194750 210888
rect 195146 210876 195152 210888
rect 195204 210876 195210 210928
rect 169938 210468 169944 210520
rect 169996 210508 170002 210520
rect 170674 210508 170680 210520
rect 169996 210480 170680 210508
rect 169996 210468 170002 210480
rect 170674 210468 170680 210480
rect 170732 210468 170738 210520
rect 220906 210468 220912 210520
rect 220964 210508 220970 210520
rect 221734 210508 221740 210520
rect 220964 210480 221740 210508
rect 220964 210468 220970 210480
rect 221734 210468 221740 210480
rect 221792 210468 221798 210520
rect 169846 210400 169852 210452
rect 169904 210440 169910 210452
rect 170306 210440 170312 210452
rect 169904 210412 170312 210440
rect 169904 210400 169910 210412
rect 170306 210400 170312 210412
rect 170364 210400 170370 210452
rect 175366 210400 175372 210452
rect 175424 210440 175430 210452
rect 176010 210440 176016 210452
rect 175424 210412 176016 210440
rect 175424 210400 175430 210412
rect 176010 210400 176016 210412
rect 176068 210400 176074 210452
rect 179506 210400 179512 210452
rect 179564 210440 179570 210452
rect 180058 210440 180064 210452
rect 179564 210412 180064 210440
rect 179564 210400 179570 210412
rect 180058 210400 180064 210412
rect 180116 210400 180122 210452
rect 180886 210400 180892 210452
rect 180944 210440 180950 210452
rect 181254 210440 181260 210452
rect 180944 210412 181260 210440
rect 180944 210400 180950 210412
rect 181254 210400 181260 210412
rect 181312 210400 181318 210452
rect 186406 210400 186412 210452
rect 186464 210440 186470 210452
rect 186590 210440 186596 210452
rect 186464 210412 186596 210440
rect 186464 210400 186470 210412
rect 186590 210400 186596 210412
rect 186648 210400 186654 210452
rect 187970 210400 187976 210452
rect 188028 210440 188034 210452
rect 188614 210440 188620 210452
rect 188028 210412 188620 210440
rect 188028 210400 188034 210412
rect 188614 210400 188620 210412
rect 188672 210400 188678 210452
rect 192018 210400 192024 210452
rect 192076 210440 192082 210452
rect 192754 210440 192760 210452
rect 192076 210412 192760 210440
rect 192076 210400 192082 210412
rect 192754 210400 192760 210412
rect 192812 210400 192818 210452
rect 193306 210400 193312 210452
rect 193364 210440 193370 210452
rect 193950 210440 193956 210452
rect 193364 210412 193956 210440
rect 193364 210400 193370 210412
rect 193950 210400 193956 210412
rect 194008 210400 194014 210452
rect 201678 210400 201684 210452
rect 201736 210440 201742 210452
rect 202506 210440 202512 210452
rect 201736 210412 202512 210440
rect 201736 210400 201742 210412
rect 202506 210400 202512 210412
rect 202564 210400 202570 210452
rect 202966 210400 202972 210452
rect 203024 210440 203030 210452
rect 203702 210440 203708 210452
rect 203024 210412 203708 210440
rect 203024 210400 203030 210412
rect 203702 210400 203708 210412
rect 203760 210400 203766 210452
rect 204346 210400 204352 210452
rect 204404 210440 204410 210452
rect 204990 210440 204996 210452
rect 204404 210412 204996 210440
rect 204404 210400 204410 210412
rect 204990 210400 204996 210412
rect 205048 210400 205054 210452
rect 215386 210400 215392 210452
rect 215444 210440 215450 210452
rect 216030 210440 216036 210452
rect 215444 210412 216036 210440
rect 215444 210400 215450 210412
rect 216030 210400 216036 210412
rect 216088 210400 216094 210452
rect 218054 210400 218060 210452
rect 218112 210440 218118 210452
rect 218790 210440 218796 210452
rect 218112 210412 218796 210440
rect 218112 210400 218118 210412
rect 218790 210400 218796 210412
rect 218848 210400 218854 210452
rect 220998 210400 221004 210452
rect 221056 210440 221062 210452
rect 221366 210440 221372 210452
rect 221056 210412 221372 210440
rect 221056 210400 221062 210412
rect 221366 210400 221372 210412
rect 221424 210400 221430 210452
rect 222286 210400 222292 210452
rect 222344 210440 222350 210452
rect 222470 210440 222476 210452
rect 222344 210412 222476 210440
rect 222344 210400 222350 210412
rect 222470 210400 222476 210412
rect 222528 210400 222534 210452
rect 224954 210400 224960 210452
rect 225012 210440 225018 210452
rect 225782 210440 225788 210452
rect 225012 210412 225788 210440
rect 225012 210400 225018 210412
rect 225782 210400 225788 210412
rect 225840 210400 225846 210452
rect 226334 210400 226340 210452
rect 226392 210440 226398 210452
rect 227070 210440 227076 210452
rect 226392 210412 227076 210440
rect 226392 210400 226398 210412
rect 227070 210400 227076 210412
rect 227128 210400 227134 210452
rect 227898 210400 227904 210452
rect 227956 210440 227962 210452
rect 228634 210440 228640 210452
rect 227956 210412 228640 210440
rect 227956 210400 227962 210412
rect 228634 210400 228640 210412
rect 228692 210400 228698 210452
rect 229094 210400 229100 210452
rect 229152 210440 229158 210452
rect 229462 210440 229468 210452
rect 229152 210412 229468 210440
rect 229152 210400 229158 210412
rect 229462 210400 229468 210412
rect 229520 210400 229526 210452
rect 230474 210400 230480 210452
rect 230532 210440 230538 210452
rect 231118 210440 231124 210452
rect 230532 210412 231124 210440
rect 230532 210400 230538 210412
rect 231118 210400 231124 210412
rect 231176 210400 231182 210452
rect 231854 210400 231860 210452
rect 231912 210440 231918 210452
rect 232774 210440 232780 210452
rect 231912 210412 232780 210440
rect 231912 210400 231918 210412
rect 232774 210400 232780 210412
rect 232832 210400 232838 210452
rect 233326 210400 233332 210452
rect 233384 210440 233390 210452
rect 233970 210440 233976 210452
rect 233384 210412 233976 210440
rect 233384 210400 233390 210412
rect 233970 210400 233976 210412
rect 234028 210400 234034 210452
rect 235994 210400 236000 210452
rect 236052 210440 236058 210452
rect 236822 210440 236828 210452
rect 236052 210412 236828 210440
rect 236052 210400 236058 210412
rect 236822 210400 236828 210412
rect 236880 210400 236886 210452
rect 242986 210400 242992 210452
rect 243044 210440 243050 210452
rect 243814 210440 243820 210452
rect 243044 210412 243820 210440
rect 243044 210400 243050 210412
rect 243814 210400 243820 210412
rect 243872 210400 243878 210452
rect 270126 210400 270132 210452
rect 270184 210440 270190 210452
rect 270310 210440 270316 210452
rect 270184 210412 270316 210440
rect 270184 210400 270190 210412
rect 270310 210400 270316 210412
rect 270368 210400 270374 210452
rect 346946 210400 346952 210452
rect 347004 210440 347010 210452
rect 347682 210440 347688 210452
rect 347004 210412 347688 210440
rect 347004 210400 347010 210412
rect 347682 210400 347688 210412
rect 347740 210400 347746 210452
rect 234614 210332 234620 210384
rect 234672 210372 234678 210384
rect 234890 210372 234896 210384
rect 234672 210344 234896 210372
rect 234672 210332 234678 210344
rect 234890 210332 234896 210344
rect 234948 210332 234954 210384
rect 207106 209788 207112 209840
rect 207164 209828 207170 209840
rect 207382 209828 207388 209840
rect 207164 209800 207388 209828
rect 207164 209788 207170 209800
rect 207382 209788 207388 209800
rect 207440 209788 207446 209840
rect 225138 209720 225144 209772
rect 225196 209760 225202 209772
rect 225414 209760 225420 209772
rect 225196 209732 225420 209760
rect 225196 209720 225202 209732
rect 225414 209720 225420 209732
rect 225472 209720 225478 209772
rect 275830 209720 275836 209772
rect 275888 209760 275894 209772
rect 276106 209760 276112 209772
rect 275888 209732 276112 209760
rect 275888 209720 275894 209732
rect 276106 209720 276112 209732
rect 276164 209720 276170 209772
rect 329374 209760 329380 209772
rect 329335 209732 329380 209760
rect 329374 209720 329380 209732
rect 329432 209720 329438 209772
rect 223574 208496 223580 208548
rect 223632 208536 223638 208548
rect 224126 208536 224132 208548
rect 223632 208508 224132 208536
rect 223632 208496 223638 208508
rect 224126 208496 224132 208508
rect 224184 208496 224190 208548
rect 183830 208360 183836 208412
rect 183888 208400 183894 208412
rect 184566 208400 184572 208412
rect 183888 208372 184572 208400
rect 183888 208360 183894 208372
rect 184566 208360 184572 208372
rect 184624 208360 184630 208412
rect 198826 208292 198832 208344
rect 198884 208332 198890 208344
rect 199654 208332 199660 208344
rect 198884 208304 199660 208332
rect 198884 208292 198890 208304
rect 199654 208292 199660 208304
rect 199712 208292 199718 208344
rect 258258 207720 258264 207732
rect 258219 207692 258264 207720
rect 258258 207680 258264 207692
rect 258316 207680 258322 207732
rect 229186 207000 229192 207052
rect 229244 207040 229250 207052
rect 229830 207040 229836 207052
rect 229244 207012 229836 207040
rect 229244 207000 229250 207012
rect 229830 207000 229836 207012
rect 229888 207000 229894 207052
rect 222194 206456 222200 206508
rect 222252 206496 222258 206508
rect 222930 206496 222936 206508
rect 222252 206468 222936 206496
rect 222252 206456 222258 206468
rect 222930 206456 222936 206468
rect 222988 206456 222994 206508
rect 230658 205844 230664 205896
rect 230716 205884 230722 205896
rect 230842 205884 230848 205896
rect 230716 205856 230848 205884
rect 230716 205844 230722 205856
rect 230842 205844 230848 205856
rect 230900 205844 230906 205896
rect 197446 205708 197452 205760
rect 197504 205748 197510 205760
rect 197630 205748 197636 205760
rect 197504 205720 197636 205748
rect 197504 205708 197510 205720
rect 197630 205708 197636 205720
rect 197688 205708 197694 205760
rect 234798 205708 234804 205760
rect 234856 205708 234862 205760
rect 182266 205640 182272 205692
rect 182324 205680 182330 205692
rect 182542 205680 182548 205692
rect 182324 205652 182548 205680
rect 182324 205640 182330 205652
rect 182542 205640 182548 205652
rect 182600 205640 182606 205692
rect 196066 205640 196072 205692
rect 196124 205680 196130 205692
rect 196342 205680 196348 205692
rect 196124 205652 196348 205680
rect 196124 205640 196130 205652
rect 196342 205640 196348 205652
rect 196400 205640 196406 205692
rect 219802 205680 219808 205692
rect 219763 205652 219808 205680
rect 219802 205640 219808 205652
rect 219860 205640 219866 205692
rect 234816 205624 234844 205708
rect 286594 205640 286600 205692
rect 286652 205640 286658 205692
rect 315850 205680 315856 205692
rect 315811 205652 315856 205680
rect 315850 205640 315856 205652
rect 315908 205640 315914 205692
rect 171410 205572 171416 205624
rect 171468 205612 171474 205624
rect 171594 205612 171600 205624
rect 171468 205584 171600 205612
rect 171468 205572 171474 205584
rect 171594 205572 171600 205584
rect 171652 205572 171658 205624
rect 234798 205572 234804 205624
rect 234856 205572 234862 205624
rect 236270 205572 236276 205624
rect 236328 205612 236334 205624
rect 236454 205612 236460 205624
rect 236328 205584 236460 205612
rect 236328 205572 236334 205584
rect 236454 205572 236460 205584
rect 236512 205572 236518 205624
rect 262582 205612 262588 205624
rect 262543 205584 262588 205612
rect 262582 205572 262588 205584
rect 262640 205572 262646 205624
rect 282638 205504 282644 205556
rect 282696 205544 282702 205556
rect 282822 205544 282828 205556
rect 282696 205516 282828 205544
rect 282696 205504 282702 205516
rect 282822 205504 282828 205516
rect 282880 205504 282886 205556
rect 286612 205544 286640 205640
rect 328089 205615 328147 205621
rect 328089 205581 328101 205615
rect 328135 205612 328147 205615
rect 328178 205612 328184 205624
rect 328135 205584 328184 205612
rect 328135 205581 328147 205584
rect 328089 205575 328147 205581
rect 328178 205572 328184 205584
rect 328236 205572 328242 205624
rect 343266 205612 343272 205624
rect 343227 205584 343272 205612
rect 343266 205572 343272 205584
rect 343324 205572 343330 205624
rect 344554 205612 344560 205624
rect 344515 205584 344560 205612
rect 344554 205572 344560 205584
rect 344612 205572 344618 205624
rect 286686 205544 286692 205556
rect 286612 205516 286692 205544
rect 286686 205504 286692 205516
rect 286744 205504 286750 205556
rect 173342 202852 173348 202904
rect 173400 202892 173406 202904
rect 173434 202892 173440 202904
rect 173400 202864 173440 202892
rect 173400 202852 173406 202864
rect 173434 202852 173440 202864
rect 173492 202852 173498 202904
rect 211893 202895 211951 202901
rect 211893 202861 211905 202895
rect 211939 202892 211951 202895
rect 211982 202892 211988 202904
rect 211939 202864 211988 202892
rect 211939 202861 211951 202864
rect 211893 202855 211951 202861
rect 211982 202852 211988 202864
rect 212040 202852 212046 202904
rect 212166 202852 212172 202904
rect 212224 202892 212230 202904
rect 212442 202892 212448 202904
rect 212224 202864 212448 202892
rect 212224 202852 212230 202864
rect 212442 202852 212448 202864
rect 212500 202852 212506 202904
rect 219802 202892 219808 202904
rect 219763 202864 219808 202892
rect 219802 202852 219808 202864
rect 219860 202852 219866 202904
rect 232130 202852 232136 202904
rect 232188 202892 232194 202904
rect 232314 202892 232320 202904
rect 232188 202864 232320 202892
rect 232188 202852 232194 202864
rect 232314 202852 232320 202864
rect 232372 202852 232378 202904
rect 258261 202895 258319 202901
rect 258261 202861 258273 202895
rect 258307 202892 258319 202895
rect 258350 202892 258356 202904
rect 258307 202864 258356 202892
rect 258307 202861 258319 202864
rect 258261 202855 258319 202861
rect 258350 202852 258356 202864
rect 258408 202852 258414 202904
rect 289170 202852 289176 202904
rect 289228 202892 289234 202904
rect 289446 202892 289452 202904
rect 289228 202864 289452 202892
rect 289228 202852 289234 202864
rect 289446 202852 289452 202864
rect 289504 202852 289510 202904
rect 315850 202892 315856 202904
rect 315811 202864 315856 202892
rect 315850 202852 315856 202864
rect 315908 202852 315914 202904
rect 352834 202852 352840 202904
rect 352892 202892 352898 202904
rect 353018 202892 353024 202904
rect 352892 202864 353024 202892
rect 352892 202852 352898 202864
rect 353018 202852 353024 202864
rect 353076 202852 353082 202904
rect 217045 201535 217103 201541
rect 217045 201501 217057 201535
rect 217091 201532 217103 201535
rect 217134 201532 217140 201544
rect 217091 201504 217140 201532
rect 217091 201501 217103 201504
rect 217045 201495 217103 201501
rect 217134 201492 217140 201504
rect 217192 201492 217198 201544
rect 184106 201424 184112 201476
rect 184164 201464 184170 201476
rect 184290 201464 184296 201476
rect 184164 201436 184296 201464
rect 184164 201424 184170 201436
rect 184290 201424 184296 201436
rect 184348 201424 184354 201476
rect 192113 201467 192171 201473
rect 192113 201433 192125 201467
rect 192159 201464 192171 201467
rect 192386 201464 192392 201476
rect 192159 201436 192392 201464
rect 192159 201433 192171 201436
rect 192113 201427 192171 201433
rect 192386 201424 192392 201436
rect 192444 201424 192450 201476
rect 282822 201464 282828 201476
rect 282783 201436 282828 201464
rect 282822 201424 282828 201436
rect 282880 201424 282886 201476
rect 329377 201467 329435 201473
rect 329377 201433 329389 201467
rect 329423 201464 329435 201467
rect 329466 201464 329472 201476
rect 329423 201436 329472 201464
rect 329423 201433 329435 201436
rect 329377 201427 329435 201433
rect 329466 201424 329472 201436
rect 329524 201424 329530 201476
rect 362497 201467 362555 201473
rect 362497 201433 362509 201467
rect 362543 201464 362555 201467
rect 362586 201464 362592 201476
rect 362543 201436 362592 201464
rect 362543 201433 362555 201436
rect 362497 201427 362555 201433
rect 362586 201424 362592 201436
rect 362644 201424 362650 201476
rect 229462 200064 229468 200116
rect 229520 200104 229526 200116
rect 229554 200104 229560 200116
rect 229520 200076 229560 200104
rect 229520 200064 229526 200076
rect 229554 200064 229560 200076
rect 229612 200064 229618 200116
rect 230842 200064 230848 200116
rect 230900 200104 230906 200116
rect 231394 200104 231400 200116
rect 230900 200076 231400 200104
rect 230900 200064 230906 200076
rect 231394 200064 231400 200076
rect 231452 200064 231458 200116
rect 277210 200104 277216 200116
rect 277171 200076 277216 200104
rect 277210 200064 277216 200076
rect 277268 200064 277274 200116
rect 232130 198132 232136 198144
rect 232056 198104 232136 198132
rect 232056 198076 232084 198104
rect 232130 198092 232136 198104
rect 232188 198092 232194 198144
rect 232038 198024 232044 198076
rect 232096 198024 232102 198076
rect 234982 198024 234988 198076
rect 235040 198064 235046 198076
rect 235626 198064 235632 198076
rect 235040 198036 235632 198064
rect 235040 198024 235046 198036
rect 235626 198024 235632 198036
rect 235684 198024 235690 198076
rect 234798 197956 234804 198008
rect 234856 197996 234862 198008
rect 235166 197996 235172 198008
rect 234856 197968 235172 197996
rect 234856 197956 234862 197968
rect 235166 197956 235172 197968
rect 235224 197956 235230 198008
rect 262398 196596 262404 196648
rect 262456 196636 262462 196648
rect 262674 196636 262680 196648
rect 262456 196608 262680 196636
rect 262456 196596 262462 196608
rect 262674 196596 262680 196608
rect 262732 196596 262738 196648
rect 315761 196095 315819 196101
rect 315761 196061 315773 196095
rect 315807 196092 315819 196095
rect 315850 196092 315856 196104
rect 315807 196064 315856 196092
rect 315807 196061 315819 196064
rect 315761 196055 315819 196061
rect 315850 196052 315856 196064
rect 315908 196052 315914 196104
rect 171502 196024 171508 196036
rect 171463 195996 171508 196024
rect 171502 195984 171508 195996
rect 171560 195984 171566 196036
rect 219802 196024 219808 196036
rect 219728 195996 219808 196024
rect 219728 195968 219756 195996
rect 219802 195984 219808 195996
rect 219860 195984 219866 196036
rect 219710 195916 219716 195968
rect 219768 195916 219774 195968
rect 275830 195236 275836 195288
rect 275888 195276 275894 195288
rect 276106 195276 276112 195288
rect 275888 195248 276112 195276
rect 275888 195236 275894 195248
rect 276106 195236 276112 195248
rect 276164 195236 276170 195288
rect 180058 195168 180064 195220
rect 180116 195208 180122 195220
rect 180150 195208 180156 195220
rect 180116 195180 180156 195208
rect 180116 195168 180122 195180
rect 180150 195168 180156 195180
rect 180208 195168 180214 195220
rect 3142 194488 3148 194540
rect 3200 194528 3206 194540
rect 19978 194528 19984 194540
rect 3200 194500 19984 194528
rect 3200 194488 3206 194500
rect 19978 194488 19984 194500
rect 20036 194488 20042 194540
rect 171502 193236 171508 193248
rect 171463 193208 171508 193236
rect 171502 193196 171508 193208
rect 171560 193196 171566 193248
rect 173158 193196 173164 193248
rect 173216 193236 173222 193248
rect 173526 193236 173532 193248
rect 173216 193208 173532 193236
rect 173216 193196 173222 193208
rect 173526 193196 173532 193208
rect 173584 193196 173590 193248
rect 203242 193196 203248 193248
rect 203300 193236 203306 193248
rect 203334 193236 203340 193248
rect 203300 193208 203340 193236
rect 203300 193196 203306 193208
rect 203334 193196 203340 193208
rect 203392 193196 203398 193248
rect 216674 193196 216680 193248
rect 216732 193236 216738 193248
rect 216950 193236 216956 193248
rect 216732 193208 216956 193236
rect 216732 193196 216738 193208
rect 216950 193196 216956 193208
rect 217008 193196 217014 193248
rect 286502 193196 286508 193248
rect 286560 193236 286566 193248
rect 286686 193236 286692 193248
rect 286560 193208 286692 193236
rect 286560 193196 286566 193208
rect 286686 193196 286692 193208
rect 286744 193196 286750 193248
rect 289262 193196 289268 193248
rect 289320 193236 289326 193248
rect 289446 193236 289452 193248
rect 289320 193208 289452 193236
rect 289320 193196 289326 193208
rect 289446 193196 289452 193208
rect 289504 193196 289510 193248
rect 192110 193168 192116 193180
rect 192071 193140 192116 193168
rect 192110 193128 192116 193140
rect 192168 193128 192174 193180
rect 217134 193128 217140 193180
rect 217192 193168 217198 193180
rect 217226 193168 217232 193180
rect 217192 193140 217232 193168
rect 217192 193128 217198 193140
rect 217226 193128 217232 193140
rect 217284 193128 217290 193180
rect 282822 193168 282828 193180
rect 282783 193140 282828 193168
rect 282822 193128 282828 193140
rect 282880 193128 282886 193180
rect 328181 193103 328239 193109
rect 328181 193069 328193 193103
rect 328227 193100 328239 193103
rect 328270 193100 328276 193112
rect 328227 193072 328276 193100
rect 328227 193069 328239 193072
rect 328181 193063 328239 193069
rect 328270 193060 328276 193072
rect 328328 193060 328334 193112
rect 315758 191876 315764 191888
rect 315719 191848 315764 191876
rect 315758 191836 315764 191848
rect 315816 191836 315822 191888
rect 362494 191876 362500 191888
rect 362455 191848 362500 191876
rect 362494 191836 362500 191848
rect 362552 191836 362558 191888
rect 262490 191808 262496 191820
rect 262451 191780 262496 191808
rect 262490 191768 262496 191780
rect 262548 191768 262554 191820
rect 283834 191768 283840 191820
rect 283892 191808 283898 191820
rect 284018 191808 284024 191820
rect 283892 191780 284024 191808
rect 283892 191768 283898 191780
rect 284018 191768 284024 191780
rect 284076 191768 284082 191820
rect 329558 191808 329564 191820
rect 329519 191780 329564 191808
rect 329558 191768 329564 191780
rect 329616 191768 329622 191820
rect 342990 191768 342996 191820
rect 343048 191808 343054 191820
rect 343174 191808 343180 191820
rect 343048 191780 343180 191808
rect 343048 191768 343054 191780
rect 343174 191768 343180 191780
rect 343232 191768 343238 191820
rect 354214 191808 354220 191820
rect 354175 191780 354220 191808
rect 354214 191768 354220 191780
rect 354272 191768 354278 191820
rect 355410 191768 355416 191820
rect 355468 191808 355474 191820
rect 355502 191808 355508 191820
rect 355468 191780 355508 191808
rect 355468 191768 355474 191780
rect 355502 191768 355508 191780
rect 355560 191768 355566 191820
rect 315669 191743 315727 191749
rect 315669 191709 315681 191743
rect 315715 191740 315727 191743
rect 315758 191740 315764 191752
rect 315715 191712 315764 191740
rect 315715 191709 315727 191712
rect 315669 191703 315727 191709
rect 315758 191700 315764 191712
rect 315816 191700 315822 191752
rect 230566 191088 230572 191140
rect 230624 191128 230630 191140
rect 230750 191128 230756 191140
rect 230624 191100 230756 191128
rect 230624 191088 230630 191100
rect 230750 191088 230756 191100
rect 230808 191088 230814 191140
rect 225230 190408 225236 190460
rect 225288 190448 225294 190460
rect 225414 190448 225420 190460
rect 225288 190420 225420 190448
rect 225288 190408 225294 190420
rect 225414 190408 225420 190420
rect 225472 190408 225478 190460
rect 270126 189864 270132 189916
rect 270184 189904 270190 189916
rect 270310 189904 270316 189916
rect 270184 189876 270316 189904
rect 270184 189864 270190 189876
rect 270310 189864 270316 189876
rect 270368 189864 270374 189916
rect 179969 189023 180027 189029
rect 179969 188989 179981 189023
rect 180015 189020 180027 189023
rect 180058 189020 180064 189032
rect 180015 188992 180064 189020
rect 180015 188989 180027 188992
rect 179969 188983 180027 188989
rect 180058 188980 180064 188992
rect 180116 188980 180122 189032
rect 178862 187796 178868 187808
rect 178236 187768 178868 187796
rect 178236 187740 178264 187768
rect 178862 187756 178868 187768
rect 178920 187756 178926 187808
rect 178218 187688 178224 187740
rect 178276 187688 178282 187740
rect 178218 186436 178224 186448
rect 178144 186408 178224 186436
rect 178144 186312 178172 186408
rect 178218 186396 178224 186408
rect 178276 186396 178282 186448
rect 231026 186436 231032 186448
rect 230952 186408 231032 186436
rect 181162 186368 181168 186380
rect 181088 186340 181168 186368
rect 181088 186312 181116 186340
rect 181162 186328 181168 186340
rect 181220 186328 181226 186380
rect 182174 186328 182180 186380
rect 182232 186368 182238 186380
rect 182232 186340 182277 186368
rect 182232 186328 182238 186340
rect 189442 186328 189448 186380
rect 189500 186328 189506 186380
rect 223942 186328 223948 186380
rect 224000 186328 224006 186380
rect 178126 186260 178132 186312
rect 178184 186260 178190 186312
rect 181070 186260 181076 186312
rect 181128 186260 181134 186312
rect 189460 186232 189488 186328
rect 189534 186232 189540 186244
rect 189460 186204 189540 186232
rect 189534 186192 189540 186204
rect 189592 186192 189598 186244
rect 223960 186232 223988 186328
rect 230952 186312 230980 186408
rect 231026 186396 231032 186408
rect 231084 186396 231090 186448
rect 230934 186260 230940 186312
rect 230992 186260 230998 186312
rect 262490 186300 262496 186312
rect 262451 186272 262496 186300
rect 262490 186260 262496 186272
rect 262548 186260 262554 186312
rect 328178 186300 328184 186312
rect 328139 186272 328184 186300
rect 328178 186260 328184 186272
rect 328236 186260 328242 186312
rect 224034 186232 224040 186244
rect 223960 186204 224040 186232
rect 224034 186192 224040 186204
rect 224092 186192 224098 186244
rect 184014 183608 184020 183660
rect 184072 183648 184078 183660
rect 184106 183648 184112 183660
rect 184072 183620 184112 183648
rect 184072 183608 184078 183620
rect 184106 183608 184112 183620
rect 184164 183608 184170 183660
rect 275830 183608 275836 183660
rect 275888 183608 275894 183660
rect 286686 183648 286692 183660
rect 286612 183620 286692 183648
rect 192110 183540 192116 183592
rect 192168 183580 192174 183592
rect 192202 183580 192208 183592
rect 192168 183552 192208 183580
rect 192168 183540 192174 183552
rect 192202 183540 192208 183552
rect 192260 183540 192266 183592
rect 232130 183540 232136 183592
rect 232188 183580 232194 183592
rect 232222 183580 232228 183592
rect 232188 183552 232228 183580
rect 232188 183540 232194 183552
rect 232222 183540 232228 183552
rect 232280 183540 232286 183592
rect 234982 183540 234988 183592
rect 235040 183580 235046 183592
rect 235074 183580 235080 183592
rect 235040 183552 235080 183580
rect 235040 183540 235046 183552
rect 235074 183540 235080 183552
rect 235132 183540 235138 183592
rect 275848 183524 275876 183608
rect 286612 183592 286640 183620
rect 286686 183608 286692 183620
rect 286744 183608 286750 183660
rect 344370 183608 344376 183660
rect 344428 183648 344434 183660
rect 344554 183648 344560 183660
rect 344428 183620 344560 183648
rect 344428 183608 344434 183620
rect 344554 183608 344560 183620
rect 344612 183608 344618 183660
rect 277210 183580 277216 183592
rect 277171 183552 277216 183580
rect 277210 183540 277216 183552
rect 277268 183540 277274 183592
rect 282730 183540 282736 183592
rect 282788 183580 282794 183592
rect 282914 183580 282920 183592
rect 282788 183552 282920 183580
rect 282788 183540 282794 183552
rect 282914 183540 282920 183552
rect 282972 183540 282978 183592
rect 286594 183540 286600 183592
rect 286652 183540 286658 183592
rect 289262 183540 289268 183592
rect 289320 183580 289326 183592
rect 289446 183580 289452 183592
rect 289320 183552 289452 183580
rect 289320 183540 289326 183552
rect 289446 183540 289452 183552
rect 289504 183540 289510 183592
rect 291654 183540 291660 183592
rect 291712 183580 291718 183592
rect 291930 183580 291936 183592
rect 291712 183552 291936 183580
rect 291712 183540 291718 183552
rect 291930 183540 291936 183552
rect 291988 183540 291994 183592
rect 275830 183472 275836 183524
rect 275888 183472 275894 183524
rect 354214 183512 354220 183524
rect 354175 183484 354220 183512
rect 354214 183472 354220 183484
rect 354272 183472 354278 183524
rect 182174 182180 182180 182232
rect 182232 182220 182238 182232
rect 315666 182220 315672 182232
rect 182232 182192 182277 182220
rect 315627 182192 315672 182220
rect 182232 182180 182238 182192
rect 315666 182180 315672 182192
rect 315724 182180 315730 182232
rect 184106 182112 184112 182164
rect 184164 182152 184170 182164
rect 184198 182152 184204 182164
rect 184164 182124 184204 182152
rect 184164 182112 184170 182124
rect 184198 182112 184204 182124
rect 184256 182112 184262 182164
rect 192202 182152 192208 182164
rect 192163 182124 192208 182152
rect 192202 182112 192208 182124
rect 192260 182112 192266 182164
rect 224034 182152 224040 182164
rect 223995 182124 224040 182152
rect 224034 182112 224040 182124
rect 224092 182112 224098 182164
rect 228266 182112 228272 182164
rect 228324 182152 228330 182164
rect 228358 182152 228364 182164
rect 228324 182124 228364 182152
rect 228324 182112 228330 182124
rect 228358 182112 228364 182124
rect 228416 182112 228422 182164
rect 229278 182112 229284 182164
rect 229336 182152 229342 182164
rect 229462 182152 229468 182164
rect 229336 182124 229468 182152
rect 229336 182112 229342 182124
rect 229462 182112 229468 182124
rect 229520 182112 229526 182164
rect 230934 182112 230940 182164
rect 230992 182152 230998 182164
rect 231026 182152 231032 182164
rect 230992 182124 231032 182152
rect 230992 182112 230998 182124
rect 231026 182112 231032 182124
rect 231084 182112 231090 182164
rect 236270 182112 236276 182164
rect 236328 182152 236334 182164
rect 236454 182152 236460 182164
rect 236328 182124 236460 182152
rect 236328 182112 236334 182124
rect 236454 182112 236460 182124
rect 236512 182112 236518 182164
rect 261110 182112 261116 182164
rect 261168 182152 261174 182164
rect 261294 182152 261300 182164
rect 261168 182124 261300 182152
rect 261168 182112 261174 182124
rect 261294 182112 261300 182124
rect 261352 182112 261358 182164
rect 277121 182155 277179 182161
rect 277121 182121 277133 182155
rect 277167 182152 277179 182155
rect 277210 182152 277216 182164
rect 277167 182124 277216 182152
rect 277167 182121 277179 182124
rect 277121 182115 277179 182121
rect 277210 182112 277216 182124
rect 277268 182112 277274 182164
rect 282822 182112 282828 182164
rect 282880 182152 282886 182164
rect 282914 182152 282920 182164
rect 282880 182124 282920 182152
rect 282880 182112 282886 182124
rect 282914 182112 282920 182124
rect 282972 182112 282978 182164
rect 285214 182152 285220 182164
rect 285175 182124 285220 182152
rect 285214 182112 285220 182124
rect 285272 182112 285278 182164
rect 354306 182152 354312 182164
rect 354267 182124 354312 182152
rect 354306 182112 354312 182124
rect 354364 182112 354370 182164
rect 355594 182152 355600 182164
rect 355555 182124 355600 182152
rect 355594 182112 355600 182124
rect 355652 182112 355658 182164
rect 360930 182112 360936 182164
rect 360988 182152 360994 182164
rect 361206 182152 361212 182164
rect 360988 182124 361212 182152
rect 360988 182112 360994 182124
rect 361206 182112 361212 182124
rect 361264 182112 361270 182164
rect 362405 182155 362463 182161
rect 362405 182121 362417 182155
rect 362451 182152 362463 182155
rect 362586 182152 362592 182164
rect 362451 182124 362592 182152
rect 362451 182121 362463 182124
rect 362405 182115 362463 182121
rect 362586 182112 362592 182124
rect 362644 182112 362650 182164
rect 262582 182084 262588 182096
rect 262543 182056 262588 182084
rect 262582 182044 262588 182056
rect 262640 182044 262646 182096
rect 182174 181976 182180 182028
rect 182232 182016 182238 182028
rect 182232 181988 182277 182016
rect 182232 181976 182238 181988
rect 329374 181568 329380 181620
rect 329432 181608 329438 181620
rect 329561 181611 329619 181617
rect 329561 181608 329573 181611
rect 329432 181580 329573 181608
rect 329432 181568 329438 181580
rect 329561 181577 329573 181580
rect 329607 181577 329619 181611
rect 329561 181571 329619 181577
rect 230566 181432 230572 181484
rect 230624 181472 230630 181484
rect 230750 181472 230756 181484
rect 230624 181444 230756 181472
rect 230624 181432 230630 181444
rect 230750 181432 230756 181444
rect 230808 181432 230814 181484
rect 270126 181432 270132 181484
rect 270184 181472 270190 181484
rect 270310 181472 270316 181484
rect 270184 181444 270316 181472
rect 270184 181432 270190 181444
rect 270310 181432 270316 181444
rect 270368 181432 270374 181484
rect 217318 180792 217324 180804
rect 217279 180764 217324 180792
rect 217318 180752 217324 180764
rect 217376 180752 217382 180804
rect 275830 180792 275836 180804
rect 275791 180764 275836 180792
rect 275830 180752 275836 180764
rect 275888 180752 275894 180804
rect 179966 179432 179972 179444
rect 179927 179404 179972 179432
rect 179966 179392 179972 179404
rect 180024 179392 180030 179444
rect 176933 179367 176991 179373
rect 176933 179333 176945 179367
rect 176979 179364 176991 179367
rect 177114 179364 177120 179376
rect 176979 179336 177120 179364
rect 176979 179333 176991 179336
rect 176933 179327 176991 179333
rect 177114 179324 177120 179336
rect 177172 179324 177178 179376
rect 181070 179364 181076 179376
rect 181031 179336 181076 179364
rect 181070 179324 181076 179336
rect 181128 179324 181134 179376
rect 291930 176740 291936 176792
rect 291988 176740 291994 176792
rect 211706 176672 211712 176724
rect 211764 176712 211770 176724
rect 211982 176712 211988 176724
rect 211764 176684 211988 176712
rect 211764 176672 211770 176684
rect 211982 176672 211988 176684
rect 212040 176672 212046 176724
rect 291948 176588 291976 176740
rect 344554 176604 344560 176656
rect 344612 176604 344618 176656
rect 355594 176644 355600 176656
rect 355555 176616 355600 176644
rect 355594 176604 355600 176616
rect 355652 176604 355658 176656
rect 182177 176579 182235 176585
rect 182177 176545 182189 176579
rect 182223 176576 182235 176579
rect 182266 176576 182272 176588
rect 182223 176548 182272 176576
rect 182223 176545 182235 176548
rect 182177 176539 182235 176545
rect 182266 176536 182272 176548
rect 182324 176536 182330 176588
rect 291930 176536 291936 176588
rect 291988 176536 291994 176588
rect 344462 176536 344468 176588
rect 344520 176576 344526 176588
rect 344572 176576 344600 176604
rect 344520 176548 344600 176576
rect 354309 176579 354367 176585
rect 344520 176536 344526 176548
rect 354309 176545 354321 176579
rect 354355 176576 354367 176579
rect 354398 176576 354404 176588
rect 354355 176548 354404 176576
rect 354355 176545 354367 176548
rect 354309 176539 354367 176545
rect 354398 176536 354404 176548
rect 354456 176536 354462 176588
rect 192202 176100 192208 176112
rect 192163 176072 192208 176100
rect 192202 176060 192208 176072
rect 192260 176060 192266 176112
rect 232130 173952 232136 174004
rect 232188 173992 232194 174004
rect 232222 173992 232228 174004
rect 232188 173964 232228 173992
rect 232188 173952 232194 173964
rect 232222 173952 232228 173964
rect 232280 173952 232286 174004
rect 173066 173884 173072 173936
rect 173124 173924 173130 173936
rect 173158 173924 173164 173936
rect 173124 173896 173164 173924
rect 173124 173884 173130 173896
rect 173158 173884 173164 173896
rect 173216 173884 173222 173936
rect 216674 173884 216680 173936
rect 216732 173924 216738 173936
rect 216950 173924 216956 173936
rect 216732 173896 216956 173924
rect 216732 173884 216738 173896
rect 216950 173884 216956 173896
rect 217008 173884 217014 173936
rect 219802 173884 219808 173936
rect 219860 173924 219866 173936
rect 219986 173924 219992 173936
rect 219860 173896 219992 173924
rect 219860 173884 219866 173896
rect 219986 173884 219992 173896
rect 220044 173884 220050 173936
rect 286502 173884 286508 173936
rect 286560 173884 286566 173936
rect 289262 173884 289268 173936
rect 289320 173924 289326 173936
rect 289446 173924 289452 173936
rect 289320 173896 289452 173924
rect 289320 173884 289326 173896
rect 289446 173884 289452 173896
rect 289504 173884 289510 173936
rect 329374 173884 329380 173936
rect 329432 173924 329438 173936
rect 329558 173924 329564 173936
rect 329432 173896 329564 173924
rect 329432 173884 329438 173896
rect 329558 173884 329564 173896
rect 329616 173884 329622 173936
rect 286520 173788 286548 173884
rect 286594 173788 286600 173800
rect 286520 173760 286600 173788
rect 286594 173748 286600 173760
rect 286652 173748 286658 173800
rect 176933 173179 176991 173185
rect 176933 173145 176945 173179
rect 176979 173176 176991 173179
rect 177114 173176 177120 173188
rect 176979 173148 177120 173176
rect 176979 173145 176991 173148
rect 176933 173139 176991 173145
rect 177114 173136 177120 173148
rect 177172 173136 177178 173188
rect 189442 172524 189448 172576
rect 189500 172564 189506 172576
rect 189534 172564 189540 172576
rect 189500 172536 189540 172564
rect 189500 172524 189506 172536
rect 189534 172524 189540 172536
rect 189592 172524 189598 172576
rect 194962 172524 194968 172576
rect 195020 172564 195026 172576
rect 195054 172564 195060 172576
rect 195020 172536 195060 172564
rect 195020 172524 195026 172536
rect 195054 172524 195060 172536
rect 195112 172524 195118 172576
rect 224034 172564 224040 172576
rect 223995 172536 224040 172564
rect 224034 172524 224040 172536
rect 224092 172524 224098 172576
rect 262582 172564 262588 172576
rect 262543 172536 262588 172564
rect 262582 172524 262588 172536
rect 262640 172524 262646 172576
rect 277118 172564 277124 172576
rect 277079 172536 277124 172564
rect 277118 172524 277124 172536
rect 277176 172524 277182 172576
rect 225414 172496 225420 172508
rect 225375 172468 225420 172496
rect 225414 172456 225420 172468
rect 225472 172456 225478 172508
rect 229370 172496 229376 172508
rect 229331 172468 229376 172496
rect 229370 172456 229376 172468
rect 229428 172456 229434 172508
rect 283834 172456 283840 172508
rect 283892 172496 283898 172508
rect 284018 172496 284024 172508
rect 283892 172468 284024 172496
rect 283892 172456 283898 172468
rect 284018 172456 284024 172468
rect 284076 172456 284082 172508
rect 345474 172456 345480 172508
rect 345532 172496 345538 172508
rect 345658 172496 345664 172508
rect 345532 172468 345664 172496
rect 345532 172456 345538 172468
rect 345658 172456 345664 172468
rect 345716 172456 345722 172508
rect 361114 172456 361120 172508
rect 361172 172496 361178 172508
rect 361390 172496 361396 172508
rect 361172 172468 361396 172496
rect 361172 172456 361178 172468
rect 361390 172456 361396 172468
rect 361448 172456 361454 172508
rect 362310 171164 362316 171216
rect 362368 171204 362374 171216
rect 362405 171207 362463 171213
rect 362405 171204 362417 171207
rect 362368 171176 362417 171204
rect 362368 171164 362374 171176
rect 362405 171173 362417 171176
rect 362451 171173 362463 171207
rect 362405 171167 362463 171173
rect 203150 171096 203156 171148
rect 203208 171136 203214 171148
rect 203242 171136 203248 171148
rect 203208 171108 203248 171136
rect 203208 171096 203214 171108
rect 203242 171096 203248 171108
rect 203300 171096 203306 171148
rect 217321 171139 217379 171145
rect 217321 171105 217333 171139
rect 217367 171136 217379 171139
rect 217410 171136 217416 171148
rect 217367 171108 217416 171136
rect 217367 171105 217379 171108
rect 217321 171099 217379 171105
rect 217410 171096 217416 171108
rect 217468 171096 217474 171148
rect 275833 171139 275891 171145
rect 275833 171105 275845 171139
rect 275879 171136 275891 171139
rect 275922 171136 275928 171148
rect 275879 171108 275928 171136
rect 275879 171105 275891 171108
rect 275833 171099 275891 171105
rect 275922 171096 275928 171108
rect 275980 171096 275986 171148
rect 182177 171071 182235 171077
rect 182177 171037 182189 171071
rect 182223 171068 182235 171071
rect 182266 171068 182272 171080
rect 182223 171040 182272 171068
rect 182223 171037 182235 171040
rect 182177 171031 182235 171037
rect 182266 171028 182272 171040
rect 182324 171028 182330 171080
rect 211706 171028 211712 171080
rect 211764 171068 211770 171080
rect 211893 171071 211951 171077
rect 211893 171068 211905 171071
rect 211764 171040 211905 171068
rect 211764 171028 211770 171040
rect 211893 171037 211905 171040
rect 211939 171037 211951 171071
rect 236362 171068 236368 171080
rect 236323 171040 236368 171068
rect 211893 171031 211951 171037
rect 236362 171028 236368 171040
rect 236420 171028 236426 171080
rect 362402 171068 362408 171080
rect 362363 171040 362408 171068
rect 362402 171028 362408 171040
rect 362460 171028 362466 171080
rect 376018 171028 376024 171080
rect 376076 171068 376082 171080
rect 580166 171068 580172 171080
rect 376076 171040 580172 171068
rect 376076 171028 376082 171040
rect 580166 171028 580172 171040
rect 580224 171028 580230 171080
rect 270126 170552 270132 170604
rect 270184 170592 270190 170604
rect 270310 170592 270316 170604
rect 270184 170564 270316 170592
rect 270184 170552 270190 170564
rect 270310 170552 270316 170564
rect 270368 170552 270374 170604
rect 181073 169779 181131 169785
rect 181073 169745 181085 169779
rect 181119 169776 181131 169779
rect 181346 169776 181352 169788
rect 181119 169748 181352 169776
rect 181119 169745 181131 169748
rect 181073 169739 181131 169745
rect 181346 169736 181352 169748
rect 181404 169736 181410 169788
rect 343266 169668 343272 169720
rect 343324 169708 343330 169720
rect 343358 169708 343364 169720
rect 343324 169680 343364 169708
rect 343324 169668 343330 169680
rect 343358 169668 343364 169680
rect 343416 169668 343422 169720
rect 318429 169167 318487 169173
rect 318429 169133 318441 169167
rect 318475 169164 318487 169167
rect 318518 169164 318524 169176
rect 318475 169136 318524 169164
rect 318475 169133 318487 169136
rect 318429 169127 318487 169133
rect 318518 169124 318524 169136
rect 318576 169124 318582 169176
rect 327994 169056 328000 169108
rect 328052 169096 328058 169108
rect 328178 169096 328184 169108
rect 328052 169068 328184 169096
rect 328052 169056 328058 169068
rect 328178 169056 328184 169068
rect 328236 169056 328242 169108
rect 329282 169056 329288 169108
rect 329340 169096 329346 169108
rect 329466 169096 329472 169108
rect 329340 169068 329472 169096
rect 329340 169056 329346 169068
rect 329466 169056 329472 169068
rect 329524 169056 329530 169108
rect 177114 168348 177120 168360
rect 177075 168320 177120 168348
rect 177114 168308 177120 168320
rect 177172 168308 177178 168360
rect 344557 167535 344615 167541
rect 344557 167501 344569 167535
rect 344603 167532 344615 167535
rect 344646 167532 344652 167544
rect 344603 167504 344652 167532
rect 344603 167501 344615 167504
rect 344557 167495 344615 167501
rect 344646 167492 344652 167504
rect 344704 167492 344710 167544
rect 232130 167084 232136 167136
rect 232188 167084 232194 167136
rect 273070 167124 273076 167136
rect 272996 167096 273076 167124
rect 232148 167000 232176 167084
rect 258166 167016 258172 167068
rect 258224 167056 258230 167068
rect 258350 167056 258356 167068
rect 258224 167028 258356 167056
rect 258224 167016 258230 167028
rect 258350 167016 258356 167028
rect 258408 167016 258414 167068
rect 232130 166948 232136 167000
rect 232188 166948 232194 167000
rect 272996 166932 273024 167096
rect 273070 167084 273076 167096
rect 273128 167084 273134 167136
rect 317046 167016 317052 167068
rect 317104 167056 317110 167068
rect 355597 167059 355655 167065
rect 317104 167028 317184 167056
rect 317104 167016 317110 167028
rect 317156 167000 317184 167028
rect 355597 167025 355609 167059
rect 355643 167056 355655 167059
rect 355686 167056 355692 167068
rect 355643 167028 355692 167056
rect 355643 167025 355655 167028
rect 355597 167019 355655 167025
rect 355686 167016 355692 167028
rect 355744 167016 355750 167068
rect 317138 166948 317144 167000
rect 317196 166948 317202 167000
rect 272978 166880 272984 166932
rect 273036 166880 273042 166932
rect 285217 166923 285275 166929
rect 285217 166889 285229 166923
rect 285263 166920 285275 166923
rect 285306 166920 285312 166932
rect 285263 166892 285312 166920
rect 285263 166889 285275 166892
rect 285217 166883 285275 166889
rect 285306 166880 285312 166892
rect 285364 166880 285370 166932
rect 2774 165452 2780 165504
rect 2832 165492 2838 165504
rect 5166 165492 5172 165504
rect 2832 165464 5172 165492
rect 2832 165452 2838 165464
rect 5166 165452 5172 165464
rect 5224 165452 5230 165504
rect 217226 164228 217232 164280
rect 217284 164268 217290 164280
rect 217410 164268 217416 164280
rect 217284 164240 217416 164268
rect 217284 164228 217290 164240
rect 217410 164228 217416 164240
rect 217468 164228 217474 164280
rect 235258 164228 235264 164280
rect 235316 164268 235322 164280
rect 235350 164268 235356 164280
rect 235316 164240 235356 164268
rect 235316 164228 235322 164240
rect 235350 164228 235356 164240
rect 235408 164228 235414 164280
rect 315666 164228 315672 164280
rect 315724 164268 315730 164280
rect 315758 164268 315764 164280
rect 315724 164240 315764 164268
rect 315724 164228 315730 164240
rect 315758 164228 315764 164240
rect 315816 164228 315822 164280
rect 318426 164268 318432 164280
rect 318387 164240 318432 164268
rect 318426 164228 318432 164240
rect 318484 164228 318490 164280
rect 354306 164228 354312 164280
rect 354364 164268 354370 164280
rect 354398 164268 354404 164280
rect 354364 164240 354404 164268
rect 354364 164228 354370 164240
rect 354398 164228 354404 164240
rect 354456 164228 354462 164280
rect 355594 164268 355600 164280
rect 355555 164240 355600 164268
rect 355594 164228 355600 164240
rect 355652 164228 355658 164280
rect 171410 164160 171416 164212
rect 171468 164200 171474 164212
rect 171594 164200 171600 164212
rect 171468 164172 171600 164200
rect 171468 164160 171474 164172
rect 171594 164160 171600 164172
rect 171652 164160 171658 164212
rect 173066 164160 173072 164212
rect 173124 164200 173130 164212
rect 173250 164200 173256 164212
rect 173124 164172 173256 164200
rect 173124 164160 173130 164172
rect 173250 164160 173256 164172
rect 173308 164160 173314 164212
rect 184014 164160 184020 164212
rect 184072 164200 184078 164212
rect 184106 164200 184112 164212
rect 184072 164172 184112 164200
rect 184072 164160 184078 164172
rect 184106 164160 184112 164172
rect 184164 164160 184170 164212
rect 189350 164160 189356 164212
rect 189408 164200 189414 164212
rect 189442 164200 189448 164212
rect 189408 164172 189448 164200
rect 189408 164160 189414 164172
rect 189442 164160 189448 164172
rect 189500 164160 189506 164212
rect 212442 164200 212448 164212
rect 212403 164172 212448 164200
rect 212442 164160 212448 164172
rect 212500 164160 212506 164212
rect 229370 164200 229376 164212
rect 229331 164172 229376 164200
rect 229370 164160 229376 164172
rect 229428 164160 229434 164212
rect 235074 164160 235080 164212
rect 235132 164160 235138 164212
rect 258258 164200 258264 164212
rect 258219 164172 258264 164200
rect 258258 164160 258264 164172
rect 258316 164160 258322 164212
rect 262306 164160 262312 164212
rect 262364 164200 262370 164212
rect 262490 164200 262496 164212
rect 262364 164172 262496 164200
rect 262364 164160 262370 164172
rect 262490 164160 262496 164172
rect 262548 164160 262554 164212
rect 286594 164160 286600 164212
rect 286652 164200 286658 164212
rect 286686 164200 286692 164212
rect 286652 164172 286692 164200
rect 286652 164160 286658 164172
rect 286686 164160 286692 164172
rect 286744 164160 286750 164212
rect 289354 164160 289360 164212
rect 289412 164200 289418 164212
rect 289446 164200 289452 164212
rect 289412 164172 289452 164200
rect 289412 164160 289418 164172
rect 289446 164160 289452 164172
rect 289504 164160 289510 164212
rect 235092 164132 235120 164160
rect 235166 164132 235172 164144
rect 235092 164104 235172 164132
rect 235166 164092 235172 164104
rect 235224 164092 235230 164144
rect 344554 162908 344560 162920
rect 344515 162880 344560 162908
rect 344554 162868 344560 162880
rect 344612 162868 344618 162920
rect 229281 162843 229339 162849
rect 229281 162809 229293 162843
rect 229327 162840 229339 162843
rect 229462 162840 229468 162852
rect 229327 162812 229468 162840
rect 229327 162809 229339 162812
rect 229281 162803 229339 162809
rect 229462 162800 229468 162812
rect 229520 162800 229526 162852
rect 261110 162840 261116 162852
rect 261071 162812 261116 162840
rect 261110 162800 261116 162812
rect 261168 162800 261174 162852
rect 275830 162800 275836 162852
rect 275888 162840 275894 162852
rect 275922 162840 275928 162852
rect 275888 162812 275928 162840
rect 275888 162800 275894 162812
rect 275922 162800 275928 162812
rect 275980 162800 275986 162852
rect 282638 162800 282644 162852
rect 282696 162840 282702 162852
rect 282822 162840 282828 162852
rect 282696 162812 282828 162840
rect 282696 162800 282702 162812
rect 282822 162800 282828 162812
rect 282880 162800 282886 162852
rect 286686 162840 286692 162852
rect 286647 162812 286692 162840
rect 286686 162800 286692 162812
rect 286744 162800 286750 162852
rect 289262 162800 289268 162852
rect 289320 162840 289326 162852
rect 289446 162840 289452 162852
rect 289320 162812 289452 162840
rect 289320 162800 289326 162812
rect 289446 162800 289452 162812
rect 289504 162800 289510 162852
rect 317138 162840 317144 162852
rect 317099 162812 317144 162840
rect 317138 162800 317144 162812
rect 317196 162800 317202 162852
rect 318426 162840 318432 162852
rect 318387 162812 318432 162840
rect 318426 162800 318432 162812
rect 318484 162800 318490 162852
rect 341978 162840 341984 162852
rect 341939 162812 341984 162840
rect 341978 162800 341984 162812
rect 342036 162800 342042 162852
rect 354306 162840 354312 162852
rect 354267 162812 354312 162840
rect 354306 162800 354312 162812
rect 354364 162800 354370 162852
rect 355505 162843 355563 162849
rect 355505 162809 355517 162843
rect 355551 162840 355563 162843
rect 355594 162840 355600 162852
rect 355551 162812 355600 162840
rect 355551 162809 355563 162812
rect 355505 162803 355563 162809
rect 355594 162800 355600 162812
rect 355652 162800 355658 162852
rect 225414 162704 225420 162716
rect 225375 162676 225420 162704
rect 225414 162664 225420 162676
rect 225472 162664 225478 162716
rect 270126 162120 270132 162172
rect 270184 162160 270190 162172
rect 270310 162160 270316 162172
rect 270184 162132 270316 162160
rect 270184 162120 270190 162132
rect 270310 162120 270316 162132
rect 270368 162120 270374 162172
rect 182174 161480 182180 161492
rect 182135 161452 182180 161480
rect 182174 161440 182180 161452
rect 182232 161440 182238 161492
rect 362402 161480 362408 161492
rect 362363 161452 362408 161480
rect 362402 161440 362408 161452
rect 362460 161440 362466 161492
rect 181070 161412 181076 161424
rect 181031 161384 181076 161412
rect 181070 161372 181076 161384
rect 181128 161372 181134 161424
rect 203150 161412 203156 161424
rect 203111 161384 203156 161412
rect 203150 161372 203156 161384
rect 203208 161372 203214 161424
rect 217137 161415 217195 161421
rect 217137 161381 217149 161415
rect 217183 161412 217195 161415
rect 217226 161412 217232 161424
rect 217183 161384 217232 161412
rect 217183 161381 217195 161384
rect 217137 161375 217195 161381
rect 217226 161372 217232 161384
rect 217284 161372 217290 161424
rect 345658 161412 345664 161424
rect 345619 161384 345664 161412
rect 345658 161372 345664 161384
rect 345716 161372 345722 161424
rect 182174 161344 182180 161356
rect 182135 161316 182180 161344
rect 182174 161304 182180 161316
rect 182232 161304 182238 161356
rect 236365 160191 236423 160197
rect 236365 160188 236377 160191
rect 236288 160160 236377 160188
rect 236288 160132 236316 160160
rect 236365 160157 236377 160160
rect 236411 160157 236423 160191
rect 236365 160151 236423 160157
rect 236270 160080 236276 160132
rect 236328 160080 236334 160132
rect 225414 160012 225420 160064
rect 225472 160052 225478 160064
rect 225598 160052 225604 160064
rect 225472 160024 225604 160052
rect 225472 160012 225478 160024
rect 225598 160012 225604 160024
rect 225656 160012 225662 160064
rect 361206 160052 361212 160064
rect 361167 160024 361212 160052
rect 361206 160012 361212 160024
rect 361264 160012 361270 160064
rect 177114 158760 177120 158772
rect 177075 158732 177120 158760
rect 177114 158720 177120 158732
rect 177172 158720 177178 158772
rect 178034 158652 178040 158704
rect 178092 158692 178098 158704
rect 178126 158692 178132 158704
rect 178092 158664 178132 158692
rect 178092 158652 178098 158664
rect 178126 158652 178132 158664
rect 178184 158652 178190 158704
rect 225598 158692 225604 158704
rect 225559 158664 225604 158692
rect 225598 158652 225604 158664
rect 225656 158652 225662 158704
rect 228358 158652 228364 158704
rect 228416 158692 228422 158704
rect 228542 158692 228548 158704
rect 228416 158664 228548 158692
rect 228416 158652 228422 158664
rect 228542 158652 228548 158664
rect 228600 158652 228606 158704
rect 343266 158692 343272 158704
rect 343227 158664 343272 158692
rect 343266 158652 343272 158664
rect 343324 158652 343330 158704
rect 272978 157972 272984 158024
rect 273036 158012 273042 158024
rect 273254 158012 273260 158024
rect 273036 157984 273260 158012
rect 273036 157972 273042 157984
rect 273254 157972 273260 157984
rect 273312 157972 273318 158024
rect 328178 157360 328184 157412
rect 328236 157360 328242 157412
rect 329466 157360 329472 157412
rect 329524 157360 329530 157412
rect 228177 157335 228235 157341
rect 228177 157301 228189 157335
rect 228223 157332 228235 157335
rect 228542 157332 228548 157344
rect 228223 157304 228548 157332
rect 228223 157301 228235 157304
rect 228177 157295 228235 157301
rect 228542 157292 228548 157304
rect 228600 157292 228606 157344
rect 258258 157332 258264 157344
rect 258219 157304 258264 157332
rect 258258 157292 258264 157304
rect 258316 157292 258322 157344
rect 291930 157292 291936 157344
rect 291988 157292 291994 157344
rect 317138 157332 317144 157344
rect 317099 157304 317144 157332
rect 317138 157292 317144 157304
rect 317196 157292 317202 157344
rect 318426 157332 318432 157344
rect 318387 157304 318432 157332
rect 318426 157292 318432 157304
rect 318484 157292 318490 157344
rect 232130 157264 232136 157276
rect 232056 157236 232136 157264
rect 232056 157140 232084 157236
rect 232130 157224 232136 157236
rect 232188 157224 232194 157276
rect 291948 157208 291976 157292
rect 328196 157264 328224 157360
rect 328270 157264 328276 157276
rect 328196 157236 328276 157264
rect 328270 157224 328276 157236
rect 328328 157224 328334 157276
rect 329484 157264 329512 157360
rect 354306 157332 354312 157344
rect 354267 157304 354312 157332
rect 354306 157292 354312 157304
rect 354364 157292 354370 157344
rect 329558 157264 329564 157276
rect 329484 157236 329564 157264
rect 329558 157224 329564 157236
rect 329616 157224 329622 157276
rect 291930 157156 291936 157208
rect 291988 157156 291994 157208
rect 232038 157088 232044 157140
rect 232096 157088 232102 157140
rect 192202 156788 192208 156800
rect 192163 156760 192208 156788
rect 192202 156748 192208 156760
rect 192260 156748 192266 156800
rect 182174 156720 182180 156732
rect 182135 156692 182180 156720
rect 182174 156680 182180 156692
rect 182232 156680 182238 156732
rect 362402 156652 362408 156664
rect 362363 156624 362408 156652
rect 362402 156612 362408 156624
rect 362460 156612 362466 156664
rect 273162 154640 273168 154692
rect 273220 154640 273226 154692
rect 211890 154612 211896 154624
rect 211851 154584 211896 154612
rect 211890 154572 211896 154584
rect 211948 154572 211954 154624
rect 212442 154612 212448 154624
rect 212403 154584 212448 154612
rect 212442 154572 212448 154584
rect 212500 154572 212506 154624
rect 273180 154556 273208 154640
rect 234982 154504 234988 154556
rect 235040 154544 235046 154556
rect 235166 154544 235172 154556
rect 235040 154516 235172 154544
rect 235040 154504 235046 154516
rect 235166 154504 235172 154516
rect 235224 154504 235230 154556
rect 273162 154504 273168 154556
rect 273220 154504 273226 154556
rect 291930 154544 291936 154556
rect 291891 154516 291936 154544
rect 291930 154504 291936 154516
rect 291988 154504 291994 154556
rect 315758 153280 315764 153332
rect 315816 153320 315822 153332
rect 315850 153320 315856 153332
rect 315816 153292 315856 153320
rect 315816 153280 315822 153292
rect 315850 153280 315856 153292
rect 315908 153280 315914 153332
rect 192110 153212 192116 153264
rect 192168 153252 192174 153264
rect 192205 153255 192263 153261
rect 192205 153252 192217 153255
rect 192168 153224 192217 153252
rect 192168 153212 192174 153224
rect 192205 153221 192217 153224
rect 192251 153221 192263 153255
rect 229278 153252 229284 153264
rect 229239 153224 229284 153252
rect 192205 153215 192263 153221
rect 229278 153212 229284 153224
rect 229336 153212 229342 153264
rect 261110 153252 261116 153264
rect 261071 153224 261116 153252
rect 261110 153212 261116 153224
rect 261168 153212 261174 153264
rect 283834 153212 283840 153264
rect 283892 153252 283898 153264
rect 283926 153252 283932 153264
rect 283892 153224 283932 153252
rect 283892 153212 283898 153224
rect 283926 153212 283932 153224
rect 283984 153212 283990 153264
rect 286686 153252 286692 153264
rect 286647 153224 286692 153252
rect 286686 153212 286692 153224
rect 286744 153212 286750 153264
rect 341978 153252 341984 153264
rect 341939 153224 341984 153252
rect 341978 153212 341984 153224
rect 342036 153212 342042 153264
rect 355502 153252 355508 153264
rect 355463 153224 355508 153252
rect 355502 153212 355508 153224
rect 355560 153212 355566 153264
rect 191098 153144 191104 153196
rect 191156 153184 191162 153196
rect 191190 153184 191196 153196
rect 191156 153156 191196 153184
rect 191156 153144 191162 153156
rect 191190 153144 191196 153156
rect 191248 153144 191254 153196
rect 230934 153184 230940 153196
rect 230895 153156 230940 153184
rect 230934 153144 230940 153156
rect 230992 153144 230998 153196
rect 231762 153144 231768 153196
rect 231820 153184 231826 153196
rect 232038 153184 232044 153196
rect 231820 153156 232044 153184
rect 231820 153144 231826 153156
rect 232038 153144 232044 153156
rect 232096 153144 232102 153196
rect 277026 153144 277032 153196
rect 277084 153184 277090 153196
rect 277118 153184 277124 153196
rect 277084 153156 277124 153184
rect 277084 153144 277090 153156
rect 277118 153144 277124 153156
rect 277176 153144 277182 153196
rect 270126 152464 270132 152516
rect 270184 152504 270190 152516
rect 270310 152504 270316 152516
rect 270184 152476 270316 152504
rect 270184 152464 270190 152476
rect 270310 152464 270316 152476
rect 270368 152464 270374 152516
rect 230566 152056 230572 152108
rect 230624 152096 230630 152108
rect 230750 152096 230756 152108
rect 230624 152068 230756 152096
rect 230624 152056 230630 152068
rect 230750 152056 230756 152068
rect 230808 152056 230814 152108
rect 179874 151784 179880 151836
rect 179932 151824 179938 151836
rect 179966 151824 179972 151836
rect 179932 151796 179972 151824
rect 179932 151784 179938 151796
rect 179966 151784 179972 151796
rect 180024 151784 180030 151836
rect 181070 151824 181076 151836
rect 181031 151796 181076 151824
rect 181070 151784 181076 151796
rect 181128 151784 181134 151836
rect 217134 151824 217140 151836
rect 217095 151796 217140 151824
rect 217134 151784 217140 151796
rect 217192 151784 217198 151836
rect 344462 151784 344468 151836
rect 344520 151824 344526 151836
rect 344554 151824 344560 151836
rect 344520 151796 344560 151824
rect 344520 151784 344526 151796
rect 344554 151784 344560 151796
rect 344612 151784 344618 151836
rect 345658 151824 345664 151836
rect 345619 151796 345664 151824
rect 345658 151784 345664 151796
rect 345716 151784 345722 151836
rect 3326 151716 3332 151768
rect 3384 151756 3390 151768
rect 21358 151756 21364 151768
rect 3384 151728 21364 151756
rect 3384 151716 3390 151728
rect 21358 151716 21364 151728
rect 21416 151716 21422 151768
rect 361209 150535 361267 150541
rect 361209 150501 361221 150535
rect 361255 150532 361267 150535
rect 361255 150504 361344 150532
rect 361255 150501 361267 150504
rect 361209 150495 361267 150501
rect 361316 150476 361344 150504
rect 361298 150424 361304 150476
rect 361356 150424 361362 150476
rect 225598 150328 225604 150340
rect 225559 150300 225604 150328
rect 225598 150288 225604 150300
rect 225656 150288 225662 150340
rect 177114 149036 177120 149048
rect 177075 149008 177120 149036
rect 177114 148996 177120 149008
rect 177172 148996 177178 149048
rect 178126 149036 178132 149048
rect 178087 149008 178132 149036
rect 178126 148996 178132 149008
rect 178184 148996 178190 149048
rect 299198 147812 299204 147824
rect 299159 147784 299204 147812
rect 299198 147772 299204 147784
rect 299256 147772 299262 147824
rect 300486 147812 300492 147824
rect 300447 147784 300492 147812
rect 300486 147772 300492 147784
rect 300544 147772 300550 147824
rect 354398 147772 354404 147824
rect 354456 147772 354462 147824
rect 184014 147704 184020 147756
rect 184072 147704 184078 147756
rect 189350 147704 189356 147756
rect 189408 147704 189414 147756
rect 200390 147704 200396 147756
rect 200448 147704 200454 147756
rect 201862 147704 201868 147756
rect 201920 147704 201926 147756
rect 273070 147704 273076 147756
rect 273128 147744 273134 147756
rect 273254 147744 273260 147756
rect 273128 147716 273260 147744
rect 273128 147704 273134 147716
rect 273254 147704 273260 147716
rect 273312 147704 273318 147756
rect 315758 147704 315764 147756
rect 315816 147704 315822 147756
rect 184032 147620 184060 147704
rect 189368 147620 189396 147704
rect 200408 147620 200436 147704
rect 201880 147620 201908 147704
rect 211890 147636 211896 147688
rect 211948 147636 211954 147688
rect 217134 147636 217140 147688
rect 217192 147636 217198 147688
rect 258166 147636 258172 147688
rect 258224 147676 258230 147688
rect 258350 147676 258356 147688
rect 258224 147648 258356 147676
rect 258224 147636 258230 147648
rect 258350 147636 258356 147648
rect 258408 147636 258414 147688
rect 184014 147568 184020 147620
rect 184072 147568 184078 147620
rect 189350 147568 189356 147620
rect 189408 147568 189414 147620
rect 200390 147568 200396 147620
rect 200448 147568 200454 147620
rect 201862 147568 201868 147620
rect 201920 147568 201926 147620
rect 211908 147608 211936 147636
rect 211982 147608 211988 147620
rect 211908 147580 211988 147608
rect 211982 147568 211988 147580
rect 212040 147568 212046 147620
rect 217152 147608 217180 147636
rect 315776 147620 315804 147704
rect 354416 147688 354444 147772
rect 317230 147676 317236 147688
rect 317191 147648 317236 147676
rect 317230 147636 317236 147648
rect 317288 147636 317294 147688
rect 328270 147676 328276 147688
rect 328231 147648 328276 147676
rect 328270 147636 328276 147648
rect 328328 147636 328334 147688
rect 354398 147636 354404 147688
rect 354456 147636 354462 147688
rect 217226 147608 217232 147620
rect 217152 147580 217232 147608
rect 217226 147568 217232 147580
rect 217284 147568 217290 147620
rect 315758 147568 315764 147620
rect 315816 147568 315822 147620
rect 291930 145024 291936 145036
rect 291891 144996 291936 145024
rect 291930 144984 291936 144996
rect 291988 144984 291994 145036
rect 224034 144916 224040 144968
rect 224092 144956 224098 144968
rect 224126 144956 224132 144968
rect 224092 144928 224132 144956
rect 224092 144916 224098 144928
rect 224126 144916 224132 144928
rect 224184 144916 224190 144968
rect 299198 144956 299204 144968
rect 299159 144928 299204 144956
rect 299198 144916 299204 144928
rect 299256 144916 299262 144968
rect 300486 144956 300492 144968
rect 300447 144928 300492 144956
rect 300486 144916 300492 144928
rect 300544 144916 300550 144968
rect 328270 144956 328276 144968
rect 328231 144928 328276 144956
rect 328270 144916 328276 144928
rect 328328 144916 328334 144968
rect 171410 144848 171416 144900
rect 171468 144888 171474 144900
rect 171594 144888 171600 144900
rect 171468 144860 171600 144888
rect 171468 144848 171474 144860
rect 171594 144848 171600 144860
rect 171652 144848 171658 144900
rect 173066 144848 173072 144900
rect 173124 144888 173130 144900
rect 173250 144888 173256 144900
rect 173124 144860 173256 144888
rect 173124 144848 173130 144860
rect 173250 144848 173256 144860
rect 173308 144848 173314 144900
rect 203150 144888 203156 144900
rect 203111 144860 203156 144888
rect 203150 144848 203156 144860
rect 203208 144848 203214 144900
rect 211893 144891 211951 144897
rect 211893 144857 211905 144891
rect 211939 144888 211951 144891
rect 211982 144888 211988 144900
rect 211939 144860 211988 144888
rect 211939 144857 211951 144860
rect 211893 144851 211951 144857
rect 211982 144848 211988 144860
rect 212040 144848 212046 144900
rect 230934 144888 230940 144900
rect 230895 144860 230940 144888
rect 230934 144848 230940 144860
rect 230992 144848 230998 144900
rect 258258 144888 258264 144900
rect 258219 144860 258264 144888
rect 258258 144848 258264 144860
rect 258316 144848 258322 144900
rect 329558 144888 329564 144900
rect 329519 144860 329564 144888
rect 329558 144848 329564 144860
rect 329616 144848 329622 144900
rect 362402 144888 362408 144900
rect 362363 144860 362408 144888
rect 362402 144848 362408 144860
rect 362460 144848 362466 144900
rect 317230 143596 317236 143608
rect 317191 143568 317236 143596
rect 317230 143556 317236 143568
rect 317288 143556 317294 143608
rect 261110 143528 261116 143540
rect 261071 143500 261116 143528
rect 261110 143488 261116 143500
rect 261168 143488 261174 143540
rect 275833 143531 275891 143537
rect 275833 143497 275845 143531
rect 275879 143528 275891 143531
rect 275922 143528 275928 143540
rect 275879 143500 275928 143528
rect 275879 143497 275891 143500
rect 275833 143491 275891 143497
rect 275922 143488 275928 143500
rect 275980 143488 275986 143540
rect 285306 143528 285312 143540
rect 285267 143500 285312 143528
rect 285306 143488 285312 143500
rect 285364 143488 285370 143540
rect 286594 143528 286600 143540
rect 286555 143500 286600 143528
rect 286594 143488 286600 143500
rect 286652 143488 286658 143540
rect 289354 143528 289360 143540
rect 289315 143500 289360 143528
rect 289354 143488 289360 143500
rect 289412 143488 289418 143540
rect 291838 143488 291844 143540
rect 291896 143528 291902 143540
rect 291930 143528 291936 143540
rect 291896 143500 291936 143528
rect 291896 143488 291902 143500
rect 291930 143488 291936 143500
rect 291988 143488 291994 143540
rect 318429 143531 318487 143537
rect 318429 143497 318441 143531
rect 318475 143528 318487 143531
rect 318518 143528 318524 143540
rect 318475 143500 318524 143528
rect 318475 143497 318487 143500
rect 318429 143491 318487 143497
rect 318518 143488 318524 143500
rect 318576 143488 318582 143540
rect 230566 142808 230572 142860
rect 230624 142848 230630 142860
rect 230750 142848 230756 142860
rect 230624 142820 230756 142848
rect 230624 142808 230630 142820
rect 230750 142808 230756 142820
rect 230808 142808 230814 142860
rect 234982 142808 234988 142860
rect 235040 142848 235046 142860
rect 235258 142848 235264 142860
rect 235040 142820 235264 142848
rect 235040 142808 235046 142820
rect 235258 142808 235264 142820
rect 235316 142808 235322 142860
rect 270126 142808 270132 142860
rect 270184 142848 270190 142860
rect 270310 142848 270316 142860
rect 270184 142820 270316 142848
rect 270184 142808 270190 142820
rect 270310 142808 270316 142820
rect 270368 142808 270374 142860
rect 236178 142196 236184 142248
rect 236236 142236 236242 142248
rect 236270 142236 236276 142248
rect 236236 142208 236276 142236
rect 236236 142196 236242 142208
rect 236270 142196 236276 142208
rect 236328 142196 236334 142248
rect 341978 142168 341984 142180
rect 341939 142140 341984 142168
rect 341978 142128 341984 142140
rect 342036 142128 342042 142180
rect 181070 142100 181076 142112
rect 181031 142072 181076 142100
rect 181070 142060 181076 142072
rect 181128 142060 181134 142112
rect 182174 142100 182180 142112
rect 182135 142072 182180 142100
rect 182174 142060 182180 142072
rect 182232 142060 182238 142112
rect 229278 142060 229284 142112
rect 229336 142100 229342 142112
rect 229370 142100 229376 142112
rect 229336 142072 229376 142100
rect 229336 142060 229342 142072
rect 229370 142060 229376 142072
rect 229428 142060 229434 142112
rect 235074 142060 235080 142112
rect 235132 142060 235138 142112
rect 236178 142060 236184 142112
rect 236236 142100 236242 142112
rect 236273 142103 236331 142109
rect 236273 142100 236285 142103
rect 236236 142072 236285 142100
rect 236236 142060 236242 142072
rect 236273 142069 236285 142072
rect 236319 142069 236331 142103
rect 315850 142100 315856 142112
rect 315811 142072 315856 142100
rect 236273 142063 236331 142069
rect 315850 142060 315856 142072
rect 315908 142060 315914 142112
rect 361390 142100 361396 142112
rect 361351 142072 361396 142100
rect 361390 142060 361396 142072
rect 361448 142060 361454 142112
rect 235092 142032 235120 142060
rect 235166 142032 235172 142044
rect 235092 142004 235172 142032
rect 235166 141992 235172 142004
rect 235224 141992 235230 142044
rect 225230 140768 225236 140820
rect 225288 140808 225294 140820
rect 225598 140808 225604 140820
rect 225288 140780 225604 140808
rect 225288 140768 225294 140780
rect 225598 140768 225604 140780
rect 225656 140768 225662 140820
rect 341978 140808 341984 140820
rect 341939 140780 341984 140808
rect 341978 140768 341984 140780
rect 342036 140768 342042 140820
rect 343269 140811 343327 140817
rect 343269 140777 343281 140811
rect 343315 140808 343327 140811
rect 343358 140808 343364 140820
rect 343315 140780 343364 140808
rect 343315 140777 343327 140780
rect 343269 140771 343327 140777
rect 343358 140768 343364 140780
rect 343416 140768 343422 140820
rect 344278 140768 344284 140820
rect 344336 140808 344342 140820
rect 344370 140808 344376 140820
rect 344336 140780 344376 140808
rect 344336 140768 344342 140780
rect 344370 140768 344376 140780
rect 344428 140768 344434 140820
rect 179966 140740 179972 140752
rect 179927 140712 179972 140740
rect 179966 140700 179972 140712
rect 180024 140700 180030 140752
rect 194873 140743 194931 140749
rect 194873 140709 194885 140743
rect 194919 140740 194931 140743
rect 194962 140740 194968 140752
rect 194919 140712 194968 140740
rect 194919 140709 194931 140712
rect 194873 140703 194931 140709
rect 194962 140700 194968 140712
rect 195020 140700 195026 140752
rect 212261 140743 212319 140749
rect 212261 140709 212273 140743
rect 212307 140740 212319 140743
rect 212350 140740 212356 140752
rect 212307 140712 212356 140740
rect 212307 140709 212319 140712
rect 212261 140703 212319 140709
rect 212350 140700 212356 140712
rect 212408 140700 212414 140752
rect 177114 139516 177120 139528
rect 177075 139488 177120 139516
rect 177114 139476 177120 139488
rect 177172 139476 177178 139528
rect 178126 139516 178132 139528
rect 178087 139488 178132 139516
rect 178126 139476 178132 139488
rect 178184 139476 178190 139528
rect 228174 139448 228180 139460
rect 228135 139420 228180 139448
rect 228174 139408 228180 139420
rect 228232 139408 228238 139460
rect 177114 139380 177120 139392
rect 177075 139352 177120 139380
rect 177114 139340 177120 139352
rect 177172 139340 177178 139392
rect 178126 139380 178132 139392
rect 178087 139352 178132 139380
rect 178126 139340 178132 139352
rect 178184 139340 178190 139392
rect 341705 139383 341763 139389
rect 341705 139349 341717 139383
rect 341751 139380 341763 139383
rect 341978 139380 341984 139392
rect 341751 139352 341984 139380
rect 341751 139349 341763 139352
rect 341705 139343 341763 139349
rect 341978 139340 341984 139352
rect 342036 139340 342042 139392
rect 232038 139204 232044 139256
rect 232096 139244 232102 139256
rect 232314 139244 232320 139256
rect 232096 139216 232320 139244
rect 232096 139204 232102 139216
rect 232314 139204 232320 139216
rect 232372 139204 232378 139256
rect 345566 138048 345572 138100
rect 345624 138088 345630 138100
rect 345842 138088 345848 138100
rect 345624 138060 345848 138088
rect 345624 138048 345630 138060
rect 345842 138048 345848 138060
rect 345900 138048 345906 138100
rect 258258 137952 258264 137964
rect 258219 137924 258264 137952
rect 258258 137912 258264 137924
rect 258316 137912 258322 137964
rect 285306 137952 285312 137964
rect 285267 137924 285312 137952
rect 285306 137912 285312 137924
rect 285364 137912 285370 137964
rect 286594 137952 286600 137964
rect 286555 137924 286600 137952
rect 286594 137912 286600 137924
rect 286652 137912 286658 137964
rect 289354 137952 289360 137964
rect 289315 137924 289360 137952
rect 289354 137912 289360 137924
rect 289412 137912 289418 137964
rect 2774 136484 2780 136536
rect 2832 136524 2838 136536
rect 5074 136524 5080 136536
rect 2832 136496 5080 136524
rect 2832 136484 2838 136496
rect 5074 136484 5080 136496
rect 5132 136484 5138 136536
rect 211890 135300 211896 135312
rect 211851 135272 211896 135300
rect 211890 135260 211896 135272
rect 211948 135260 211954 135312
rect 329558 135300 329564 135312
rect 329519 135272 329564 135300
rect 329558 135260 329564 135272
rect 329616 135260 329622 135312
rect 183922 135192 183928 135244
rect 183980 135232 183986 135244
rect 184014 135232 184020 135244
rect 183980 135204 184020 135232
rect 183980 135192 183986 135204
rect 184014 135192 184020 135204
rect 184072 135192 184078 135244
rect 231026 135192 231032 135244
rect 231084 135232 231090 135244
rect 231210 135232 231216 135244
rect 231084 135204 231216 135232
rect 231084 135192 231090 135204
rect 231210 135192 231216 135204
rect 231268 135192 231274 135244
rect 272978 135192 272984 135244
rect 273036 135232 273042 135244
rect 273070 135232 273076 135244
rect 273036 135204 273076 135232
rect 273036 135192 273042 135204
rect 273070 135192 273076 135204
rect 273128 135192 273134 135244
rect 317138 135192 317144 135244
rect 317196 135232 317202 135244
rect 317230 135232 317236 135244
rect 317196 135204 317236 135232
rect 317196 135192 317202 135204
rect 317230 135192 317236 135204
rect 317288 135192 317294 135244
rect 203061 134011 203119 134017
rect 203061 133977 203073 134011
rect 203107 134008 203119 134011
rect 203242 134008 203248 134020
rect 203107 133980 203248 134008
rect 203107 133977 203119 133980
rect 203061 133971 203119 133977
rect 203242 133968 203248 133980
rect 203300 133968 203306 134020
rect 318426 134008 318432 134020
rect 318387 133980 318432 134008
rect 318426 133968 318432 133980
rect 318484 133968 318490 134020
rect 217134 133900 217140 133952
rect 217192 133940 217198 133952
rect 217226 133940 217232 133952
rect 217192 133912 217232 133940
rect 217192 133900 217198 133912
rect 217226 133900 217232 133912
rect 217284 133900 217290 133952
rect 261110 133940 261116 133952
rect 261071 133912 261116 133940
rect 261110 133900 261116 133912
rect 261168 133900 261174 133952
rect 275830 133940 275836 133952
rect 275791 133912 275836 133940
rect 275830 133900 275836 133912
rect 275888 133900 275894 133952
rect 201773 133875 201831 133881
rect 201773 133841 201785 133875
rect 201819 133872 201831 133875
rect 201862 133872 201868 133884
rect 201819 133844 201868 133872
rect 201819 133841 201831 133844
rect 201773 133835 201831 133841
rect 201862 133832 201868 133844
rect 201920 133832 201926 133884
rect 277210 133872 277216 133884
rect 277171 133844 277216 133872
rect 277210 133832 277216 133844
rect 277268 133832 277274 133884
rect 284018 133832 284024 133884
rect 284076 133872 284082 133884
rect 284294 133872 284300 133884
rect 284076 133844 284300 133872
rect 284076 133832 284082 133844
rect 284294 133832 284300 133844
rect 284352 133832 284358 133884
rect 291746 133832 291752 133884
rect 291804 133872 291810 133884
rect 291930 133872 291936 133884
rect 291804 133844 291936 133872
rect 291804 133832 291810 133844
rect 291930 133832 291936 133844
rect 291988 133832 291994 133884
rect 318426 133872 318432 133884
rect 318387 133844 318432 133872
rect 318426 133832 318432 133844
rect 318484 133832 318490 133884
rect 225322 133764 225328 133816
rect 225380 133804 225386 133816
rect 225506 133804 225512 133816
rect 225380 133776 225512 133804
rect 225380 133764 225386 133776
rect 225506 133764 225512 133776
rect 225564 133764 225570 133816
rect 228266 133764 228272 133816
rect 228324 133804 228330 133816
rect 228450 133804 228456 133816
rect 228324 133776 228456 133804
rect 228324 133764 228330 133776
rect 228450 133764 228456 133776
rect 228508 133764 228514 133816
rect 181073 132583 181131 132589
rect 181073 132549 181085 132583
rect 181119 132580 181131 132583
rect 181162 132580 181168 132592
rect 181119 132552 181168 132580
rect 181119 132549 181131 132552
rect 181073 132543 181131 132549
rect 181162 132540 181168 132552
rect 181220 132540 181226 132592
rect 203058 132512 203064 132524
rect 203019 132484 203064 132512
rect 203058 132472 203064 132484
rect 203116 132472 203122 132524
rect 315850 132512 315856 132524
rect 315811 132484 315856 132512
rect 315850 132472 315856 132484
rect 315908 132472 315914 132524
rect 343266 132472 343272 132524
rect 343324 132512 343330 132524
rect 343358 132512 343364 132524
rect 343324 132484 343364 132512
rect 343324 132472 343330 132484
rect 343358 132472 343364 132484
rect 343416 132472 343422 132524
rect 361390 132512 361396 132524
rect 361351 132484 361396 132512
rect 361390 132472 361396 132484
rect 361448 132472 361454 132524
rect 181073 132447 181131 132453
rect 181073 132413 181085 132447
rect 181119 132444 181131 132447
rect 181162 132444 181168 132456
rect 181119 132416 181168 132444
rect 181119 132413 181131 132416
rect 181073 132407 181131 132413
rect 181162 132404 181168 132416
rect 181220 132404 181226 132456
rect 345566 132444 345572 132456
rect 345527 132416 345572 132444
rect 345566 132404 345572 132416
rect 345624 132404 345630 132456
rect 344278 132336 344284 132388
rect 344336 132376 344342 132388
rect 344554 132376 344560 132388
rect 344336 132348 344560 132376
rect 344336 132336 344342 132348
rect 344554 132336 344560 132348
rect 344612 132336 344618 132388
rect 270126 131928 270132 131980
rect 270184 131968 270190 131980
rect 270310 131968 270316 131980
rect 270184 131940 270316 131968
rect 270184 131928 270190 131940
rect 270310 131928 270316 131940
rect 270368 131928 270374 131980
rect 179969 131223 180027 131229
rect 179969 131189 179981 131223
rect 180015 131220 180027 131223
rect 180015 131192 180196 131220
rect 180015 131189 180027 131192
rect 179969 131183 180027 131189
rect 180168 131164 180196 131192
rect 180150 131112 180156 131164
rect 180208 131112 180214 131164
rect 194870 131152 194876 131164
rect 194831 131124 194876 131152
rect 194870 131112 194876 131124
rect 194928 131112 194934 131164
rect 212261 131155 212319 131161
rect 212261 131121 212273 131155
rect 212307 131152 212319 131155
rect 212350 131152 212356 131164
rect 212307 131124 212356 131152
rect 212307 131121 212319 131124
rect 212261 131115 212319 131121
rect 212350 131112 212356 131124
rect 212408 131112 212414 131164
rect 343266 131084 343272 131096
rect 343227 131056 343272 131084
rect 343266 131044 343272 131056
rect 343324 131044 343330 131096
rect 177114 129792 177120 129804
rect 177075 129764 177120 129792
rect 177114 129752 177120 129764
rect 177172 129752 177178 129804
rect 178129 129795 178187 129801
rect 178129 129761 178141 129795
rect 178175 129792 178187 129795
rect 178402 129792 178408 129804
rect 178175 129764 178408 129792
rect 178175 129761 178187 129764
rect 178129 129755 178187 129761
rect 178402 129752 178408 129764
rect 178460 129752 178466 129804
rect 341702 129792 341708 129804
rect 341663 129764 341708 129792
rect 341702 129752 341708 129764
rect 341760 129752 341766 129804
rect 299198 128500 299204 128512
rect 299159 128472 299204 128500
rect 299198 128460 299204 128472
rect 299256 128460 299262 128512
rect 300486 128500 300492 128512
rect 300447 128472 300492 128500
rect 300486 128460 300492 128472
rect 300544 128460 300550 128512
rect 191098 128432 191104 128444
rect 191024 128404 191104 128432
rect 189350 128324 189356 128376
rect 189408 128324 189414 128376
rect 189368 128296 189396 128324
rect 191024 128308 191052 128404
rect 191098 128392 191104 128404
rect 191156 128392 191162 128444
rect 211890 128324 211896 128376
rect 211948 128324 211954 128376
rect 258166 128324 258172 128376
rect 258224 128364 258230 128376
rect 258350 128364 258356 128376
rect 258224 128336 258356 128364
rect 258224 128324 258230 128336
rect 258350 128324 258356 128336
rect 258408 128324 258414 128376
rect 328270 128364 328276 128376
rect 328231 128336 328276 128364
rect 328270 128324 328276 128336
rect 328328 128324 328334 128376
rect 354398 128364 354404 128376
rect 354359 128336 354404 128364
rect 354398 128324 354404 128336
rect 354456 128324 354462 128376
rect 355686 128364 355692 128376
rect 355647 128336 355692 128364
rect 355686 128324 355692 128336
rect 355744 128324 355750 128376
rect 189442 128296 189448 128308
rect 189368 128268 189448 128296
rect 189442 128256 189448 128268
rect 189500 128256 189506 128308
rect 191006 128256 191012 128308
rect 191064 128256 191070 128308
rect 211908 128296 211936 128324
rect 211982 128296 211988 128308
rect 211908 128268 211988 128296
rect 211982 128256 211988 128268
rect 212040 128256 212046 128308
rect 179966 127644 179972 127696
rect 180024 127684 180030 127696
rect 180150 127684 180156 127696
rect 180024 127656 180156 127684
rect 180024 127644 180030 127656
rect 180150 127644 180156 127656
rect 180208 127644 180214 127696
rect 362310 127644 362316 127696
rect 362368 127684 362374 127696
rect 362586 127684 362592 127696
rect 362368 127656 362592 127684
rect 362368 127644 362374 127656
rect 362586 127644 362592 127656
rect 362644 127644 362650 127696
rect 285306 125604 285312 125656
rect 285364 125644 285370 125656
rect 285398 125644 285404 125656
rect 285364 125616 285404 125644
rect 285364 125604 285370 125616
rect 285398 125604 285404 125616
rect 285456 125604 285462 125656
rect 286594 125604 286600 125656
rect 286652 125644 286658 125656
rect 286686 125644 286692 125656
rect 286652 125616 286692 125644
rect 286652 125604 286658 125616
rect 286686 125604 286692 125616
rect 286744 125604 286750 125656
rect 289354 125604 289360 125656
rect 289412 125644 289418 125656
rect 289446 125644 289452 125656
rect 289412 125616 289452 125644
rect 289412 125604 289418 125616
rect 289446 125604 289452 125616
rect 289504 125604 289510 125656
rect 171410 125576 171416 125588
rect 171371 125548 171416 125576
rect 171410 125536 171416 125548
rect 171468 125536 171474 125588
rect 173066 125576 173072 125588
rect 173027 125548 173072 125576
rect 173066 125536 173072 125548
rect 173124 125536 173130 125588
rect 183922 125536 183928 125588
rect 183980 125576 183986 125588
rect 184106 125576 184112 125588
rect 183980 125548 184112 125576
rect 183980 125536 183986 125548
rect 184106 125536 184112 125548
rect 184164 125536 184170 125588
rect 191006 125536 191012 125588
rect 191064 125576 191070 125588
rect 191190 125576 191196 125588
rect 191064 125548 191196 125576
rect 191064 125536 191070 125548
rect 191190 125536 191196 125548
rect 191248 125536 191254 125588
rect 211893 125579 211951 125585
rect 211893 125545 211905 125579
rect 211939 125576 211951 125579
rect 211982 125576 211988 125588
rect 211939 125548 211988 125576
rect 211939 125545 211951 125548
rect 211893 125539 211951 125545
rect 211982 125536 211988 125548
rect 212040 125536 212046 125588
rect 235074 125536 235080 125588
rect 235132 125536 235138 125588
rect 258258 125576 258264 125588
rect 258219 125548 258264 125576
rect 258258 125536 258264 125548
rect 258316 125536 258322 125588
rect 318426 125576 318432 125588
rect 318387 125548 318432 125576
rect 318426 125536 318432 125548
rect 318484 125536 318490 125588
rect 329558 125576 329564 125588
rect 329519 125548 329564 125576
rect 329558 125536 329564 125548
rect 329616 125536 329622 125588
rect 355778 125536 355784 125588
rect 355836 125536 355842 125588
rect 235092 125508 235120 125536
rect 235166 125508 235172 125520
rect 235092 125480 235172 125508
rect 235166 125468 235172 125480
rect 235224 125468 235230 125520
rect 355796 125452 355824 125536
rect 355778 125400 355784 125452
rect 355836 125400 355842 125452
rect 182174 124176 182180 124228
rect 182232 124216 182238 124228
rect 182232 124188 182277 124216
rect 182232 124176 182238 124188
rect 194870 124176 194876 124228
rect 194928 124216 194934 124228
rect 194962 124216 194968 124228
rect 194928 124188 194968 124216
rect 194928 124176 194934 124188
rect 194962 124176 194968 124188
rect 195020 124176 195026 124228
rect 201770 124216 201776 124228
rect 201731 124188 201776 124216
rect 201770 124176 201776 124188
rect 201828 124176 201834 124228
rect 232222 124176 232228 124228
rect 232280 124216 232286 124228
rect 232314 124216 232320 124228
rect 232280 124188 232320 124216
rect 232280 124176 232286 124188
rect 232314 124176 232320 124188
rect 232372 124176 232378 124228
rect 277210 124216 277216 124228
rect 277171 124188 277216 124216
rect 277210 124176 277216 124188
rect 277268 124176 277274 124228
rect 299198 124216 299204 124228
rect 299159 124188 299204 124216
rect 299198 124176 299204 124188
rect 299256 124176 299262 124228
rect 300486 124216 300492 124228
rect 300447 124188 300492 124216
rect 300486 124176 300492 124188
rect 300544 124176 300550 124228
rect 328270 124216 328276 124228
rect 328231 124188 328276 124216
rect 328270 124176 328276 124188
rect 328328 124176 328334 124228
rect 354398 124216 354404 124228
rect 354359 124188 354404 124216
rect 354398 124176 354404 124188
rect 354456 124176 354462 124228
rect 355686 124216 355692 124228
rect 355647 124188 355692 124216
rect 355686 124176 355692 124188
rect 355744 124176 355750 124228
rect 361298 124176 361304 124228
rect 361356 124216 361362 124228
rect 361390 124216 361396 124228
rect 361356 124188 361396 124216
rect 361356 124176 361362 124188
rect 361390 124176 361396 124188
rect 361448 124176 361454 124228
rect 192202 124108 192208 124160
rect 192260 124148 192266 124160
rect 192294 124148 192300 124160
rect 192260 124120 192300 124148
rect 192260 124108 192266 124120
rect 192294 124108 192300 124120
rect 192352 124108 192358 124160
rect 200298 124148 200304 124160
rect 200259 124120 200304 124148
rect 200298 124108 200304 124120
rect 200356 124108 200362 124160
rect 203058 124148 203064 124160
rect 203019 124120 203064 124148
rect 203058 124108 203064 124120
rect 203116 124108 203122 124160
rect 231029 124151 231087 124157
rect 231029 124117 231041 124151
rect 231075 124148 231087 124151
rect 231118 124148 231124 124160
rect 231075 124120 231124 124148
rect 231075 124117 231087 124120
rect 231029 124111 231087 124117
rect 231118 124108 231124 124120
rect 231176 124108 231182 124160
rect 261110 124148 261116 124160
rect 261071 124120 261116 124148
rect 261110 124108 261116 124120
rect 261168 124108 261174 124160
rect 275922 124108 275928 124160
rect 275980 124148 275986 124160
rect 276014 124148 276020 124160
rect 275980 124120 276020 124148
rect 275980 124108 275986 124120
rect 276014 124108 276020 124120
rect 276072 124108 276078 124160
rect 291930 124148 291936 124160
rect 291891 124120 291936 124148
rect 291930 124108 291936 124120
rect 291988 124108 291994 124160
rect 318518 124148 318524 124160
rect 318479 124120 318524 124148
rect 318518 124108 318524 124120
rect 318576 124108 318582 124160
rect 270126 123496 270132 123548
rect 270184 123536 270190 123548
rect 270310 123536 270316 123548
rect 270184 123508 270316 123536
rect 270184 123496 270190 123508
rect 270310 123496 270316 123508
rect 270368 123496 270374 123548
rect 181070 122856 181076 122868
rect 181031 122828 181076 122856
rect 181070 122816 181076 122828
rect 181128 122816 181134 122868
rect 345566 122856 345572 122868
rect 345527 122828 345572 122856
rect 345566 122816 345572 122828
rect 345624 122816 345630 122868
rect 182174 122788 182180 122800
rect 182135 122760 182180 122788
rect 182174 122748 182180 122760
rect 182232 122748 182238 122800
rect 192294 122788 192300 122800
rect 192255 122760 192300 122788
rect 192294 122748 192300 122760
rect 192352 122748 192358 122800
rect 225230 122748 225236 122800
rect 225288 122788 225294 122800
rect 225322 122788 225328 122800
rect 225288 122760 225328 122788
rect 225288 122748 225294 122760
rect 225322 122748 225328 122760
rect 225380 122748 225386 122800
rect 229189 122791 229247 122797
rect 229189 122757 229201 122791
rect 229235 122788 229247 122791
rect 229278 122788 229284 122800
rect 229235 122760 229284 122788
rect 229235 122757 229247 122760
rect 229189 122751 229247 122757
rect 229278 122748 229284 122760
rect 229336 122748 229342 122800
rect 232225 122791 232283 122797
rect 232225 122757 232237 122791
rect 232271 122788 232283 122791
rect 232314 122788 232320 122800
rect 232271 122760 232320 122788
rect 232271 122757 232283 122760
rect 232225 122751 232283 122757
rect 232314 122748 232320 122760
rect 232372 122748 232378 122800
rect 344462 122748 344468 122800
rect 344520 122788 344526 122800
rect 344554 122788 344560 122800
rect 344520 122760 344560 122788
rect 344520 122748 344526 122760
rect 344554 122748 344560 122760
rect 344612 122748 344618 122800
rect 181070 122680 181076 122732
rect 181128 122720 181134 122732
rect 181165 122723 181223 122729
rect 181165 122720 181177 122723
rect 181128 122692 181177 122720
rect 181128 122680 181134 122692
rect 181165 122689 181177 122692
rect 181211 122689 181223 122723
rect 181165 122683 181223 122689
rect 2774 122272 2780 122324
rect 2832 122312 2838 122324
rect 4982 122312 4988 122324
rect 2832 122284 4988 122312
rect 2832 122272 2838 122284
rect 4982 122272 4988 122284
rect 5040 122272 5046 122324
rect 343266 121496 343272 121508
rect 343227 121468 343272 121496
rect 343266 121456 343272 121468
rect 343324 121456 343330 121508
rect 180981 121431 181039 121437
rect 180981 121397 180993 121431
rect 181027 121428 181039 121431
rect 181165 121431 181223 121437
rect 181165 121428 181177 121431
rect 181027 121400 181177 121428
rect 181027 121397 181039 121400
rect 180981 121391 181039 121397
rect 181165 121397 181177 121400
rect 181211 121397 181223 121431
rect 181165 121391 181223 121397
rect 212261 121431 212319 121437
rect 212261 121397 212273 121431
rect 212307 121428 212319 121431
rect 212350 121428 212356 121440
rect 212307 121400 212356 121428
rect 212307 121397 212319 121400
rect 212261 121391 212319 121397
rect 212350 121388 212356 121400
rect 212408 121388 212414 121440
rect 362310 121428 362316 121440
rect 362271 121400 362316 121428
rect 362310 121388 362316 121400
rect 362368 121388 362374 121440
rect 236270 120680 236276 120692
rect 236231 120652 236276 120680
rect 236270 120640 236276 120652
rect 236328 120640 236334 120692
rect 178310 120068 178316 120080
rect 178271 120040 178316 120068
rect 178310 120028 178316 120040
rect 178368 120028 178374 120080
rect 277210 118776 277216 118788
rect 277171 118748 277216 118776
rect 277210 118736 277216 118748
rect 277268 118736 277274 118788
rect 315850 118776 315856 118788
rect 315811 118748 315856 118776
rect 315850 118736 315856 118748
rect 315908 118736 315914 118788
rect 235258 118708 235264 118720
rect 235219 118680 235264 118708
rect 235258 118668 235264 118680
rect 235316 118668 235322 118720
rect 258258 118640 258264 118652
rect 258219 118612 258264 118640
rect 258258 118600 258264 118612
rect 258316 118600 258322 118652
rect 182174 118028 182180 118040
rect 182135 118000 182180 118028
rect 182174 117988 182180 118000
rect 182232 117988 182238 118040
rect 229189 118031 229247 118037
rect 229189 117997 229201 118031
rect 229235 118028 229247 118031
rect 229278 118028 229284 118040
rect 229235 118000 229284 118028
rect 229235 117997 229247 118000
rect 229189 117991 229247 117997
rect 229278 117988 229284 118000
rect 229336 117988 229342 118040
rect 171410 115988 171416 116000
rect 171371 115960 171416 115988
rect 171410 115948 171416 115960
rect 171468 115948 171474 116000
rect 173066 115988 173072 116000
rect 173027 115960 173072 115988
rect 173066 115948 173072 115960
rect 173124 115948 173130 116000
rect 194962 115988 194968 116000
rect 194888 115960 194968 115988
rect 194888 115932 194916 115960
rect 194962 115948 194968 115960
rect 195020 115948 195026 116000
rect 201770 115948 201776 116000
rect 201828 115988 201834 116000
rect 201862 115988 201868 116000
rect 201828 115960 201868 115988
rect 201828 115948 201834 115960
rect 201862 115948 201868 115960
rect 201920 115948 201926 116000
rect 211890 115988 211896 116000
rect 211851 115960 211896 115988
rect 211890 115948 211896 115960
rect 211948 115948 211954 116000
rect 235258 115988 235264 116000
rect 235219 115960 235264 115988
rect 235258 115948 235264 115960
rect 235316 115948 235322 116000
rect 282733 115991 282791 115997
rect 282733 115957 282745 115991
rect 282779 115988 282791 115991
rect 282822 115988 282828 116000
rect 282779 115960 282828 115988
rect 282779 115957 282791 115960
rect 282733 115951 282791 115957
rect 282822 115948 282828 115960
rect 282880 115948 282886 116000
rect 329558 115988 329564 116000
rect 329519 115960 329564 115988
rect 329558 115948 329564 115960
rect 329616 115948 329622 116000
rect 361206 115948 361212 116000
rect 361264 115988 361270 116000
rect 361298 115988 361304 116000
rect 361264 115960 361304 115988
rect 361264 115948 361270 115960
rect 361298 115948 361304 115960
rect 361356 115948 361362 116000
rect 184014 115920 184020 115932
rect 183975 115892 184020 115920
rect 184014 115880 184020 115892
rect 184072 115880 184078 115932
rect 189350 115880 189356 115932
rect 189408 115920 189414 115932
rect 189442 115920 189448 115932
rect 189408 115892 189448 115920
rect 189408 115880 189414 115892
rect 189442 115880 189448 115892
rect 189500 115880 189506 115932
rect 194870 115880 194876 115932
rect 194928 115880 194934 115932
rect 273070 115920 273076 115932
rect 273031 115892 273076 115920
rect 273070 115880 273076 115892
rect 273128 115880 273134 115932
rect 286410 115880 286416 115932
rect 286468 115920 286474 115932
rect 286686 115920 286692 115932
rect 286468 115892 286692 115920
rect 286468 115880 286474 115892
rect 286686 115880 286692 115892
rect 286744 115880 286750 115932
rect 289170 115880 289176 115932
rect 289228 115920 289234 115932
rect 289446 115920 289452 115932
rect 289228 115892 289452 115920
rect 289228 115880 289234 115892
rect 289446 115880 289452 115892
rect 289504 115880 289510 115932
rect 362310 115920 362316 115932
rect 362271 115892 362316 115920
rect 362310 115880 362316 115892
rect 362368 115880 362374 115932
rect 200301 115855 200359 115861
rect 200301 115821 200313 115855
rect 200347 115852 200359 115855
rect 200574 115852 200580 115864
rect 200347 115824 200580 115852
rect 200347 115821 200359 115824
rect 200301 115815 200359 115821
rect 200574 115812 200580 115824
rect 200632 115812 200638 115864
rect 354217 114631 354275 114637
rect 354217 114597 354229 114631
rect 354263 114628 354275 114631
rect 354398 114628 354404 114640
rect 354263 114600 354404 114628
rect 354263 114597 354275 114600
rect 354217 114591 354275 114597
rect 354398 114588 354404 114600
rect 354456 114588 354462 114640
rect 203061 114563 203119 114569
rect 203061 114529 203073 114563
rect 203107 114560 203119 114563
rect 203242 114560 203248 114572
rect 203107 114532 203248 114560
rect 203107 114529 203119 114532
rect 203061 114523 203119 114529
rect 203242 114520 203248 114532
rect 203300 114520 203306 114572
rect 231026 114560 231032 114572
rect 230987 114532 231032 114560
rect 231026 114520 231032 114532
rect 231084 114520 231090 114572
rect 261110 114560 261116 114572
rect 261071 114532 261116 114560
rect 261110 114520 261116 114532
rect 261168 114520 261174 114572
rect 277213 114563 277271 114569
rect 277213 114529 277225 114563
rect 277259 114529 277271 114563
rect 282730 114560 282736 114572
rect 282691 114532 282736 114560
rect 277213 114523 277271 114529
rect 194870 114492 194876 114504
rect 194831 114464 194876 114492
rect 194870 114452 194876 114464
rect 194928 114452 194934 114504
rect 201862 114492 201868 114504
rect 201823 114464 201868 114492
rect 201862 114452 201868 114464
rect 201920 114452 201926 114504
rect 277228 114433 277256 114523
rect 282730 114520 282736 114532
rect 282788 114520 282794 114572
rect 291930 114560 291936 114572
rect 291891 114532 291936 114560
rect 291930 114520 291936 114532
rect 291988 114520 291994 114572
rect 315850 114560 315856 114572
rect 315811 114532 315856 114560
rect 315850 114520 315856 114532
rect 315908 114520 315914 114572
rect 318518 114560 318524 114572
rect 318479 114532 318524 114560
rect 318518 114520 318524 114532
rect 318576 114520 318582 114572
rect 328178 114520 328184 114572
rect 328236 114560 328242 114572
rect 328270 114560 328276 114572
rect 328236 114532 328276 114560
rect 328236 114520 328242 114532
rect 328270 114520 328276 114532
rect 328328 114520 328334 114572
rect 277213 114427 277271 114433
rect 277213 114393 277225 114427
rect 277259 114393 277271 114427
rect 277213 114387 277271 114393
rect 230750 113840 230756 113892
rect 230808 113880 230814 113892
rect 230934 113880 230940 113892
rect 230808 113852 230940 113880
rect 230808 113840 230814 113852
rect 230934 113840 230940 113852
rect 230992 113840 230998 113892
rect 270126 113840 270132 113892
rect 270184 113880 270190 113892
rect 270310 113880 270316 113892
rect 270184 113852 270316 113880
rect 270184 113840 270190 113852
rect 270310 113840 270316 113852
rect 270368 113840 270374 113892
rect 232222 113200 232228 113212
rect 232183 113172 232228 113200
rect 232222 113160 232228 113172
rect 232280 113160 232286 113212
rect 341794 113160 341800 113212
rect 341852 113200 341858 113212
rect 341886 113200 341892 113212
rect 341852 113172 341892 113200
rect 341852 113160 341858 113172
rect 341886 113160 341892 113172
rect 341944 113160 341950 113212
rect 354214 113200 354220 113212
rect 354175 113172 354220 113200
rect 354214 113160 354220 113172
rect 354272 113160 354278 113212
rect 212261 113135 212319 113141
rect 212261 113101 212273 113135
rect 212307 113132 212319 113135
rect 212350 113132 212356 113144
rect 212307 113104 212356 113132
rect 212307 113101 212319 113104
rect 212261 113095 212319 113101
rect 212350 113092 212356 113104
rect 212408 113092 212414 113144
rect 219805 113135 219863 113141
rect 219805 113101 219817 113135
rect 219851 113132 219863 113135
rect 219894 113132 219900 113144
rect 219851 113104 219900 113132
rect 219851 113101 219863 113104
rect 219805 113095 219863 113101
rect 219894 113092 219900 113104
rect 219952 113092 219958 113144
rect 355594 113132 355600 113144
rect 355555 113104 355600 113132
rect 355594 113092 355600 113104
rect 355652 113092 355658 113144
rect 341886 113064 341892 113076
rect 341847 113036 341892 113064
rect 341886 113024 341892 113036
rect 341944 113024 341950 113076
rect 180981 111911 181039 111917
rect 180981 111877 180993 111911
rect 181027 111908 181039 111911
rect 181070 111908 181076 111920
rect 181027 111880 181076 111908
rect 181027 111877 181039 111880
rect 180981 111871 181039 111877
rect 181070 111868 181076 111880
rect 181128 111868 181134 111920
rect 217042 111800 217048 111852
rect 217100 111840 217106 111852
rect 217226 111840 217232 111852
rect 217100 111812 217232 111840
rect 217100 111800 217106 111812
rect 217226 111800 217232 111812
rect 217284 111800 217290 111852
rect 181070 111772 181076 111784
rect 181031 111744 181076 111772
rect 181070 111732 181076 111744
rect 181128 111732 181134 111784
rect 217042 111704 217048 111716
rect 217003 111676 217048 111704
rect 217042 111664 217048 111676
rect 217100 111664 217106 111716
rect 230750 111052 230756 111104
rect 230808 111092 230814 111104
rect 231026 111092 231032 111104
rect 230808 111064 231032 111092
rect 230808 111052 230814 111064
rect 231026 111052 231032 111064
rect 231084 111052 231090 111104
rect 176930 110440 176936 110492
rect 176988 110480 176994 110492
rect 177114 110480 177120 110492
rect 176988 110452 177120 110480
rect 176988 110440 176994 110452
rect 177114 110440 177120 110452
rect 177172 110440 177178 110492
rect 178313 110483 178371 110489
rect 178313 110449 178325 110483
rect 178359 110480 178371 110483
rect 178494 110480 178500 110492
rect 178359 110452 178500 110480
rect 178359 110449 178371 110452
rect 178313 110443 178371 110449
rect 178494 110440 178500 110452
rect 178552 110440 178558 110492
rect 192297 110415 192355 110421
rect 192297 110381 192309 110415
rect 192343 110412 192355 110415
rect 192386 110412 192392 110424
rect 192343 110384 192392 110412
rect 192343 110381 192355 110384
rect 192297 110375 192355 110381
rect 192386 110372 192392 110384
rect 192444 110372 192450 110424
rect 317230 109732 317236 109744
rect 317191 109704 317236 109732
rect 317230 109692 317236 109704
rect 317288 109692 317294 109744
rect 354214 109692 354220 109744
rect 354272 109732 354278 109744
rect 354401 109735 354459 109741
rect 354401 109732 354413 109735
rect 354272 109704 354413 109732
rect 354272 109692 354278 109704
rect 354401 109701 354413 109704
rect 354447 109701 354459 109735
rect 354401 109695 354459 109701
rect 318337 109395 318395 109401
rect 318337 109361 318349 109395
rect 318383 109392 318395 109395
rect 318518 109392 318524 109404
rect 318383 109364 318524 109392
rect 318383 109361 318395 109364
rect 318337 109355 318395 109361
rect 318518 109352 318524 109364
rect 318576 109352 318582 109404
rect 300486 109188 300492 109200
rect 300447 109160 300492 109188
rect 300486 109148 300492 109160
rect 300544 109148 300550 109200
rect 236362 109120 236368 109132
rect 236288 109092 236368 109120
rect 182174 109012 182180 109064
rect 182232 109012 182238 109064
rect 211890 109012 211896 109064
rect 211948 109012 211954 109064
rect 3326 108944 3332 108996
rect 3384 108984 3390 108996
rect 28258 108984 28264 108996
rect 3384 108956 28264 108984
rect 3384 108944 3390 108956
rect 28258 108944 28264 108956
rect 28316 108944 28322 108996
rect 182192 108928 182220 109012
rect 211908 108984 211936 109012
rect 236288 108996 236316 109092
rect 236362 109080 236368 109092
rect 236420 109080 236426 109132
rect 285398 109120 285404 109132
rect 285324 109092 285404 109120
rect 258166 109012 258172 109064
rect 258224 109052 258230 109064
rect 258350 109052 258356 109064
rect 258224 109024 258356 109052
rect 258224 109012 258230 109024
rect 258350 109012 258356 109024
rect 258408 109012 258414 109064
rect 285324 108996 285352 109092
rect 285398 109080 285404 109092
rect 285456 109080 285462 109132
rect 315850 109120 315856 109132
rect 315811 109092 315856 109120
rect 315850 109080 315856 109092
rect 315908 109080 315914 109132
rect 328270 109012 328276 109064
rect 328328 109012 328334 109064
rect 211982 108984 211988 108996
rect 211908 108956 211988 108984
rect 211982 108944 211988 108956
rect 212040 108944 212046 108996
rect 236270 108944 236276 108996
rect 236328 108944 236334 108996
rect 285306 108944 285312 108996
rect 285364 108944 285370 108996
rect 328288 108928 328316 109012
rect 182174 108876 182180 108928
rect 182232 108876 182238 108928
rect 328270 108876 328276 108928
rect 328328 108876 328334 108928
rect 184017 108851 184075 108857
rect 184017 108817 184029 108851
rect 184063 108848 184075 108851
rect 184106 108848 184112 108860
rect 184063 108820 184112 108848
rect 184063 108817 184075 108820
rect 184017 108811 184075 108817
rect 184106 108808 184112 108820
rect 184164 108808 184170 108860
rect 178126 106904 178132 106956
rect 178184 106944 178190 106956
rect 178494 106944 178500 106956
rect 178184 106916 178500 106944
rect 178184 106904 178190 106916
rect 178494 106904 178500 106916
rect 178552 106904 178558 106956
rect 273070 106332 273076 106344
rect 273031 106304 273076 106332
rect 273070 106292 273076 106304
rect 273128 106292 273134 106344
rect 171410 106264 171416 106276
rect 171371 106236 171416 106264
rect 171410 106224 171416 106236
rect 171468 106224 171474 106276
rect 173066 106264 173072 106276
rect 173027 106236 173072 106264
rect 173066 106224 173072 106236
rect 173124 106224 173130 106276
rect 211893 106267 211951 106273
rect 211893 106233 211905 106267
rect 211939 106264 211951 106267
rect 211982 106264 211988 106276
rect 211939 106236 211988 106264
rect 211939 106233 211951 106236
rect 211893 106227 211951 106233
rect 211982 106224 211988 106236
rect 212040 106224 212046 106276
rect 235074 106224 235080 106276
rect 235132 106224 235138 106276
rect 236270 106264 236276 106276
rect 236231 106236 236276 106264
rect 236270 106224 236276 106236
rect 236328 106224 236334 106276
rect 258258 106264 258264 106276
rect 258219 106236 258264 106264
rect 258258 106224 258264 106236
rect 258316 106224 258322 106276
rect 329558 106264 329564 106276
rect 329519 106236 329564 106264
rect 329558 106224 329564 106236
rect 329616 106224 329622 106276
rect 235092 106196 235120 106224
rect 235166 106196 235172 106208
rect 235092 106168 235172 106196
rect 235166 106156 235172 106168
rect 235224 106156 235230 106208
rect 270126 105408 270132 105460
rect 270184 105448 270190 105460
rect 270310 105448 270316 105460
rect 270184 105420 270316 105448
rect 270184 105408 270190 105420
rect 270310 105408 270316 105420
rect 270368 105408 270374 105460
rect 277210 104972 277216 104984
rect 277171 104944 277216 104972
rect 277210 104932 277216 104944
rect 277268 104932 277274 104984
rect 176930 104864 176936 104916
rect 176988 104904 176994 104916
rect 177022 104904 177028 104916
rect 176988 104876 177028 104904
rect 176988 104864 176994 104876
rect 177022 104864 177028 104876
rect 177080 104864 177086 104916
rect 194873 104907 194931 104913
rect 194873 104873 194885 104907
rect 194919 104904 194931 104907
rect 194962 104904 194968 104916
rect 194919 104876 194968 104904
rect 194919 104873 194931 104876
rect 194873 104867 194931 104873
rect 194962 104864 194968 104876
rect 195020 104864 195026 104916
rect 201865 104907 201923 104913
rect 201865 104873 201877 104907
rect 201911 104904 201923 104907
rect 202046 104904 202052 104916
rect 201911 104876 202052 104904
rect 201911 104873 201923 104876
rect 201865 104867 201923 104873
rect 202046 104864 202052 104876
rect 202104 104864 202110 104916
rect 315850 104904 315856 104916
rect 315811 104876 315856 104904
rect 315850 104864 315856 104876
rect 315908 104864 315914 104916
rect 318334 104904 318340 104916
rect 318295 104876 318340 104904
rect 318334 104864 318340 104876
rect 318392 104864 318398 104916
rect 261110 104836 261116 104848
rect 261071 104808 261116 104836
rect 261110 104796 261116 104808
rect 261168 104796 261174 104848
rect 275833 104839 275891 104845
rect 275833 104805 275845 104839
rect 275879 104836 275891 104839
rect 275922 104836 275928 104848
rect 275879 104808 275928 104836
rect 275879 104805 275891 104808
rect 275833 104799 275891 104805
rect 275922 104796 275928 104808
rect 275980 104796 275986 104848
rect 277121 104839 277179 104845
rect 277121 104805 277133 104839
rect 277167 104836 277179 104839
rect 277210 104836 277216 104848
rect 277167 104808 277216 104836
rect 277167 104805 277179 104808
rect 277121 104799 277179 104805
rect 277210 104796 277216 104808
rect 277268 104796 277274 104848
rect 282730 104836 282736 104848
rect 282691 104808 282736 104836
rect 282730 104796 282736 104808
rect 282788 104796 282794 104848
rect 283929 104839 283987 104845
rect 283929 104805 283941 104839
rect 283975 104836 283987 104839
rect 284018 104836 284024 104848
rect 283975 104808 284024 104836
rect 283975 104805 283987 104808
rect 283929 104799 283987 104805
rect 284018 104796 284024 104808
rect 284076 104796 284082 104848
rect 182174 104728 182180 104780
rect 182232 104768 182238 104780
rect 182232 104740 182277 104768
rect 182232 104728 182238 104740
rect 230750 104184 230756 104236
rect 230808 104224 230814 104236
rect 230934 104224 230940 104236
rect 230808 104196 230940 104224
rect 230808 104184 230814 104196
rect 230934 104184 230940 104196
rect 230992 104184 230998 104236
rect 219802 103612 219808 103624
rect 219763 103584 219808 103612
rect 219802 103572 219808 103584
rect 219860 103572 219866 103624
rect 299198 103544 299204 103556
rect 299159 103516 299204 103544
rect 299198 103504 299204 103516
rect 299256 103504 299262 103556
rect 300486 103544 300492 103556
rect 300447 103516 300492 103544
rect 300486 103504 300492 103516
rect 300544 103504 300550 103556
rect 341889 103547 341947 103553
rect 341889 103513 341901 103547
rect 341935 103544 341947 103547
rect 341978 103544 341984 103556
rect 341935 103516 341984 103544
rect 341935 103513 341947 103516
rect 341889 103507 341947 103513
rect 341978 103504 341984 103516
rect 342036 103504 342042 103556
rect 355597 103547 355655 103553
rect 355597 103513 355609 103547
rect 355643 103544 355655 103547
rect 355686 103544 355692 103556
rect 355643 103516 355692 103544
rect 355643 103513 355655 103516
rect 355597 103507 355655 103513
rect 355686 103504 355692 103516
rect 355744 103504 355750 103556
rect 219713 103479 219771 103485
rect 219713 103445 219725 103479
rect 219759 103476 219771 103479
rect 219802 103476 219808 103488
rect 219759 103448 219808 103476
rect 219759 103445 219771 103448
rect 219713 103439 219771 103445
rect 219802 103436 219808 103448
rect 219860 103436 219866 103488
rect 344465 103479 344523 103485
rect 344465 103445 344477 103479
rect 344511 103476 344523 103479
rect 344554 103476 344560 103488
rect 344511 103448 344560 103476
rect 344511 103445 344523 103448
rect 344465 103439 344523 103445
rect 344554 103436 344560 103448
rect 344612 103436 344618 103488
rect 181070 102252 181076 102264
rect 181031 102224 181076 102252
rect 181070 102212 181076 102224
rect 181128 102212 181134 102264
rect 299198 102252 299204 102264
rect 299159 102224 299204 102252
rect 299198 102212 299204 102224
rect 299256 102212 299262 102264
rect 217045 102187 217103 102193
rect 217045 102153 217057 102187
rect 217091 102184 217103 102187
rect 217226 102184 217232 102196
rect 217091 102156 217232 102184
rect 217091 102153 217103 102156
rect 217045 102147 217103 102153
rect 217226 102144 217232 102156
rect 217284 102144 217290 102196
rect 177022 102116 177028 102128
rect 176983 102088 177028 102116
rect 177022 102076 177028 102088
rect 177080 102076 177086 102128
rect 179966 102116 179972 102128
rect 179927 102088 179972 102116
rect 179966 102076 179972 102088
rect 180024 102076 180030 102128
rect 181070 102076 181076 102128
rect 181128 102116 181134 102128
rect 181438 102116 181444 102128
rect 181128 102088 181444 102116
rect 181128 102076 181134 102088
rect 181438 102076 181444 102088
rect 181496 102076 181502 102128
rect 298922 102076 298928 102128
rect 298980 102116 298986 102128
rect 299198 102116 299204 102128
rect 298980 102088 299204 102116
rect 298980 102076 298986 102088
rect 299198 102076 299204 102088
rect 299256 102076 299262 102128
rect 177942 102008 177948 102060
rect 178000 102048 178006 102060
rect 178126 102048 178132 102060
rect 178000 102020 178132 102048
rect 178000 102008 178006 102020
rect 178126 102008 178132 102020
rect 178184 102008 178190 102060
rect 211893 100079 211951 100085
rect 211893 100045 211905 100079
rect 211939 100076 211951 100079
rect 211982 100076 211988 100088
rect 211939 100048 211988 100076
rect 211939 100045 211951 100048
rect 211893 100039 211951 100045
rect 211982 100036 211988 100048
rect 212040 100036 212046 100088
rect 225322 99668 225328 99680
rect 225283 99640 225328 99668
rect 225322 99628 225328 99640
rect 225380 99628 225386 99680
rect 224034 99532 224040 99544
rect 223995 99504 224040 99532
rect 224034 99492 224040 99504
rect 224092 99492 224098 99544
rect 235258 99396 235264 99408
rect 235219 99368 235264 99396
rect 235258 99356 235264 99368
rect 235316 99356 235322 99408
rect 182177 99331 182235 99337
rect 182177 99297 182189 99331
rect 182223 99328 182235 99331
rect 182266 99328 182272 99340
rect 182223 99300 182272 99328
rect 182223 99297 182235 99300
rect 182177 99291 182235 99297
rect 182266 99288 182272 99300
rect 182324 99288 182330 99340
rect 258258 99328 258264 99340
rect 258219 99300 258264 99328
rect 258258 99288 258264 99300
rect 258316 99288 258322 99340
rect 315758 96948 315764 96960
rect 315719 96920 315764 96948
rect 315758 96908 315764 96920
rect 315816 96908 315822 96960
rect 171410 96676 171416 96688
rect 171371 96648 171416 96676
rect 171410 96636 171416 96648
rect 171468 96636 171474 96688
rect 173066 96676 173072 96688
rect 173027 96648 173072 96676
rect 173066 96636 173072 96648
rect 173124 96636 173130 96688
rect 235258 96676 235264 96688
rect 235219 96648 235264 96676
rect 235258 96636 235264 96648
rect 235316 96636 235322 96688
rect 236273 96679 236331 96685
rect 236273 96645 236285 96679
rect 236319 96676 236331 96679
rect 236362 96676 236368 96688
rect 236319 96648 236368 96676
rect 236319 96645 236331 96648
rect 236273 96639 236331 96645
rect 236362 96636 236368 96648
rect 236420 96636 236426 96688
rect 291930 96636 291936 96688
rect 291988 96676 291994 96688
rect 292022 96676 292028 96688
rect 291988 96648 292028 96676
rect 291988 96636 291994 96648
rect 292022 96636 292028 96648
rect 292080 96636 292086 96688
rect 317230 96676 317236 96688
rect 317191 96648 317236 96676
rect 317230 96636 317236 96648
rect 317288 96636 317294 96688
rect 329558 96676 329564 96688
rect 329519 96648 329564 96676
rect 329558 96636 329564 96648
rect 329616 96636 329622 96688
rect 354398 96676 354404 96688
rect 354359 96648 354404 96676
rect 354398 96636 354404 96648
rect 354456 96636 354462 96688
rect 232038 96568 232044 96620
rect 232096 96608 232102 96620
rect 232222 96608 232228 96620
rect 232096 96580 232228 96608
rect 232096 96568 232102 96580
rect 232222 96568 232228 96580
rect 232280 96568 232286 96620
rect 235166 96568 235172 96620
rect 235224 96608 235230 96620
rect 235350 96608 235356 96620
rect 235224 96580 235356 96608
rect 235224 96568 235230 96580
rect 235350 96568 235356 96580
rect 235408 96568 235414 96620
rect 217226 95384 217232 95396
rect 217187 95356 217232 95384
rect 217226 95344 217232 95356
rect 217284 95344 217290 95396
rect 191006 95208 191012 95260
rect 191064 95248 191070 95260
rect 191190 95248 191196 95260
rect 191064 95220 191196 95248
rect 191064 95208 191070 95220
rect 191190 95208 191196 95220
rect 191248 95208 191254 95260
rect 192386 95208 192392 95260
rect 192444 95208 192450 95260
rect 224037 95251 224095 95257
rect 224037 95217 224049 95251
rect 224083 95248 224095 95251
rect 224126 95248 224132 95260
rect 224083 95220 224132 95248
rect 224083 95217 224095 95220
rect 224037 95211 224095 95217
rect 224126 95208 224132 95220
rect 224184 95208 224190 95260
rect 225322 95248 225328 95260
rect 225283 95220 225328 95248
rect 225322 95208 225328 95220
rect 225380 95208 225386 95260
rect 261110 95248 261116 95260
rect 261071 95220 261116 95248
rect 261110 95208 261116 95220
rect 261168 95208 261174 95260
rect 275830 95248 275836 95260
rect 275791 95220 275836 95248
rect 275830 95208 275836 95220
rect 275888 95208 275894 95260
rect 277118 95248 277124 95260
rect 277079 95220 277124 95248
rect 277118 95208 277124 95220
rect 277176 95208 277182 95260
rect 282730 95248 282736 95260
rect 282691 95220 282736 95248
rect 282730 95208 282736 95220
rect 282788 95208 282794 95260
rect 283926 95248 283932 95260
rect 283887 95220 283932 95248
rect 283926 95208 283932 95220
rect 283984 95208 283990 95260
rect 192404 95124 192432 95208
rect 194873 95183 194931 95189
rect 194873 95149 194885 95183
rect 194919 95180 194931 95183
rect 194962 95180 194968 95192
rect 194919 95152 194968 95180
rect 194919 95149 194931 95152
rect 194873 95143 194931 95149
rect 194962 95140 194968 95152
rect 195020 95140 195026 95192
rect 178034 95072 178040 95124
rect 178092 95112 178098 95124
rect 178092 95084 178137 95112
rect 178092 95072 178098 95084
rect 192386 95072 192392 95124
rect 192444 95072 192450 95124
rect 230750 94528 230756 94580
rect 230808 94568 230814 94580
rect 230934 94568 230940 94580
rect 230808 94540 230940 94568
rect 230808 94528 230814 94540
rect 230934 94528 230940 94540
rect 230992 94528 230998 94580
rect 270126 94528 270132 94580
rect 270184 94568 270190 94580
rect 270310 94568 270316 94580
rect 270184 94540 270316 94568
rect 270184 94528 270190 94540
rect 270310 94528 270316 94540
rect 270368 94528 270374 94580
rect 219710 93888 219716 93900
rect 219671 93860 219716 93888
rect 219710 93848 219716 93860
rect 219768 93848 219774 93900
rect 343082 93848 343088 93900
rect 343140 93888 343146 93900
rect 343174 93888 343180 93900
rect 343140 93860 343180 93888
rect 343140 93848 343146 93860
rect 343174 93848 343180 93860
rect 343232 93848 343238 93900
rect 344462 93888 344468 93900
rect 344423 93860 344468 93888
rect 344462 93848 344468 93860
rect 344520 93848 344526 93900
rect 182177 93823 182235 93829
rect 182177 93789 182189 93823
rect 182223 93820 182235 93823
rect 182266 93820 182272 93832
rect 182223 93792 182272 93820
rect 182223 93789 182235 93792
rect 182177 93783 182235 93789
rect 182266 93780 182272 93792
rect 182324 93780 182330 93832
rect 355686 93820 355692 93832
rect 355647 93792 355692 93820
rect 355686 93780 355692 93792
rect 355744 93780 355750 93832
rect 361206 93820 361212 93832
rect 361167 93792 361212 93820
rect 361206 93780 361212 93792
rect 361264 93780 361270 93832
rect 177025 92531 177083 92537
rect 177025 92497 177037 92531
rect 177071 92528 177083 92531
rect 177114 92528 177120 92540
rect 177071 92500 177120 92528
rect 177071 92497 177083 92500
rect 177025 92491 177083 92497
rect 177114 92488 177120 92500
rect 177172 92488 177178 92540
rect 179966 92528 179972 92540
rect 179927 92500 179972 92528
rect 179966 92488 179972 92500
rect 180024 92488 180030 92540
rect 178037 91103 178095 91109
rect 178037 91069 178049 91103
rect 178083 91100 178095 91103
rect 178126 91100 178132 91112
rect 178083 91072 178132 91100
rect 178083 91069 178095 91072
rect 178037 91063 178095 91069
rect 178126 91060 178132 91072
rect 178184 91060 178190 91112
rect 192110 90380 192116 90432
rect 192168 90420 192174 90432
rect 192386 90420 192392 90432
rect 192168 90392 192392 90420
rect 192168 90380 192174 90392
rect 192386 90380 192392 90392
rect 192444 90380 192450 90432
rect 236362 89768 236368 89820
rect 236420 89768 236426 89820
rect 236380 89684 236408 89768
rect 258166 89700 258172 89752
rect 258224 89740 258230 89752
rect 258350 89740 258356 89752
rect 258224 89712 258356 89740
rect 258224 89700 258230 89712
rect 258350 89700 258356 89712
rect 258408 89700 258414 89752
rect 236362 89632 236368 89684
rect 236420 89632 236426 89684
rect 191190 87020 191196 87032
rect 191116 86992 191196 87020
rect 191116 86964 191144 86992
rect 191190 86980 191196 86992
rect 191248 86980 191254 87032
rect 315758 87020 315764 87032
rect 315719 86992 315764 87020
rect 315758 86980 315764 86992
rect 315816 86980 315822 87032
rect 171410 86952 171416 86964
rect 171371 86924 171416 86952
rect 171410 86912 171416 86924
rect 171468 86912 171474 86964
rect 173066 86952 173072 86964
rect 173027 86924 173072 86952
rect 173066 86912 173072 86924
rect 173124 86912 173130 86964
rect 191098 86912 191104 86964
rect 191156 86912 191162 86964
rect 201862 86952 201868 86964
rect 201823 86924 201868 86952
rect 201862 86912 201868 86924
rect 201920 86912 201926 86964
rect 211890 86912 211896 86964
rect 211948 86952 211954 86964
rect 211982 86952 211988 86964
rect 211948 86924 211988 86952
rect 211948 86912 211954 86924
rect 211982 86912 211988 86924
rect 212040 86912 212046 86964
rect 225230 86912 225236 86964
rect 225288 86952 225294 86964
rect 225322 86952 225328 86964
rect 225288 86924 225328 86952
rect 225288 86912 225294 86924
rect 225322 86912 225328 86924
rect 225380 86912 225386 86964
rect 228174 86912 228180 86964
rect 228232 86952 228238 86964
rect 228266 86952 228272 86964
rect 228232 86924 228272 86952
rect 228232 86912 228238 86924
rect 228266 86912 228272 86924
rect 228324 86912 228330 86964
rect 229278 86912 229284 86964
rect 229336 86912 229342 86964
rect 235074 86912 235080 86964
rect 235132 86912 235138 86964
rect 236270 86952 236276 86964
rect 236231 86924 236276 86952
rect 236270 86912 236276 86924
rect 236328 86912 236334 86964
rect 258258 86952 258264 86964
rect 258219 86924 258264 86952
rect 258258 86912 258264 86924
rect 258316 86912 258322 86964
rect 262309 86955 262367 86961
rect 262309 86921 262321 86955
rect 262355 86952 262367 86955
rect 262398 86952 262404 86964
rect 262355 86924 262404 86952
rect 262355 86921 262367 86924
rect 262309 86915 262367 86921
rect 262398 86912 262404 86924
rect 262456 86912 262462 86964
rect 229296 86884 229324 86912
rect 229370 86884 229376 86896
rect 229296 86856 229376 86884
rect 229370 86844 229376 86856
rect 229428 86844 229434 86896
rect 235092 86884 235120 86912
rect 235166 86884 235172 86896
rect 235092 86856 235172 86884
rect 235166 86844 235172 86856
rect 235224 86844 235230 86896
rect 270126 86096 270132 86148
rect 270184 86136 270190 86148
rect 270310 86136 270316 86148
rect 270184 86108 270316 86136
rect 270184 86096 270190 86108
rect 270310 86096 270316 86108
rect 270368 86096 270374 86148
rect 200390 85660 200396 85672
rect 200316 85632 200396 85660
rect 200316 85604 200344 85632
rect 200390 85620 200396 85632
rect 200448 85620 200454 85672
rect 177022 85552 177028 85604
rect 177080 85592 177086 85604
rect 177114 85592 177120 85604
rect 177080 85564 177120 85592
rect 177080 85552 177086 85564
rect 177114 85552 177120 85564
rect 177172 85552 177178 85604
rect 194870 85592 194876 85604
rect 194831 85564 194876 85592
rect 194870 85552 194876 85564
rect 194928 85552 194934 85604
rect 200298 85552 200304 85604
rect 200356 85552 200362 85604
rect 224034 85552 224040 85604
rect 224092 85592 224098 85604
rect 224126 85592 224132 85604
rect 224092 85564 224132 85592
rect 224092 85552 224098 85564
rect 224126 85552 224132 85564
rect 224184 85552 224190 85604
rect 362310 85552 362316 85604
rect 362368 85592 362374 85604
rect 362494 85592 362500 85604
rect 362368 85564 362500 85592
rect 362368 85552 362374 85564
rect 362494 85552 362500 85564
rect 362552 85552 362558 85604
rect 212258 85484 212264 85536
rect 212316 85524 212322 85536
rect 212442 85524 212448 85536
rect 212316 85496 212448 85524
rect 212316 85484 212322 85496
rect 212442 85484 212448 85496
rect 212500 85484 212506 85536
rect 228174 85484 228180 85536
rect 228232 85524 228238 85536
rect 228266 85524 228272 85536
rect 228232 85496 228272 85524
rect 228232 85484 228238 85496
rect 228266 85484 228272 85496
rect 228324 85484 228330 85536
rect 260929 85527 260987 85533
rect 260929 85493 260941 85527
rect 260975 85524 260987 85527
rect 261110 85524 261116 85536
rect 260975 85496 261116 85524
rect 260975 85493 260987 85496
rect 260929 85487 260987 85493
rect 261110 85484 261116 85496
rect 261168 85484 261174 85536
rect 283926 85524 283932 85536
rect 283887 85496 283932 85524
rect 283926 85484 283932 85496
rect 283984 85484 283990 85536
rect 289265 85527 289323 85533
rect 289265 85493 289277 85527
rect 289311 85524 289323 85527
rect 289354 85524 289360 85536
rect 289311 85496 289360 85524
rect 289311 85493 289323 85496
rect 289265 85487 289323 85493
rect 289354 85484 289360 85496
rect 289412 85484 289418 85536
rect 361206 85524 361212 85536
rect 361167 85496 361212 85524
rect 361206 85484 361212 85496
rect 361264 85484 361270 85536
rect 230750 84872 230756 84924
rect 230808 84912 230814 84924
rect 230934 84912 230940 84924
rect 230808 84884 230940 84912
rect 230808 84872 230814 84884
rect 230934 84872 230940 84884
rect 230992 84872 230998 84924
rect 341978 84328 341984 84380
rect 342036 84328 342042 84380
rect 341996 84244 342024 84328
rect 182174 84232 182180 84244
rect 182135 84204 182180 84232
rect 182174 84192 182180 84204
rect 182232 84192 182238 84244
rect 217226 84232 217232 84244
rect 217187 84204 217232 84232
rect 217226 84192 217232 84204
rect 217284 84192 217290 84244
rect 219526 84192 219532 84244
rect 219584 84232 219590 84244
rect 219802 84232 219808 84244
rect 219584 84204 219808 84232
rect 219584 84192 219590 84204
rect 219802 84192 219808 84204
rect 219860 84192 219866 84244
rect 341978 84192 341984 84244
rect 342036 84192 342042 84244
rect 355686 84232 355692 84244
rect 355647 84204 355692 84232
rect 355686 84192 355692 84204
rect 355744 84192 355750 84244
rect 191098 84164 191104 84176
rect 191059 84136 191104 84164
rect 191098 84124 191104 84136
rect 191156 84124 191162 84176
rect 192202 84124 192208 84176
rect 192260 84164 192266 84176
rect 192297 84167 192355 84173
rect 192297 84164 192309 84167
rect 192260 84136 192309 84164
rect 192260 84124 192266 84136
rect 192297 84133 192309 84136
rect 192343 84133 192355 84167
rect 192297 84127 192355 84133
rect 275738 84124 275744 84176
rect 275796 84164 275802 84176
rect 275922 84164 275928 84176
rect 275796 84136 275928 84164
rect 275796 84124 275802 84136
rect 275922 84124 275928 84136
rect 275980 84124 275986 84176
rect 343266 84164 343272 84176
rect 343227 84136 343272 84164
rect 343266 84124 343272 84136
rect 343324 84124 343330 84176
rect 345566 84164 345572 84176
rect 345527 84136 345572 84164
rect 345566 84124 345572 84136
rect 345624 84124 345630 84176
rect 361298 84164 361304 84176
rect 361259 84136 361304 84164
rect 361298 84124 361304 84136
rect 361356 84124 361362 84176
rect 362313 84167 362371 84173
rect 362313 84133 362325 84167
rect 362359 84164 362371 84167
rect 362494 84164 362500 84176
rect 362359 84136 362500 84164
rect 362359 84133 362371 84136
rect 362313 84127 362371 84133
rect 362494 84124 362500 84136
rect 362552 84124 362558 84176
rect 179966 82804 179972 82816
rect 179927 82776 179972 82804
rect 179966 82764 179972 82776
rect 180024 82764 180030 82816
rect 178126 81376 178132 81388
rect 178087 81348 178132 81376
rect 178126 81336 178132 81348
rect 178184 81336 178190 81388
rect 203058 80696 203064 80708
rect 203019 80668 203064 80696
rect 203058 80656 203064 80668
rect 203116 80656 203122 80708
rect 235258 80084 235264 80096
rect 235219 80056 235264 80084
rect 235258 80044 235264 80056
rect 235316 80044 235322 80096
rect 291930 80084 291936 80096
rect 291856 80056 291936 80084
rect 291856 80028 291884 80056
rect 291930 80044 291936 80056
rect 291988 80044 291994 80096
rect 291838 79976 291844 80028
rect 291896 79976 291902 80028
rect 344554 79336 344560 79348
rect 344515 79308 344560 79336
rect 344554 79296 344560 79308
rect 344612 79296 344618 79348
rect 361301 79339 361359 79345
rect 361301 79305 361313 79339
rect 361347 79336 361359 79339
rect 361390 79336 361396 79348
rect 361347 79308 361396 79336
rect 361347 79305 361359 79308
rect 361301 79299 361359 79305
rect 361390 79296 361396 79308
rect 361448 79296 361454 79348
rect 318245 77571 318303 77577
rect 318245 77537 318257 77571
rect 318291 77568 318303 77571
rect 318518 77568 318524 77580
rect 318291 77540 318524 77568
rect 318291 77537 318303 77540
rect 318245 77531 318303 77537
rect 318518 77528 318524 77540
rect 318576 77528 318582 77580
rect 229370 77460 229376 77512
rect 229428 77460 229434 77512
rect 229388 77376 229416 77460
rect 224034 77364 224040 77376
rect 223960 77336 224040 77364
rect 171410 77296 171416 77308
rect 171371 77268 171416 77296
rect 171410 77256 171416 77268
rect 171468 77256 171474 77308
rect 173066 77296 173072 77308
rect 173027 77268 173072 77296
rect 173066 77256 173072 77268
rect 173124 77256 173130 77308
rect 200298 77256 200304 77308
rect 200356 77296 200362 77308
rect 200390 77296 200396 77308
rect 200356 77268 200396 77296
rect 200356 77256 200362 77268
rect 200390 77256 200396 77268
rect 200448 77256 200454 77308
rect 201862 77296 201868 77308
rect 201823 77268 201868 77296
rect 201862 77256 201868 77268
rect 201920 77256 201926 77308
rect 223960 77240 223988 77336
rect 224034 77324 224040 77336
rect 224092 77324 224098 77376
rect 229370 77324 229376 77376
rect 229428 77324 229434 77376
rect 282733 77367 282791 77373
rect 282733 77333 282745 77367
rect 282779 77364 282791 77367
rect 282822 77364 282828 77376
rect 282779 77336 282828 77364
rect 282779 77333 282791 77336
rect 282733 77327 282791 77333
rect 282822 77324 282828 77336
rect 282880 77324 282886 77376
rect 232222 77296 232228 77308
rect 232183 77268 232228 77296
rect 232222 77256 232228 77268
rect 232280 77256 232286 77308
rect 235258 77296 235264 77308
rect 235219 77268 235264 77296
rect 235258 77256 235264 77268
rect 235316 77256 235322 77308
rect 258261 77299 258319 77305
rect 258261 77265 258273 77299
rect 258307 77296 258319 77299
rect 258350 77296 258356 77308
rect 258307 77268 258356 77296
rect 258307 77265 258319 77268
rect 258261 77259 258319 77265
rect 258350 77256 258356 77268
rect 258408 77256 258414 77308
rect 262306 77296 262312 77308
rect 262267 77268 262312 77296
rect 262306 77256 262312 77268
rect 262364 77256 262370 77308
rect 182358 77188 182364 77240
rect 182416 77188 182422 77240
rect 194870 77228 194876 77240
rect 194831 77200 194876 77228
rect 194870 77188 194876 77200
rect 194928 77188 194934 77240
rect 223942 77188 223948 77240
rect 224000 77188 224006 77240
rect 182376 77104 182404 77188
rect 182358 77052 182364 77104
rect 182416 77052 182422 77104
rect 189350 75896 189356 75948
rect 189408 75936 189414 75948
rect 189442 75936 189448 75948
rect 189408 75908 189448 75936
rect 189408 75896 189414 75908
rect 189442 75896 189448 75908
rect 189500 75896 189506 75948
rect 217134 75896 217140 75948
rect 217192 75936 217198 75948
rect 217318 75936 217324 75948
rect 217192 75908 217324 75936
rect 217192 75896 217198 75908
rect 217318 75896 217324 75908
rect 217376 75896 217382 75948
rect 232222 75936 232228 75948
rect 232183 75908 232228 75936
rect 232222 75896 232228 75908
rect 232280 75896 232286 75948
rect 236273 75939 236331 75945
rect 236273 75905 236285 75939
rect 236319 75936 236331 75939
rect 236454 75936 236460 75948
rect 236319 75908 236460 75936
rect 236319 75905 236331 75908
rect 236273 75899 236331 75905
rect 236454 75896 236460 75908
rect 236512 75896 236518 75948
rect 260926 75936 260932 75948
rect 260887 75908 260932 75936
rect 260926 75896 260932 75908
rect 260984 75896 260990 75948
rect 282730 75936 282736 75948
rect 282691 75908 282736 75936
rect 282730 75896 282736 75908
rect 282788 75896 282794 75948
rect 283929 75939 283987 75945
rect 283929 75905 283941 75939
rect 283975 75936 283987 75939
rect 284018 75936 284024 75948
rect 283975 75908 284024 75936
rect 283975 75905 283987 75908
rect 283929 75899 283987 75905
rect 284018 75896 284024 75908
rect 284076 75896 284082 75948
rect 289262 75936 289268 75948
rect 289223 75908 289268 75936
rect 289262 75896 289268 75908
rect 289320 75896 289326 75948
rect 318242 75936 318248 75948
rect 318203 75908 318248 75936
rect 318242 75896 318248 75908
rect 318300 75896 318306 75948
rect 184014 75868 184020 75880
rect 183975 75840 184020 75868
rect 184014 75828 184020 75840
rect 184072 75828 184078 75880
rect 355962 75868 355968 75880
rect 355923 75840 355968 75868
rect 355962 75828 355968 75840
rect 356020 75828 356026 75880
rect 217134 75800 217140 75812
rect 217095 75772 217140 75800
rect 217134 75760 217140 75772
rect 217192 75760 217198 75812
rect 355870 75760 355876 75812
rect 355928 75760 355934 75812
rect 355778 75692 355784 75744
rect 355836 75692 355842 75744
rect 355796 75608 355824 75692
rect 355888 75676 355916 75760
rect 355870 75624 355876 75676
rect 355928 75624 355934 75676
rect 355778 75556 355784 75608
rect 355836 75556 355842 75608
rect 230750 75216 230756 75268
rect 230808 75256 230814 75268
rect 230934 75256 230940 75268
rect 230808 75228 230940 75256
rect 230808 75216 230814 75228
rect 230934 75216 230940 75228
rect 230992 75216 230998 75268
rect 270126 75216 270132 75268
rect 270184 75256 270190 75268
rect 270310 75256 270316 75268
rect 270184 75228 270316 75256
rect 270184 75216 270190 75228
rect 270310 75216 270316 75228
rect 270368 75216 270374 75268
rect 277118 74604 277124 74656
rect 277176 74644 277182 74656
rect 277210 74644 277216 74656
rect 277176 74616 277216 74644
rect 277176 74604 277182 74616
rect 277210 74604 277216 74616
rect 277268 74604 277274 74656
rect 341978 74644 341984 74656
rect 341939 74616 341984 74644
rect 341978 74604 341984 74616
rect 342036 74604 342042 74656
rect 191101 74579 191159 74585
rect 191101 74545 191113 74579
rect 191147 74576 191159 74579
rect 191282 74576 191288 74588
rect 191147 74548 191288 74576
rect 191147 74545 191159 74548
rect 191101 74539 191159 74545
rect 191282 74536 191288 74548
rect 191340 74536 191346 74588
rect 343269 74579 343327 74585
rect 343269 74545 343281 74579
rect 343315 74576 343327 74579
rect 343358 74576 343364 74588
rect 343315 74548 343364 74576
rect 343315 74545 343327 74548
rect 343269 74539 343327 74545
rect 343358 74536 343364 74548
rect 343416 74536 343422 74588
rect 345569 74579 345627 74585
rect 345569 74545 345581 74579
rect 345615 74576 345627 74579
rect 345658 74576 345664 74588
rect 345615 74548 345664 74576
rect 345615 74545 345627 74548
rect 345569 74539 345627 74545
rect 345658 74536 345664 74548
rect 345716 74536 345722 74588
rect 181254 74508 181260 74520
rect 181215 74480 181260 74508
rect 181254 74468 181260 74480
rect 181312 74468 181318 74520
rect 341978 73284 341984 73296
rect 341939 73256 341984 73284
rect 341978 73244 341984 73256
rect 342036 73244 342042 73296
rect 179966 73216 179972 73228
rect 179927 73188 179972 73216
rect 179966 73176 179972 73188
rect 180024 73176 180030 73228
rect 203058 71108 203064 71120
rect 203019 71080 203064 71108
rect 203058 71068 203064 71080
rect 203116 71068 203122 71120
rect 211890 70456 211896 70508
rect 211948 70456 211954 70508
rect 219713 70499 219771 70505
rect 219713 70465 219725 70499
rect 219759 70496 219771 70499
rect 219802 70496 219808 70508
rect 219759 70468 219808 70496
rect 219759 70465 219771 70468
rect 219713 70459 219771 70465
rect 219802 70456 219808 70468
rect 219860 70456 219866 70508
rect 211908 70372 211936 70456
rect 258166 70388 258172 70440
rect 258224 70428 258230 70440
rect 258224 70400 258304 70428
rect 258224 70388 258230 70400
rect 258276 70372 258304 70400
rect 211890 70320 211896 70372
rect 211948 70320 211954 70372
rect 258258 70320 258264 70372
rect 258316 70320 258322 70372
rect 329558 67736 329564 67788
rect 329616 67736 329622 67788
rect 235166 67708 235172 67720
rect 235092 67680 235172 67708
rect 235092 67652 235120 67680
rect 235166 67668 235172 67680
rect 235224 67668 235230 67720
rect 329576 67652 329604 67736
rect 225230 67600 225236 67652
rect 225288 67640 225294 67652
rect 225322 67640 225328 67652
rect 225288 67612 225328 67640
rect 225288 67600 225294 67612
rect 225322 67600 225328 67612
rect 225380 67600 225386 67652
rect 232038 67600 232044 67652
rect 232096 67640 232102 67652
rect 232222 67640 232228 67652
rect 232096 67612 232228 67640
rect 232096 67600 232102 67612
rect 232222 67600 232228 67612
rect 232280 67600 232286 67652
rect 235074 67600 235080 67652
rect 235132 67600 235138 67652
rect 236270 67600 236276 67652
rect 236328 67640 236334 67652
rect 236454 67640 236460 67652
rect 236328 67612 236460 67640
rect 236328 67600 236334 67612
rect 236454 67600 236460 67612
rect 236512 67600 236518 67652
rect 282730 67600 282736 67652
rect 282788 67640 282794 67652
rect 282822 67640 282828 67652
rect 282788 67612 282828 67640
rect 282788 67600 282794 67612
rect 282822 67600 282828 67612
rect 282880 67600 282886 67652
rect 285214 67600 285220 67652
rect 285272 67640 285278 67652
rect 285306 67640 285312 67652
rect 285272 67612 285312 67640
rect 285272 67600 285278 67612
rect 285306 67600 285312 67612
rect 285364 67600 285370 67652
rect 286502 67600 286508 67652
rect 286560 67640 286566 67652
rect 286594 67640 286600 67652
rect 286560 67612 286600 67640
rect 286560 67600 286566 67612
rect 286594 67600 286600 67612
rect 286652 67600 286658 67652
rect 289262 67600 289268 67652
rect 289320 67640 289326 67652
rect 289354 67640 289360 67652
rect 289320 67612 289360 67640
rect 289320 67600 289326 67612
rect 289354 67600 289360 67612
rect 289412 67600 289418 67652
rect 317046 67600 317052 67652
rect 317104 67640 317110 67652
rect 317230 67640 317236 67652
rect 317104 67612 317236 67640
rect 317104 67600 317110 67612
rect 317230 67600 317236 67612
rect 317288 67600 317294 67652
rect 329558 67600 329564 67652
rect 329616 67600 329622 67652
rect 344554 67640 344560 67652
rect 344515 67612 344560 67640
rect 344554 67600 344560 67612
rect 344612 67600 344618 67652
rect 362310 67640 362316 67652
rect 362271 67612 362316 67640
rect 362310 67600 362316 67612
rect 362368 67600 362374 67652
rect 171410 67572 171416 67584
rect 171371 67544 171416 67572
rect 171410 67532 171416 67544
rect 171468 67532 171474 67584
rect 173066 67572 173072 67584
rect 173027 67544 173072 67572
rect 173066 67532 173072 67544
rect 173124 67532 173130 67584
rect 223942 67532 223948 67584
rect 224000 67532 224006 67584
rect 229278 67532 229284 67584
rect 229336 67532 229342 67584
rect 223960 67504 223988 67532
rect 224034 67504 224040 67516
rect 223960 67476 224040 67504
rect 224034 67464 224040 67476
rect 224092 67464 224098 67516
rect 229296 67504 229324 67532
rect 229370 67504 229376 67516
rect 229296 67476 229376 67504
rect 229370 67464 229376 67476
rect 229428 67464 229434 67516
rect 362218 67464 362224 67516
rect 362276 67504 362282 67516
rect 362310 67504 362316 67516
rect 362276 67476 362316 67504
rect 362276 67464 362282 67476
rect 362310 67464 362316 67476
rect 362368 67464 362374 67516
rect 355962 67368 355968 67380
rect 355923 67340 355968 67368
rect 355962 67328 355968 67340
rect 356020 67328 356026 67380
rect 184017 66283 184075 66289
rect 184017 66249 184029 66283
rect 184063 66280 184075 66283
rect 184106 66280 184112 66292
rect 184063 66252 184112 66280
rect 184063 66249 184075 66252
rect 184017 66243 184075 66249
rect 184106 66240 184112 66252
rect 184164 66240 184170 66292
rect 192202 66240 192208 66292
rect 192260 66280 192266 66292
rect 192297 66283 192355 66289
rect 192297 66280 192309 66283
rect 192260 66252 192309 66280
rect 192260 66240 192266 66252
rect 192297 66249 192309 66252
rect 192343 66249 192355 66283
rect 192297 66243 192355 66249
rect 194873 66283 194931 66289
rect 194873 66249 194885 66283
rect 194919 66280 194931 66283
rect 194962 66280 194968 66292
rect 194919 66252 194968 66280
rect 194919 66249 194931 66252
rect 194873 66243 194931 66249
rect 194962 66240 194968 66252
rect 195020 66240 195026 66292
rect 217137 66283 217195 66289
rect 217137 66249 217149 66283
rect 217183 66280 217195 66283
rect 217226 66280 217232 66292
rect 217183 66252 217232 66280
rect 217183 66249 217195 66252
rect 217137 66243 217195 66249
rect 217226 66240 217232 66252
rect 217284 66240 217290 66292
rect 219710 66280 219716 66292
rect 219671 66252 219716 66280
rect 219710 66240 219716 66252
rect 219768 66240 219774 66292
rect 203058 66172 203064 66224
rect 203116 66212 203122 66224
rect 203334 66212 203340 66224
rect 203116 66184 203340 66212
rect 203116 66172 203122 66184
rect 203334 66172 203340 66184
rect 203392 66172 203398 66224
rect 212258 66172 212264 66224
rect 212316 66212 212322 66224
rect 212350 66212 212356 66224
rect 212316 66184 212356 66212
rect 212316 66172 212322 66184
rect 212350 66172 212356 66184
rect 212408 66172 212414 66224
rect 235074 66172 235080 66224
rect 235132 66172 235138 66224
rect 275830 66172 275836 66224
rect 275888 66172 275894 66224
rect 283929 66215 283987 66221
rect 283929 66181 283941 66215
rect 283975 66212 283987 66215
rect 284018 66212 284024 66224
rect 283975 66184 284024 66212
rect 283975 66181 283987 66184
rect 283929 66175 283987 66181
rect 284018 66172 284024 66184
rect 284076 66172 284082 66224
rect 285306 66212 285312 66224
rect 285267 66184 285312 66212
rect 285306 66172 285312 66184
rect 285364 66172 285370 66224
rect 286594 66212 286600 66224
rect 286555 66184 286600 66212
rect 286594 66172 286600 66184
rect 286652 66172 286658 66224
rect 289354 66212 289360 66224
rect 289315 66184 289360 66212
rect 289354 66172 289360 66184
rect 289412 66172 289418 66224
rect 291930 66172 291936 66224
rect 291988 66212 291994 66224
rect 329558 66212 329564 66224
rect 291988 66184 292068 66212
rect 329519 66184 329564 66212
rect 291988 66172 291994 66184
rect 235092 66144 235120 66172
rect 235166 66144 235172 66156
rect 235092 66116 235172 66144
rect 235166 66104 235172 66116
rect 235224 66104 235230 66156
rect 275848 66144 275876 66172
rect 292040 66156 292068 66184
rect 329558 66172 329564 66184
rect 329616 66172 329622 66224
rect 276014 66144 276020 66156
rect 275848 66116 276020 66144
rect 276014 66104 276020 66116
rect 276072 66104 276078 66156
rect 292022 66104 292028 66156
rect 292080 66104 292086 66156
rect 230750 65940 230756 65952
rect 230711 65912 230756 65940
rect 230750 65900 230756 65912
rect 230808 65900 230814 65952
rect 234982 65492 234988 65544
rect 235040 65532 235046 65544
rect 235258 65532 235264 65544
rect 235040 65504 235264 65532
rect 235040 65492 235046 65504
rect 235258 65492 235264 65504
rect 235316 65492 235322 65544
rect 270126 65492 270132 65544
rect 270184 65532 270190 65544
rect 270310 65532 270316 65544
rect 270184 65504 270316 65532
rect 270184 65492 270190 65504
rect 270310 65492 270316 65504
rect 270368 65492 270374 65544
rect 181070 64880 181076 64932
rect 181128 64920 181134 64932
rect 181257 64923 181315 64929
rect 181257 64920 181269 64923
rect 181128 64892 181269 64920
rect 181128 64880 181134 64892
rect 181257 64889 181269 64892
rect 181303 64889 181315 64923
rect 181257 64883 181315 64889
rect 341886 64880 341892 64932
rect 341944 64880 341950 64932
rect 203061 64855 203119 64861
rect 203061 64821 203073 64855
rect 203107 64852 203119 64855
rect 203334 64852 203340 64864
rect 203107 64824 203340 64852
rect 203107 64821 203119 64824
rect 203061 64815 203119 64821
rect 203334 64812 203340 64824
rect 203392 64812 203398 64864
rect 341904 64784 341932 64880
rect 344465 64855 344523 64861
rect 344465 64821 344477 64855
rect 344511 64852 344523 64855
rect 344554 64852 344560 64864
rect 344511 64824 344560 64852
rect 344511 64821 344523 64824
rect 344465 64815 344523 64821
rect 344554 64812 344560 64824
rect 344612 64812 344618 64864
rect 355597 64855 355655 64861
rect 355597 64821 355609 64855
rect 355643 64852 355655 64855
rect 355686 64852 355692 64864
rect 355643 64824 355692 64852
rect 355643 64821 355655 64824
rect 355597 64815 355655 64821
rect 355686 64812 355692 64824
rect 355744 64812 355750 64864
rect 341978 64784 341984 64796
rect 341904 64756 341984 64784
rect 341978 64744 341984 64756
rect 342036 64744 342042 64796
rect 178129 63563 178187 63569
rect 178129 63529 178141 63563
rect 178175 63560 178187 63563
rect 178310 63560 178316 63572
rect 178175 63532 178316 63560
rect 178175 63529 178187 63532
rect 178129 63523 178187 63529
rect 178310 63520 178316 63532
rect 178368 63520 178374 63572
rect 177022 63492 177028 63504
rect 176983 63464 177028 63492
rect 177022 63452 177028 63464
rect 177080 63452 177086 63504
rect 179966 63492 179972 63504
rect 179927 63464 179972 63492
rect 179966 63452 179972 63464
rect 180024 63452 180030 63504
rect 275741 63495 275799 63501
rect 275741 63461 275753 63495
rect 275787 63492 275799 63495
rect 275922 63492 275928 63504
rect 275787 63464 275928 63492
rect 275787 63461 275799 63464
rect 275741 63455 275799 63461
rect 275922 63452 275928 63464
rect 275980 63452 275986 63504
rect 277121 63495 277179 63501
rect 277121 63461 277133 63495
rect 277167 63492 277179 63495
rect 277210 63492 277216 63504
rect 277167 63464 277216 63492
rect 277167 63461 277179 63464
rect 277121 63455 277179 63461
rect 277210 63452 277216 63464
rect 277268 63452 277274 63504
rect 341978 63492 341984 63504
rect 341904 63464 341984 63492
rect 341904 63436 341932 63464
rect 341978 63452 341984 63464
rect 342036 63452 342042 63504
rect 343174 63452 343180 63504
rect 343232 63492 343238 63504
rect 343358 63492 343364 63504
rect 343232 63464 343364 63492
rect 343232 63452 343238 63464
rect 343358 63452 343364 63464
rect 343416 63452 343422 63504
rect 341886 63384 341892 63436
rect 341944 63384 341950 63436
rect 200390 61452 200396 61464
rect 200351 61424 200396 61452
rect 200390 61412 200396 61424
rect 200448 61412 200454 61464
rect 201862 61452 201868 61464
rect 201823 61424 201868 61452
rect 201862 61412 201868 61424
rect 201920 61412 201926 61464
rect 262398 60664 262404 60716
rect 262456 60704 262462 60716
rect 262582 60704 262588 60716
rect 262456 60676 262588 60704
rect 262456 60664 262462 60676
rect 262582 60664 262588 60676
rect 262640 60664 262646 60716
rect 234982 60596 234988 60648
rect 235040 60636 235046 60648
rect 235258 60636 235264 60648
rect 235040 60608 235264 60636
rect 235040 60596 235046 60608
rect 235258 60596 235264 60608
rect 235316 60596 235322 60648
rect 345566 59984 345572 60036
rect 345624 60024 345630 60036
rect 345661 60027 345719 60033
rect 345661 60024 345673 60027
rect 345624 59996 345673 60024
rect 345624 59984 345630 59996
rect 345661 59993 345673 59996
rect 345707 59993 345719 60027
rect 345661 59987 345719 59993
rect 181070 58664 181076 58676
rect 181031 58636 181076 58664
rect 181070 58624 181076 58636
rect 181128 58624 181134 58676
rect 354398 58148 354404 58200
rect 354456 58148 354462 58200
rect 354416 58064 354444 58148
rect 354398 58012 354404 58064
rect 354456 58012 354462 58064
rect 171410 57984 171416 57996
rect 171371 57956 171416 57984
rect 171410 57944 171416 57956
rect 171468 57944 171474 57996
rect 173066 57984 173072 57996
rect 173027 57956 173072 57984
rect 173066 57944 173072 57956
rect 173124 57944 173130 57996
rect 315758 57944 315764 57996
rect 315816 57984 315822 57996
rect 315850 57984 315856 57996
rect 315816 57956 315856 57984
rect 315816 57944 315822 57956
rect 315850 57944 315856 57956
rect 315908 57944 315914 57996
rect 328178 57944 328184 57996
rect 328236 57984 328242 57996
rect 328270 57984 328276 57996
rect 328236 57956 328276 57984
rect 328236 57944 328242 57956
rect 328270 57944 328276 57956
rect 328328 57944 328334 57996
rect 177025 57919 177083 57925
rect 177025 57885 177037 57919
rect 177071 57916 177083 57919
rect 177114 57916 177120 57928
rect 177071 57888 177120 57916
rect 177071 57885 177083 57888
rect 177025 57879 177083 57885
rect 177114 57876 177120 57888
rect 177172 57876 177178 57928
rect 183922 57876 183928 57928
rect 183980 57916 183986 57928
rect 184106 57916 184112 57928
rect 183980 57888 184112 57916
rect 183980 57876 183986 57888
rect 184106 57876 184112 57888
rect 184164 57876 184170 57928
rect 261018 57876 261024 57928
rect 261076 57916 261082 57928
rect 261110 57916 261116 57928
rect 261076 57888 261116 57916
rect 261076 57876 261082 57888
rect 261110 57876 261116 57888
rect 261168 57876 261174 57928
rect 262493 57919 262551 57925
rect 262493 57885 262505 57919
rect 262539 57916 262551 57919
rect 262582 57916 262588 57928
rect 262539 57888 262588 57916
rect 262539 57885 262551 57888
rect 262493 57879 262551 57885
rect 262582 57876 262588 57888
rect 262640 57876 262646 57928
rect 318334 57876 318340 57928
rect 318392 57916 318398 57928
rect 318518 57916 318524 57928
rect 318392 57888 318524 57916
rect 318392 57876 318398 57888
rect 318518 57876 318524 57888
rect 318576 57876 318582 57928
rect 354309 57919 354367 57925
rect 354309 57885 354321 57919
rect 354355 57916 354367 57919
rect 354398 57916 354404 57928
rect 354355 57888 354404 57916
rect 354355 57885 354367 57888
rect 354309 57879 354367 57885
rect 354398 57876 354404 57888
rect 354456 57876 354462 57928
rect 362310 57916 362316 57928
rect 362271 57888 362316 57916
rect 362310 57876 362316 57888
rect 362368 57876 362374 57928
rect 283926 56692 283932 56704
rect 283887 56664 283932 56692
rect 283926 56652 283932 56664
rect 283984 56652 283990 56704
rect 219710 56584 219716 56636
rect 219768 56624 219774 56636
rect 219802 56624 219808 56636
rect 219768 56596 219808 56624
rect 219768 56584 219774 56596
rect 219802 56584 219808 56596
rect 219860 56584 219866 56636
rect 230753 56627 230811 56633
rect 230753 56593 230765 56627
rect 230799 56624 230811 56627
rect 231026 56624 231032 56636
rect 230799 56596 231032 56624
rect 230799 56593 230811 56596
rect 230753 56587 230811 56593
rect 231026 56584 231032 56596
rect 231084 56584 231090 56636
rect 285309 56627 285367 56633
rect 285309 56593 285321 56627
rect 285355 56624 285367 56627
rect 285398 56624 285404 56636
rect 285355 56596 285404 56624
rect 285355 56593 285367 56596
rect 285309 56587 285367 56593
rect 285398 56584 285404 56596
rect 285456 56584 285462 56636
rect 286597 56627 286655 56633
rect 286597 56593 286609 56627
rect 286643 56624 286655 56627
rect 286686 56624 286692 56636
rect 286643 56596 286692 56624
rect 286643 56593 286655 56596
rect 286597 56587 286655 56593
rect 286686 56584 286692 56596
rect 286744 56584 286750 56636
rect 289357 56627 289415 56633
rect 289357 56593 289369 56627
rect 289403 56624 289415 56627
rect 289446 56624 289452 56636
rect 289403 56596 289452 56624
rect 289403 56593 289415 56596
rect 289357 56587 289415 56593
rect 289446 56584 289452 56596
rect 289504 56584 289510 56636
rect 329558 56624 329564 56636
rect 329519 56596 329564 56624
rect 329558 56584 329564 56596
rect 329616 56584 329622 56636
rect 225230 56516 225236 56568
rect 225288 56556 225294 56568
rect 225506 56556 225512 56568
rect 225288 56528 225512 56556
rect 225288 56516 225294 56528
rect 225506 56516 225512 56528
rect 225564 56516 225570 56568
rect 261018 56516 261024 56568
rect 261076 56516 261082 56568
rect 283926 56556 283932 56568
rect 283887 56528 283932 56556
rect 283926 56516 283932 56528
rect 283984 56516 283990 56568
rect 318334 56556 318340 56568
rect 318295 56528 318340 56556
rect 318334 56516 318340 56528
rect 318392 56516 318398 56568
rect 231026 56448 231032 56500
rect 231084 56488 231090 56500
rect 231394 56488 231400 56500
rect 231084 56460 231400 56488
rect 231084 56448 231090 56460
rect 231394 56448 231400 56460
rect 231452 56448 231458 56500
rect 261036 56488 261064 56516
rect 261202 56488 261208 56500
rect 261036 56460 261208 56488
rect 261202 56448 261208 56460
rect 261260 56448 261266 56500
rect 203058 55264 203064 55276
rect 203019 55236 203064 55264
rect 203058 55224 203064 55236
rect 203116 55224 203122 55276
rect 344462 55264 344468 55276
rect 344423 55236 344468 55264
rect 344462 55224 344468 55236
rect 344520 55224 344526 55276
rect 183922 55196 183928 55208
rect 183883 55168 183928 55196
rect 183922 55156 183928 55168
rect 183980 55156 183986 55208
rect 228174 55196 228180 55208
rect 228135 55168 228180 55196
rect 228174 55156 228180 55168
rect 228232 55156 228238 55208
rect 270126 54612 270132 54664
rect 270184 54652 270190 54664
rect 270310 54652 270316 54664
rect 270184 54624 270316 54652
rect 270184 54612 270190 54624
rect 270310 54612 270316 54624
rect 270368 54612 270374 54664
rect 201865 53975 201923 53981
rect 201865 53941 201877 53975
rect 201911 53972 201923 53975
rect 202046 53972 202052 53984
rect 201911 53944 202052 53972
rect 201911 53941 201923 53944
rect 201865 53935 201923 53941
rect 202046 53932 202052 53944
rect 202104 53932 202110 53984
rect 178034 53796 178040 53848
rect 178092 53836 178098 53848
rect 178126 53836 178132 53848
rect 178092 53808 178132 53836
rect 178092 53796 178098 53808
rect 178126 53796 178132 53808
rect 178184 53796 178190 53848
rect 179966 53836 179972 53848
rect 179927 53808 179972 53836
rect 179966 53796 179972 53808
rect 180024 53796 180030 53848
rect 181073 53839 181131 53845
rect 181073 53805 181085 53839
rect 181119 53836 181131 53839
rect 181162 53836 181168 53848
rect 181119 53808 181168 53836
rect 181119 53805 181131 53808
rect 181073 53799 181131 53805
rect 181162 53796 181168 53808
rect 181220 53796 181226 53848
rect 275738 53836 275744 53848
rect 275699 53808 275744 53836
rect 275738 53796 275744 53808
rect 275796 53796 275802 53848
rect 275738 53116 275744 53168
rect 275796 53156 275802 53168
rect 275922 53156 275928 53168
rect 275796 53128 275928 53156
rect 275796 53116 275802 53128
rect 275922 53116 275928 53128
rect 275980 53116 275986 53168
rect 327902 53116 327908 53168
rect 327960 53156 327966 53168
rect 328270 53156 328276 53168
rect 327960 53128 328276 53156
rect 327960 53116 327966 53128
rect 328270 53116 328276 53128
rect 328328 53116 328334 53168
rect 344462 51756 344468 51808
rect 344520 51796 344526 51808
rect 344557 51799 344615 51805
rect 344557 51796 344569 51799
rect 344520 51768 344569 51796
rect 344520 51756 344526 51768
rect 344557 51765 344569 51768
rect 344603 51765 344615 51799
rect 344557 51759 344615 51765
rect 192202 51116 192208 51128
rect 192128 51088 192208 51116
rect 192128 51060 192156 51088
rect 192202 51076 192208 51088
rect 192260 51076 192266 51128
rect 224034 51076 224040 51128
rect 224092 51076 224098 51128
rect 229370 51076 229376 51128
rect 229428 51076 229434 51128
rect 232130 51116 232136 51128
rect 232056 51088 232136 51116
rect 192110 51008 192116 51060
rect 192168 51008 192174 51060
rect 224052 50992 224080 51076
rect 229388 50992 229416 51076
rect 232056 51060 232084 51088
rect 232130 51076 232136 51088
rect 232188 51076 232194 51128
rect 235258 51076 235264 51128
rect 235316 51076 235322 51128
rect 273070 51116 273076 51128
rect 272996 51088 273076 51116
rect 232038 51008 232044 51060
rect 232096 51008 232102 51060
rect 235276 51048 235304 51076
rect 272996 51060 273024 51088
rect 273070 51076 273076 51088
rect 273128 51076 273134 51128
rect 235350 51048 235356 51060
rect 235276 51020 235356 51048
rect 235350 51008 235356 51020
rect 235408 51008 235414 51060
rect 272978 51008 272984 51060
rect 273036 51008 273042 51060
rect 291838 51008 291844 51060
rect 291896 51048 291902 51060
rect 292022 51048 292028 51060
rect 291896 51020 292028 51048
rect 291896 51008 291902 51020
rect 292022 51008 292028 51020
rect 292080 51008 292086 51060
rect 224034 50940 224040 50992
rect 224092 50940 224098 50992
rect 229370 50940 229376 50992
rect 229428 50940 229434 50992
rect 2774 50124 2780 50176
rect 2832 50164 2838 50176
rect 4890 50164 4896 50176
rect 2832 50136 4896 50164
rect 2832 50124 2838 50136
rect 4890 50124 4896 50136
rect 4948 50124 4954 50176
rect 235166 48396 235172 48408
rect 235092 48368 235172 48396
rect 235092 48340 235120 48368
rect 235166 48356 235172 48368
rect 235224 48356 235230 48408
rect 354306 48396 354312 48408
rect 354267 48368 354312 48396
rect 354306 48356 354312 48368
rect 354364 48356 354370 48408
rect 200393 48331 200451 48337
rect 200393 48297 200405 48331
rect 200439 48328 200451 48331
rect 200482 48328 200488 48340
rect 200439 48300 200488 48328
rect 200439 48297 200451 48300
rect 200393 48291 200451 48297
rect 200482 48288 200488 48300
rect 200540 48288 200546 48340
rect 235074 48288 235080 48340
rect 235132 48288 235138 48340
rect 258258 48288 258264 48340
rect 258316 48328 258322 48340
rect 258350 48328 258356 48340
rect 258316 48300 258356 48328
rect 258316 48288 258322 48300
rect 258350 48288 258356 48300
rect 258408 48288 258414 48340
rect 262490 48328 262496 48340
rect 262451 48300 262496 48328
rect 262490 48288 262496 48300
rect 262548 48288 262554 48340
rect 277121 48331 277179 48337
rect 277121 48297 277133 48331
rect 277167 48328 277179 48331
rect 277210 48328 277216 48340
rect 277167 48300 277216 48328
rect 277167 48297 277179 48300
rect 277121 48291 277179 48297
rect 277210 48288 277216 48300
rect 277268 48288 277274 48340
rect 285306 48288 285312 48340
rect 285364 48328 285370 48340
rect 285398 48328 285404 48340
rect 285364 48300 285404 48328
rect 285364 48288 285370 48300
rect 285398 48288 285404 48300
rect 285456 48288 285462 48340
rect 286594 48288 286600 48340
rect 286652 48328 286658 48340
rect 286686 48328 286692 48340
rect 286652 48300 286692 48328
rect 286652 48288 286658 48300
rect 286686 48288 286692 48300
rect 286744 48288 286750 48340
rect 289354 48288 289360 48340
rect 289412 48328 289418 48340
rect 289446 48328 289452 48340
rect 289412 48300 289452 48328
rect 289412 48288 289418 48300
rect 289446 48288 289452 48300
rect 289504 48288 289510 48340
rect 355594 48328 355600 48340
rect 355555 48300 355600 48328
rect 355594 48288 355600 48300
rect 355652 48288 355658 48340
rect 362313 48331 362371 48337
rect 362313 48297 362325 48331
rect 362359 48328 362371 48331
rect 362494 48328 362500 48340
rect 362359 48300 362500 48328
rect 362359 48297 362371 48300
rect 362313 48291 362371 48297
rect 362494 48288 362500 48300
rect 362552 48288 362558 48340
rect 171410 48260 171416 48272
rect 171371 48232 171416 48260
rect 171410 48220 171416 48232
rect 171468 48220 171474 48272
rect 189442 48220 189448 48272
rect 189500 48260 189506 48272
rect 189534 48260 189540 48272
rect 189500 48232 189540 48260
rect 189500 48220 189506 48232
rect 189534 48220 189540 48232
rect 189592 48220 189598 48272
rect 211890 48220 211896 48272
rect 211948 48260 211954 48272
rect 211982 48260 211988 48272
rect 211948 48232 211988 48260
rect 211948 48220 211954 48232
rect 211982 48220 211988 48232
rect 212040 48220 212046 48272
rect 212442 48260 212448 48272
rect 212403 48232 212448 48260
rect 212442 48220 212448 48232
rect 212500 48220 212506 48272
rect 275830 48220 275836 48272
rect 275888 48260 275894 48272
rect 275922 48260 275928 48272
rect 275888 48232 275928 48260
rect 275888 48220 275894 48232
rect 275922 48220 275928 48232
rect 275980 48220 275986 48272
rect 282730 48220 282736 48272
rect 282788 48260 282794 48272
rect 282822 48260 282828 48272
rect 282788 48232 282828 48260
rect 282788 48220 282794 48232
rect 282822 48220 282828 48232
rect 282880 48220 282886 48272
rect 354306 48260 354312 48272
rect 354267 48232 354312 48260
rect 354306 48220 354312 48232
rect 354364 48220 354370 48272
rect 291746 48152 291752 48204
rect 291804 48192 291810 48204
rect 291838 48192 291844 48204
rect 291804 48164 291844 48192
rect 291804 48152 291810 48164
rect 291838 48152 291844 48164
rect 291896 48152 291902 48204
rect 270126 47404 270132 47456
rect 270184 47444 270190 47456
rect 270310 47444 270316 47456
rect 270184 47416 270316 47444
rect 270184 47404 270190 47416
rect 270310 47404 270316 47416
rect 270368 47404 270374 47456
rect 283929 46971 283987 46977
rect 283929 46937 283941 46971
rect 283975 46968 283987 46971
rect 284018 46968 284024 46980
rect 283975 46940 284024 46968
rect 283975 46937 283987 46940
rect 283929 46931 283987 46937
rect 284018 46928 284024 46940
rect 284076 46928 284082 46980
rect 318337 46971 318395 46977
rect 318337 46937 318349 46971
rect 318383 46968 318395 46971
rect 318426 46968 318432 46980
rect 318383 46940 318432 46968
rect 318383 46937 318395 46940
rect 318337 46931 318395 46937
rect 318426 46928 318432 46940
rect 318484 46928 318490 46980
rect 345658 46928 345664 46980
rect 345716 46968 345722 46980
rect 345716 46940 345761 46968
rect 345716 46928 345722 46940
rect 194962 46860 194968 46912
rect 195020 46900 195026 46912
rect 195146 46900 195152 46912
rect 195020 46872 195152 46900
rect 195020 46860 195026 46872
rect 195146 46860 195152 46872
rect 195204 46860 195210 46912
rect 228177 46903 228235 46909
rect 228177 46869 228189 46903
rect 228223 46900 228235 46903
rect 228266 46900 228272 46912
rect 228223 46872 228272 46900
rect 228223 46869 228235 46872
rect 228177 46863 228235 46869
rect 228266 46860 228272 46872
rect 228324 46860 228330 46912
rect 232038 46900 232044 46912
rect 231999 46872 232044 46900
rect 232038 46860 232044 46872
rect 232096 46860 232102 46912
rect 261202 46860 261208 46912
rect 261260 46900 261266 46912
rect 261294 46900 261300 46912
rect 261260 46872 261300 46900
rect 261260 46860 261266 46872
rect 261294 46860 261300 46872
rect 261352 46860 261358 46912
rect 317138 46900 317144 46912
rect 317099 46872 317144 46900
rect 317138 46860 317144 46872
rect 317196 46860 317202 46912
rect 179966 45636 179972 45688
rect 180024 45636 180030 45688
rect 181162 45676 181168 45688
rect 181088 45648 181168 45676
rect 179984 45549 180012 45636
rect 181088 45620 181116 45648
rect 181162 45636 181168 45648
rect 181220 45636 181226 45688
rect 181070 45568 181076 45620
rect 181128 45568 181134 45620
rect 183922 45608 183928 45620
rect 183883 45580 183928 45608
rect 183922 45568 183928 45580
rect 183980 45568 183986 45620
rect 341886 45568 341892 45620
rect 341944 45568 341950 45620
rect 179969 45543 180027 45549
rect 179969 45509 179981 45543
rect 180015 45509 180027 45543
rect 179969 45503 180027 45509
rect 201865 45543 201923 45549
rect 201865 45509 201877 45543
rect 201911 45540 201923 45543
rect 201954 45540 201960 45552
rect 201911 45512 201960 45540
rect 201911 45509 201923 45512
rect 201865 45503 201923 45509
rect 201954 45500 201960 45512
rect 202012 45500 202018 45552
rect 228174 45500 228180 45552
rect 228232 45540 228238 45552
rect 228266 45540 228272 45552
rect 228232 45512 228272 45540
rect 228232 45500 228238 45512
rect 228266 45500 228272 45512
rect 228324 45500 228330 45552
rect 231210 45500 231216 45552
rect 231268 45540 231274 45552
rect 231302 45540 231308 45552
rect 231268 45512 231308 45540
rect 231268 45500 231274 45512
rect 231302 45500 231308 45512
rect 231360 45500 231366 45552
rect 272978 45500 272984 45552
rect 273036 45540 273042 45552
rect 273073 45543 273131 45549
rect 273073 45540 273085 45543
rect 273036 45512 273085 45540
rect 273036 45500 273042 45512
rect 273073 45509 273085 45512
rect 273119 45509 273131 45543
rect 273073 45503 273131 45509
rect 341904 45484 341932 45568
rect 341886 45432 341892 45484
rect 341944 45432 341950 45484
rect 190914 44140 190920 44192
rect 190972 44180 190978 44192
rect 191098 44180 191104 44192
rect 190972 44152 191104 44180
rect 190972 44140 190978 44152
rect 191098 44140 191104 44152
rect 191156 44140 191162 44192
rect 181073 44115 181131 44121
rect 181073 44081 181085 44115
rect 181119 44112 181131 44115
rect 181346 44112 181352 44124
rect 181119 44084 181352 44112
rect 181119 44081 181131 44084
rect 181073 44075 181131 44081
rect 181346 44072 181352 44084
rect 181404 44072 181410 44124
rect 219802 42480 219808 42492
rect 219763 42452 219808 42480
rect 219802 42440 219808 42452
rect 219860 42440 219866 42492
rect 329377 42143 329435 42149
rect 329377 42109 329389 42143
rect 329423 42140 329435 42143
rect 329466 42140 329472 42152
rect 329423 42112 329472 42140
rect 329423 42109 329435 42112
rect 329377 42103 329435 42109
rect 329466 42100 329472 42112
rect 329524 42100 329530 42152
rect 182174 41460 182180 41472
rect 182135 41432 182180 41460
rect 182174 41420 182180 41432
rect 182232 41420 182238 41472
rect 234798 41420 234804 41472
rect 234856 41460 234862 41472
rect 235074 41460 235080 41472
rect 234856 41432 235080 41460
rect 234856 41420 234862 41432
rect 235074 41420 235080 41432
rect 235132 41420 235138 41472
rect 236270 41420 236276 41472
rect 236328 41420 236334 41472
rect 236288 41336 236316 41420
rect 262398 41352 262404 41404
rect 262456 41392 262462 41404
rect 262582 41392 262588 41404
rect 262456 41364 262588 41392
rect 262456 41352 262462 41364
rect 262582 41352 262588 41364
rect 262640 41352 262646 41404
rect 236270 41284 236276 41336
rect 236328 41284 236334 41336
rect 344554 41120 344560 41132
rect 344515 41092 344560 41120
rect 344554 41080 344560 41092
rect 344612 41080 344618 41132
rect 354306 41120 354312 41132
rect 354267 41092 354312 41120
rect 354306 41080 354312 41092
rect 354364 41080 354370 41132
rect 189534 40712 189540 40724
rect 189495 40684 189540 40712
rect 189534 40672 189540 40684
rect 189592 40672 189598 40724
rect 367094 40264 367100 40316
rect 367152 40304 367158 40316
rect 369946 40304 369952 40316
rect 367152 40276 369952 40304
rect 367152 40264 367158 40276
rect 369946 40264 369952 40276
rect 370004 40264 370010 40316
rect 270494 40196 270500 40248
rect 270552 40236 270558 40248
rect 275738 40236 275744 40248
rect 270552 40208 275744 40236
rect 270552 40196 270558 40208
rect 275738 40196 275744 40208
rect 275796 40196 275802 40248
rect 398742 40196 398748 40248
rect 398800 40236 398806 40248
rect 405642 40236 405648 40248
rect 398800 40208 405648 40236
rect 398800 40196 398806 40208
rect 405642 40196 405648 40208
rect 405700 40196 405706 40248
rect 212442 40060 212448 40112
rect 212500 40100 212506 40112
rect 220722 40100 220728 40112
rect 212500 40072 220728 40100
rect 212500 40060 212506 40072
rect 220722 40060 220728 40072
rect 220780 40060 220786 40112
rect 201494 39924 201500 39976
rect 201552 39964 201558 39976
rect 201862 39964 201868 39976
rect 201552 39936 201868 39964
rect 201552 39924 201558 39936
rect 201862 39924 201868 39936
rect 201920 39924 201926 39976
rect 284110 38700 284116 38752
rect 284168 38700 284174 38752
rect 284202 38700 284208 38752
rect 284260 38700 284266 38752
rect 171410 38672 171416 38684
rect 171371 38644 171416 38672
rect 171410 38632 171416 38644
rect 171468 38632 171474 38684
rect 191190 38672 191196 38684
rect 191116 38644 191196 38672
rect 191116 38616 191144 38644
rect 191190 38632 191196 38644
rect 191248 38632 191254 38684
rect 230750 38632 230756 38684
rect 230808 38672 230814 38684
rect 230934 38672 230940 38684
rect 230808 38644 230940 38672
rect 230808 38632 230814 38644
rect 230934 38632 230940 38644
rect 230992 38632 230998 38684
rect 284128 38616 284156 38700
rect 284220 38616 284248 38700
rect 191098 38564 191104 38616
rect 191156 38564 191162 38616
rect 211890 38564 211896 38616
rect 211948 38604 211954 38616
rect 211982 38604 211988 38616
rect 211948 38576 211988 38604
rect 211948 38564 211954 38576
rect 211982 38564 211988 38576
rect 212040 38564 212046 38616
rect 229278 38564 229284 38616
rect 229336 38604 229342 38616
rect 229370 38604 229376 38616
rect 229336 38576 229376 38604
rect 229336 38564 229342 38576
rect 229370 38564 229376 38576
rect 229428 38564 229434 38616
rect 235074 38564 235080 38616
rect 235132 38604 235138 38616
rect 235258 38604 235264 38616
rect 235132 38576 235264 38604
rect 235132 38564 235138 38576
rect 235258 38564 235264 38576
rect 235316 38564 235322 38616
rect 258261 38607 258319 38613
rect 258261 38573 258273 38607
rect 258307 38604 258319 38607
rect 258350 38604 258356 38616
rect 258307 38576 258356 38604
rect 258307 38573 258319 38576
rect 258261 38567 258319 38573
rect 258350 38564 258356 38576
rect 258408 38564 258414 38616
rect 275830 38604 275836 38616
rect 275791 38576 275836 38604
rect 275830 38564 275836 38576
rect 275888 38564 275894 38616
rect 284110 38564 284116 38616
rect 284168 38564 284174 38616
rect 284202 38564 284208 38616
rect 284260 38564 284266 38616
rect 344646 38604 344652 38616
rect 344607 38576 344652 38604
rect 344646 38564 344652 38576
rect 344704 38564 344710 38616
rect 283926 38496 283932 38548
rect 283984 38536 283990 38548
rect 284294 38536 284300 38548
rect 283984 38508 284300 38536
rect 283984 38496 283990 38508
rect 284294 38496 284300 38508
rect 284352 38496 284358 38548
rect 328270 37408 328276 37460
rect 328328 37408 328334 37460
rect 328288 37324 328316 37408
rect 200390 37272 200396 37324
rect 200448 37312 200454 37324
rect 200482 37312 200488 37324
rect 200448 37284 200488 37312
rect 200448 37272 200454 37284
rect 200482 37272 200488 37284
rect 200540 37272 200546 37324
rect 212350 37272 212356 37324
rect 212408 37312 212414 37324
rect 212445 37315 212503 37321
rect 212445 37312 212457 37315
rect 212408 37284 212457 37312
rect 212408 37272 212414 37284
rect 212445 37281 212457 37284
rect 212491 37281 212503 37315
rect 212445 37275 212503 37281
rect 217134 37272 217140 37324
rect 217192 37312 217198 37324
rect 217226 37312 217232 37324
rect 217192 37284 217232 37312
rect 217192 37272 217198 37284
rect 217226 37272 217232 37284
rect 217284 37272 217290 37324
rect 225230 37272 225236 37324
rect 225288 37312 225294 37324
rect 225506 37312 225512 37324
rect 225288 37284 225512 37312
rect 225288 37272 225294 37284
rect 225506 37272 225512 37284
rect 225564 37272 225570 37324
rect 232038 37312 232044 37324
rect 231999 37284 232044 37312
rect 232038 37272 232044 37284
rect 232096 37272 232102 37324
rect 282730 37272 282736 37324
rect 282788 37312 282794 37324
rect 282822 37312 282828 37324
rect 282788 37284 282828 37312
rect 282788 37272 282794 37284
rect 282822 37272 282828 37284
rect 282880 37272 282886 37324
rect 317141 37315 317199 37321
rect 317141 37281 317153 37315
rect 317187 37312 317199 37315
rect 317230 37312 317236 37324
rect 317187 37284 317236 37312
rect 317187 37281 317199 37284
rect 317141 37275 317199 37281
rect 317230 37272 317236 37284
rect 317288 37272 317294 37324
rect 328270 37272 328276 37324
rect 328328 37272 328334 37324
rect 329374 37312 329380 37324
rect 329335 37284 329380 37312
rect 329374 37272 329380 37284
rect 329432 37272 329438 37324
rect 343358 37312 343364 37324
rect 343319 37284 343364 37312
rect 343358 37272 343364 37284
rect 343416 37272 343422 37324
rect 272978 37136 272984 37188
rect 273036 37176 273042 37188
rect 273073 37179 273131 37185
rect 273073 37176 273085 37179
rect 273036 37148 273085 37176
rect 273036 37136 273042 37148
rect 273073 37145 273085 37148
rect 273119 37145 273131 37179
rect 273073 37139 273131 37145
rect 178126 35912 178132 35964
rect 178184 35952 178190 35964
rect 178218 35952 178224 35964
rect 178184 35924 178224 35952
rect 178184 35912 178190 35924
rect 178218 35912 178224 35924
rect 178276 35912 178282 35964
rect 179969 35955 180027 35961
rect 179969 35921 179981 35955
rect 180015 35952 180027 35955
rect 180058 35952 180064 35964
rect 180015 35924 180064 35952
rect 180015 35921 180027 35924
rect 179969 35915 180027 35921
rect 180058 35912 180064 35924
rect 180116 35912 180122 35964
rect 219805 35955 219863 35961
rect 219805 35921 219817 35955
rect 219851 35952 219863 35955
rect 219986 35952 219992 35964
rect 219851 35924 219992 35952
rect 219851 35921 219863 35924
rect 219805 35915 219863 35921
rect 219986 35912 219992 35924
rect 220044 35912 220050 35964
rect 2774 35844 2780 35896
rect 2832 35884 2838 35896
rect 4798 35884 4804 35896
rect 2832 35856 4804 35884
rect 2832 35844 2838 35856
rect 4798 35844 4804 35856
rect 4856 35844 4862 35896
rect 270126 35300 270132 35352
rect 270184 35340 270190 35352
rect 270310 35340 270316 35352
rect 270184 35312 270316 35340
rect 270184 35300 270190 35312
rect 270310 35300 270316 35312
rect 270368 35300 270374 35352
rect 284110 33804 284116 33856
rect 284168 33804 284174 33856
rect 318426 33804 318432 33856
rect 318484 33804 318490 33856
rect 284128 33720 284156 33804
rect 318444 33776 318472 33804
rect 318518 33776 318524 33788
rect 318444 33748 318524 33776
rect 318518 33736 318524 33748
rect 318576 33736 318582 33788
rect 284110 33668 284116 33720
rect 284168 33668 284174 33720
rect 275833 33235 275891 33241
rect 275833 33201 275845 33235
rect 275879 33232 275891 33235
rect 275922 33232 275928 33244
rect 275879 33204 275928 33232
rect 275879 33201 275891 33204
rect 275833 33195 275891 33201
rect 275922 33192 275928 33204
rect 275980 33192 275986 33244
rect 196066 31832 196072 31884
rect 196124 31832 196130 31884
rect 266538 31832 266544 31884
rect 266596 31832 266602 31884
rect 362405 31875 362463 31881
rect 362405 31841 362417 31875
rect 362451 31872 362463 31875
rect 362586 31872 362592 31884
rect 362451 31844 362592 31872
rect 362451 31841 362463 31844
rect 362405 31835 362463 31841
rect 362586 31832 362592 31844
rect 362644 31832 362650 31884
rect 178218 31804 178224 31816
rect 178144 31776 178224 31804
rect 178144 31748 178172 31776
rect 178218 31764 178224 31776
rect 178276 31764 178282 31816
rect 180058 31804 180064 31816
rect 179984 31776 180064 31804
rect 179984 31748 180012 31776
rect 180058 31764 180064 31776
rect 180116 31764 180122 31816
rect 196084 31748 196112 31832
rect 234798 31804 234804 31816
rect 234724 31776 234804 31804
rect 234724 31748 234752 31776
rect 234798 31764 234804 31776
rect 234856 31764 234862 31816
rect 266556 31748 266584 31832
rect 285398 31804 285404 31816
rect 285324 31776 285404 31804
rect 285324 31748 285352 31776
rect 285398 31764 285404 31776
rect 285456 31764 285462 31816
rect 286686 31804 286692 31816
rect 286612 31776 286692 31804
rect 286612 31748 286640 31776
rect 286686 31764 286692 31776
rect 286744 31764 286750 31816
rect 291838 31764 291844 31816
rect 291896 31764 291902 31816
rect 328089 31807 328147 31813
rect 328089 31773 328101 31807
rect 328135 31804 328147 31807
rect 328178 31804 328184 31816
rect 328135 31776 328184 31804
rect 328135 31773 328147 31776
rect 328089 31767 328147 31773
rect 328178 31764 328184 31776
rect 328236 31764 328242 31816
rect 361301 31807 361359 31813
rect 361301 31773 361313 31807
rect 361347 31804 361359 31807
rect 361390 31804 361396 31816
rect 361347 31776 361396 31804
rect 361347 31773 361359 31776
rect 361301 31767 361359 31773
rect 361390 31764 361396 31776
rect 361448 31764 361454 31816
rect 178126 31696 178132 31748
rect 178184 31696 178190 31748
rect 179966 31696 179972 31748
rect 180024 31696 180030 31748
rect 196066 31696 196072 31748
rect 196124 31696 196130 31748
rect 234706 31696 234712 31748
rect 234764 31696 234770 31748
rect 258258 31736 258264 31748
rect 258219 31708 258264 31736
rect 258258 31696 258264 31708
rect 258316 31696 258322 31748
rect 266538 31696 266544 31748
rect 266596 31696 266602 31748
rect 285306 31696 285312 31748
rect 285364 31696 285370 31748
rect 286594 31696 286600 31748
rect 286652 31696 286658 31748
rect 291856 31736 291884 31764
rect 291930 31736 291936 31748
rect 291856 31708 291936 31736
rect 291930 31696 291936 31708
rect 291988 31696 291994 31748
rect 370498 30268 370504 30320
rect 370556 30308 370562 30320
rect 580258 30308 580264 30320
rect 370556 30280 580264 30308
rect 370556 30268 370562 30280
rect 580258 30268 580264 30280
rect 580316 30268 580322 30320
rect 231302 29084 231308 29096
rect 231136 29056 231308 29084
rect 231136 28960 231164 29056
rect 231302 29044 231308 29056
rect 231360 29044 231366 29096
rect 232038 28976 232044 29028
rect 232096 29016 232102 29028
rect 232130 29016 232136 29028
rect 232096 28988 232136 29016
rect 232096 28976 232102 28988
rect 232130 28976 232136 28988
rect 232188 28976 232194 29028
rect 261110 28976 261116 29028
rect 261168 29016 261174 29028
rect 261202 29016 261208 29028
rect 261168 28988 261208 29016
rect 261168 28976 261174 28988
rect 261202 28976 261208 28988
rect 261260 28976 261266 29028
rect 284018 28976 284024 29028
rect 284076 29016 284082 29028
rect 284294 29016 284300 29028
rect 284076 28988 284300 29016
rect 284076 28976 284082 28988
rect 284294 28976 284300 28988
rect 284352 28976 284358 29028
rect 289262 28976 289268 29028
rect 289320 29016 289326 29028
rect 289446 29016 289452 29028
rect 289320 28988 289452 29016
rect 289320 28976 289326 28988
rect 289446 28976 289452 28988
rect 289504 28976 289510 29028
rect 317138 28976 317144 29028
rect 317196 29016 317202 29028
rect 317230 29016 317236 29028
rect 317196 28988 317236 29016
rect 317196 28976 317202 28988
rect 317230 28976 317236 28988
rect 317288 28976 317294 29028
rect 344646 29016 344652 29028
rect 344607 28988 344652 29016
rect 344646 28976 344652 28988
rect 344704 28976 344710 29028
rect 361298 29016 361304 29028
rect 361259 28988 361304 29016
rect 361298 28976 361304 28988
rect 361356 28976 361362 29028
rect 362402 29016 362408 29028
rect 362363 28988 362408 29016
rect 362402 28976 362408 28988
rect 362460 28976 362466 29028
rect 171321 28951 171379 28957
rect 171321 28917 171333 28951
rect 171367 28948 171379 28951
rect 171410 28948 171416 28960
rect 171367 28920 171416 28948
rect 171367 28917 171379 28920
rect 171321 28911 171379 28917
rect 171410 28908 171416 28920
rect 171468 28908 171474 28960
rect 173066 28908 173072 28960
rect 173124 28948 173130 28960
rect 173158 28948 173164 28960
rect 173124 28920 173164 28948
rect 173124 28908 173130 28920
rect 173158 28908 173164 28920
rect 173216 28908 173222 28960
rect 184014 28908 184020 28960
rect 184072 28948 184078 28960
rect 184106 28948 184112 28960
rect 184072 28920 184112 28948
rect 184072 28908 184078 28920
rect 184106 28908 184112 28920
rect 184164 28908 184170 28960
rect 203150 28908 203156 28960
rect 203208 28948 203214 28960
rect 203242 28948 203248 28960
rect 203208 28920 203248 28948
rect 203208 28908 203214 28920
rect 203242 28908 203248 28920
rect 203300 28908 203306 28960
rect 231118 28908 231124 28960
rect 231176 28908 231182 28960
rect 236362 28948 236368 28960
rect 236323 28920 236368 28948
rect 236362 28908 236368 28920
rect 236420 28908 236426 28960
rect 329466 28948 329472 28960
rect 329427 28920 329472 28948
rect 329466 28908 329472 28920
rect 329524 28908 329530 28960
rect 317138 28880 317144 28892
rect 317099 28852 317144 28880
rect 317138 28840 317144 28852
rect 317196 28840 317202 28892
rect 343358 28472 343364 28484
rect 343319 28444 343364 28472
rect 343358 28432 343364 28444
rect 343416 28432 343422 28484
rect 272978 27684 272984 27736
rect 273036 27724 273042 27736
rect 273036 27696 273116 27724
rect 273036 27684 273042 27696
rect 273088 27668 273116 27696
rect 182174 27616 182180 27668
rect 182232 27656 182238 27668
rect 189534 27656 189540 27668
rect 182232 27628 182277 27656
rect 189495 27628 189540 27656
rect 182232 27616 182238 27628
rect 189534 27616 189540 27628
rect 189592 27616 189598 27668
rect 200390 27656 200396 27668
rect 200351 27628 200396 27656
rect 200390 27616 200396 27628
rect 200448 27616 200454 27668
rect 201862 27656 201868 27668
rect 201823 27628 201868 27656
rect 201862 27616 201868 27628
rect 201920 27616 201926 27668
rect 219802 27616 219808 27668
rect 219860 27656 219866 27668
rect 219986 27656 219992 27668
rect 219860 27628 219992 27656
rect 219860 27616 219866 27628
rect 219986 27616 219992 27628
rect 220044 27616 220050 27668
rect 273070 27616 273076 27668
rect 273128 27616 273134 27668
rect 328086 27656 328092 27668
rect 328047 27628 328092 27656
rect 328086 27616 328092 27628
rect 328144 27616 328150 27668
rect 212074 27548 212080 27600
rect 212132 27588 212138 27600
rect 212166 27588 212172 27600
rect 212132 27560 212172 27588
rect 212132 27548 212138 27560
rect 212166 27548 212172 27560
rect 212224 27548 212230 27600
rect 212258 27548 212264 27600
rect 212316 27588 212322 27600
rect 261110 27588 261116 27600
rect 212316 27560 212361 27588
rect 261071 27560 261116 27588
rect 212316 27548 212322 27560
rect 261110 27548 261116 27560
rect 261168 27548 261174 27600
rect 268746 27588 268752 27600
rect 268707 27560 268752 27588
rect 268746 27548 268752 27560
rect 268804 27548 268810 27600
rect 275922 27588 275928 27600
rect 275883 27560 275928 27588
rect 275922 27548 275928 27560
rect 275980 27548 275986 27600
rect 277121 27591 277179 27597
rect 277121 27557 277133 27591
rect 277167 27588 277179 27591
rect 277210 27588 277216 27600
rect 277167 27560 277216 27588
rect 277167 27557 277179 27560
rect 277121 27551 277179 27557
rect 277210 27548 277216 27560
rect 277268 27548 277274 27600
rect 343269 27591 343327 27597
rect 343269 27557 343281 27591
rect 343315 27588 343327 27591
rect 343358 27588 343364 27600
rect 343315 27560 343364 27588
rect 343315 27557 343327 27560
rect 343269 27551 343327 27557
rect 343358 27548 343364 27560
rect 343416 27548 343422 27600
rect 344557 27591 344615 27597
rect 344557 27557 344569 27591
rect 344603 27588 344615 27591
rect 344646 27588 344652 27600
rect 344603 27560 344652 27588
rect 344603 27557 344615 27560
rect 344557 27551 344615 27557
rect 344646 27548 344652 27560
rect 344704 27548 344710 27600
rect 345658 27588 345664 27600
rect 345619 27560 345664 27588
rect 345658 27548 345664 27560
rect 345716 27548 345722 27600
rect 354309 27591 354367 27597
rect 354309 27557 354321 27591
rect 354355 27588 354367 27591
rect 354398 27588 354404 27600
rect 354355 27560 354404 27588
rect 354355 27557 354367 27560
rect 354309 27551 354367 27557
rect 354398 27548 354404 27560
rect 354456 27548 354462 27600
rect 355505 27591 355563 27597
rect 355505 27557 355517 27591
rect 355551 27588 355563 27591
rect 355686 27588 355692 27600
rect 355551 27560 355692 27588
rect 355551 27557 355563 27560
rect 355505 27551 355563 27557
rect 355686 27548 355692 27560
rect 355744 27548 355750 27600
rect 361209 27591 361267 27597
rect 361209 27557 361221 27591
rect 361255 27588 361267 27591
rect 361298 27588 361304 27600
rect 361255 27560 361304 27588
rect 361255 27557 361267 27560
rect 361209 27551 361267 27557
rect 361298 27548 361304 27560
rect 361356 27548 361362 27600
rect 270126 26868 270132 26920
rect 270184 26908 270190 26920
rect 270310 26908 270316 26920
rect 270184 26880 270316 26908
rect 270184 26868 270190 26880
rect 270310 26868 270316 26880
rect 270368 26868 270374 26920
rect 230934 26596 230940 26648
rect 230992 26636 230998 26648
rect 231118 26636 231124 26648
rect 230992 26608 231124 26636
rect 230992 26596 230998 26608
rect 231118 26596 231124 26608
rect 231176 26596 231182 26648
rect 181070 26296 181076 26308
rect 181031 26268 181076 26296
rect 181070 26256 181076 26268
rect 181128 26256 181134 26308
rect 200390 26296 200396 26308
rect 200351 26268 200396 26296
rect 200390 26256 200396 26268
rect 200448 26256 200454 26308
rect 178126 26228 178132 26240
rect 178087 26200 178132 26228
rect 178126 26188 178132 26200
rect 178184 26188 178190 26240
rect 179966 26228 179972 26240
rect 179927 26200 179972 26228
rect 179966 26188 179972 26200
rect 180024 26188 180030 26240
rect 182174 26188 182180 26240
rect 182232 26228 182238 26240
rect 182450 26228 182456 26240
rect 182232 26200 182456 26228
rect 182232 26188 182238 26200
rect 182450 26188 182456 26200
rect 182508 26188 182514 26240
rect 194870 26228 194876 26240
rect 194831 26200 194876 26228
rect 194870 26188 194876 26200
rect 194928 26188 194934 26240
rect 181162 26120 181168 26172
rect 181220 26160 181226 26172
rect 181346 26160 181352 26172
rect 181220 26132 181352 26160
rect 181220 26120 181226 26132
rect 181346 26120 181352 26132
rect 181404 26120 181410 26172
rect 234706 25100 234712 25152
rect 234764 25140 234770 25152
rect 235166 25140 235172 25152
rect 234764 25112 235172 25140
rect 234764 25100 234770 25112
rect 235166 25100 235172 25112
rect 235224 25100 235230 25152
rect 266538 23604 266544 23656
rect 266596 23644 266602 23656
rect 266814 23644 266820 23656
rect 266596 23616 266820 23644
rect 266596 23604 266602 23616
rect 266814 23604 266820 23616
rect 266872 23604 266878 23656
rect 200390 22108 200396 22160
rect 200448 22108 200454 22160
rect 217134 22108 217140 22160
rect 217192 22108 217198 22160
rect 291930 22108 291936 22160
rect 291988 22108 291994 22160
rect 200408 22024 200436 22108
rect 214098 22040 214104 22092
rect 214156 22080 214162 22092
rect 214282 22080 214288 22092
rect 214156 22052 214288 22080
rect 214156 22040 214162 22052
rect 214282 22040 214288 22052
rect 214340 22040 214346 22092
rect 217152 22024 217180 22108
rect 262398 22040 262404 22092
rect 262456 22080 262462 22092
rect 262582 22080 262588 22092
rect 262456 22052 262588 22080
rect 262456 22040 262462 22052
rect 262582 22040 262588 22052
rect 262640 22040 262646 22092
rect 291948 22024 291976 22108
rect 200390 21972 200396 22024
rect 200448 21972 200454 22024
rect 217134 21972 217140 22024
rect 217192 21972 217198 22024
rect 291930 21972 291936 22024
rect 291988 21972 291994 22024
rect 171318 19360 171324 19372
rect 171279 19332 171324 19360
rect 171318 19320 171324 19332
rect 171376 19320 171382 19372
rect 223942 19320 223948 19372
rect 224000 19360 224006 19372
rect 224034 19360 224040 19372
rect 224000 19332 224040 19360
rect 224000 19320 224006 19332
rect 224034 19320 224040 19332
rect 224092 19320 224098 19372
rect 229278 19320 229284 19372
rect 229336 19360 229342 19372
rect 229370 19360 229376 19372
rect 229336 19332 229376 19360
rect 229336 19320 229342 19332
rect 229370 19320 229376 19332
rect 229428 19320 229434 19372
rect 236362 19360 236368 19372
rect 236323 19332 236368 19360
rect 236362 19320 236368 19332
rect 236420 19320 236426 19372
rect 317141 19363 317199 19369
rect 317141 19329 317153 19363
rect 317187 19360 317199 19363
rect 317230 19360 317236 19372
rect 317187 19332 317236 19360
rect 317187 19329 317199 19332
rect 317141 19323 317199 19329
rect 317230 19320 317236 19332
rect 317288 19320 317294 19372
rect 329469 19363 329527 19369
rect 329469 19329 329481 19363
rect 329515 19360 329527 19363
rect 329558 19360 329564 19372
rect 329515 19332 329564 19360
rect 329515 19329 329527 19332
rect 329469 19323 329527 19329
rect 329558 19320 329564 19332
rect 329616 19320 329622 19372
rect 192113 19295 192171 19301
rect 192113 19261 192125 19295
rect 192159 19292 192171 19295
rect 192202 19292 192208 19304
rect 192159 19264 192208 19292
rect 192159 19261 192171 19264
rect 192113 19255 192171 19261
rect 192202 19252 192208 19264
rect 192260 19252 192266 19304
rect 212258 19292 212264 19304
rect 212219 19264 212264 19292
rect 212258 19252 212264 19264
rect 212316 19252 212322 19304
rect 214282 19292 214288 19304
rect 214243 19264 214288 19292
rect 214282 19252 214288 19264
rect 214340 19252 214346 19304
rect 291841 19295 291899 19301
rect 291841 19261 291853 19295
rect 291887 19292 291899 19295
rect 291930 19292 291936 19304
rect 291887 19264 291936 19292
rect 291887 19261 291899 19264
rect 291841 19255 291899 19261
rect 291930 19252 291936 19264
rect 291988 19252 291994 19304
rect 328181 19295 328239 19301
rect 328181 19261 328193 19295
rect 328227 19292 328239 19295
rect 328270 19292 328276 19304
rect 328227 19264 328276 19292
rect 328227 19261 328239 19264
rect 328181 19255 328239 19261
rect 328270 19252 328276 19264
rect 328328 19252 328334 19304
rect 352926 19292 352932 19304
rect 352887 19264 352932 19292
rect 352926 19252 352932 19264
rect 352984 19252 352990 19304
rect 362497 19295 362555 19301
rect 362497 19261 362509 19295
rect 362543 19292 362555 19295
rect 362586 19292 362592 19304
rect 362543 19264 362592 19292
rect 362543 19261 362555 19264
rect 362497 19255 362555 19261
rect 362586 19252 362592 19264
rect 362644 19252 362650 19304
rect 341886 18408 341892 18420
rect 341847 18380 341892 18408
rect 341886 18368 341892 18380
rect 341944 18368 341950 18420
rect 219710 18028 219716 18080
rect 219768 18068 219774 18080
rect 219768 18040 219848 18068
rect 219768 18028 219774 18040
rect 219820 18012 219848 18040
rect 182358 18000 182364 18012
rect 182319 17972 182364 18000
rect 182358 17960 182364 17972
rect 182416 17960 182422 18012
rect 219802 17960 219808 18012
rect 219860 17960 219866 18012
rect 261110 18000 261116 18012
rect 261071 17972 261116 18000
rect 261110 17960 261116 17972
rect 261168 17960 261174 18012
rect 268746 18000 268752 18012
rect 268707 17972 268752 18000
rect 268746 17960 268752 17972
rect 268804 17960 268810 18012
rect 272794 17960 272800 18012
rect 272852 18000 272858 18012
rect 272886 18000 272892 18012
rect 272852 17972 272892 18000
rect 272852 17960 272858 17972
rect 272886 17960 272892 17972
rect 272944 17960 272950 18012
rect 275922 18000 275928 18012
rect 275883 17972 275928 18000
rect 275922 17960 275928 17972
rect 275980 17960 275986 18012
rect 345658 18000 345664 18012
rect 345619 17972 345664 18000
rect 345658 17960 345664 17972
rect 345716 17960 345722 18012
rect 354306 18000 354312 18012
rect 354267 17972 354312 18000
rect 354306 17960 354312 17972
rect 354364 17960 354370 18012
rect 355502 18000 355508 18012
rect 355463 17972 355508 18000
rect 355502 17960 355508 17972
rect 355560 17960 355566 18012
rect 361206 18000 361212 18012
rect 361167 17972 361212 18000
rect 361206 17960 361212 17972
rect 361264 17960 361270 18012
rect 169754 17892 169760 17944
rect 169812 17932 169818 17944
rect 228085 17935 228143 17941
rect 228085 17932 228097 17935
rect 169812 17904 182220 17932
rect 169812 17892 169818 17904
rect 182192 17864 182220 17904
rect 184676 17904 228097 17932
rect 184676 17864 184704 17904
rect 228085 17901 228097 17904
rect 228131 17901 228143 17935
rect 228085 17895 228143 17901
rect 228269 17935 228327 17941
rect 228269 17901 228281 17935
rect 228315 17932 228327 17935
rect 579614 17932 579620 17944
rect 228315 17904 579620 17932
rect 228315 17901 228327 17904
rect 228269 17895 228327 17901
rect 579614 17892 579620 17904
rect 579672 17892 579678 17944
rect 182192 17836 184704 17864
rect 182358 17796 182364 17808
rect 182319 17768 182364 17796
rect 182358 17756 182364 17768
rect 182416 17756 182422 17808
rect 270126 17212 270132 17264
rect 270184 17252 270190 17264
rect 270310 17252 270316 17264
rect 270184 17224 270316 17252
rect 270184 17212 270190 17224
rect 270310 17212 270316 17224
rect 270368 17212 270374 17264
rect 230566 16736 230572 16788
rect 230624 16776 230630 16788
rect 230750 16776 230756 16788
rect 230624 16748 230756 16776
rect 230624 16736 230630 16748
rect 230750 16736 230756 16748
rect 230808 16736 230814 16788
rect 177114 16708 177120 16720
rect 177040 16680 177120 16708
rect 177040 16652 177068 16680
rect 177114 16668 177120 16680
rect 177172 16668 177178 16720
rect 177022 16600 177028 16652
rect 177080 16600 177086 16652
rect 178126 16640 178132 16652
rect 178087 16612 178132 16640
rect 178126 16600 178132 16612
rect 178184 16600 178190 16652
rect 179966 16640 179972 16652
rect 179927 16612 179972 16640
rect 179966 16600 179972 16612
rect 180024 16600 180030 16652
rect 194873 16643 194931 16649
rect 194873 16609 194885 16643
rect 194919 16640 194931 16643
rect 194962 16640 194968 16652
rect 194919 16612 194968 16640
rect 194919 16609 194931 16612
rect 194873 16603 194931 16609
rect 194962 16600 194968 16612
rect 195020 16600 195026 16652
rect 296438 14696 296444 14748
rect 296496 14736 296502 14748
rect 367094 14736 367100 14748
rect 296496 14708 367100 14736
rect 296496 14696 296502 14708
rect 367094 14696 367100 14708
rect 367152 14696 367158 14748
rect 297726 14628 297732 14680
rect 297784 14668 297790 14680
rect 371234 14668 371240 14680
rect 297784 14640 371240 14668
rect 297784 14628 297790 14640
rect 371234 14628 371240 14640
rect 371292 14628 371298 14680
rect 299106 14560 299112 14612
rect 299164 14600 299170 14612
rect 375190 14600 375196 14612
rect 299164 14572 375196 14600
rect 299164 14560 299170 14572
rect 375190 14560 375196 14572
rect 375248 14560 375254 14612
rect 300394 14492 300400 14544
rect 300452 14532 300458 14544
rect 378134 14532 378140 14544
rect 300452 14504 378140 14532
rect 300452 14492 300458 14504
rect 378134 14492 378140 14504
rect 378192 14492 378198 14544
rect 358538 14424 358544 14476
rect 358596 14464 358602 14476
rect 546494 14464 546500 14476
rect 358596 14436 546500 14464
rect 358596 14424 358602 14436
rect 546494 14424 546500 14436
rect 546552 14424 546558 14476
rect 341889 13787 341947 13793
rect 341889 13753 341901 13787
rect 341935 13784 341947 13787
rect 499574 13784 499580 13796
rect 341935 13756 499580 13784
rect 341935 13753 341947 13756
rect 341889 13747 341947 13753
rect 499574 13744 499580 13756
rect 499632 13744 499638 13796
rect 343269 13719 343327 13725
rect 343269 13685 343281 13719
rect 343315 13716 343327 13719
rect 502334 13716 502340 13728
rect 343315 13688 502340 13716
rect 343315 13685 343327 13688
rect 343269 13679 343327 13685
rect 502334 13676 502340 13688
rect 502392 13676 502398 13728
rect 344557 13651 344615 13657
rect 344557 13617 344569 13651
rect 344603 13648 344615 13651
rect 506474 13648 506480 13660
rect 344603 13620 506480 13648
rect 344603 13617 344615 13620
rect 344557 13611 344615 13617
rect 506474 13608 506480 13620
rect 506532 13608 506538 13660
rect 346118 13540 346124 13592
rect 346176 13580 346182 13592
rect 510614 13580 510620 13592
rect 346176 13552 510620 13580
rect 346176 13540 346182 13552
rect 510614 13540 510620 13552
rect 510672 13540 510678 13592
rect 347406 13472 347412 13524
rect 347464 13512 347470 13524
rect 517514 13512 517520 13524
rect 347464 13484 517520 13512
rect 347464 13472 347470 13484
rect 517514 13472 517520 13484
rect 517572 13472 517578 13524
rect 348878 13404 348884 13456
rect 348936 13444 348942 13456
rect 520274 13444 520280 13456
rect 348936 13416 520280 13444
rect 348936 13404 348942 13416
rect 520274 13404 520280 13416
rect 520332 13404 520338 13456
rect 350258 13336 350264 13388
rect 350316 13376 350322 13388
rect 524414 13376 524420 13388
rect 350316 13348 524420 13376
rect 350316 13336 350322 13348
rect 524414 13336 524420 13348
rect 524472 13336 524478 13388
rect 351546 13268 351552 13320
rect 351604 13308 351610 13320
rect 528554 13308 528560 13320
rect 351604 13280 528560 13308
rect 351604 13268 351610 13280
rect 528554 13268 528560 13280
rect 528612 13268 528618 13320
rect 354306 13200 354312 13252
rect 354364 13240 354370 13252
rect 535454 13240 535460 13252
rect 354364 13212 535460 13240
rect 354364 13200 354370 13212
rect 535454 13200 535460 13212
rect 535512 13200 535518 13252
rect 355502 13132 355508 13184
rect 355560 13172 355566 13184
rect 538214 13172 538220 13184
rect 355560 13144 538220 13172
rect 355560 13132 355566 13144
rect 538214 13132 538220 13144
rect 538272 13132 538278 13184
rect 289262 13104 289268 13116
rect 289223 13076 289268 13104
rect 289262 13064 289268 13076
rect 289320 13064 289326 13116
rect 357158 13064 357164 13116
rect 357216 13104 357222 13116
rect 542354 13104 542360 13116
rect 357216 13076 542360 13104
rect 357216 13064 357222 13076
rect 542354 13064 542360 13076
rect 542412 13064 542418 13116
rect 340506 12996 340512 13048
rect 340564 13036 340570 13048
rect 495434 13036 495440 13048
rect 340564 13008 495440 13036
rect 340564 12996 340570 13008
rect 495434 12996 495440 13008
rect 495492 12996 495498 13048
rect 339218 12928 339224 12980
rect 339276 12968 339282 12980
rect 492674 12968 492680 12980
rect 339276 12940 492680 12968
rect 339276 12928 339282 12940
rect 492674 12928 492680 12940
rect 492732 12928 492738 12980
rect 337838 12860 337844 12912
rect 337896 12900 337902 12912
rect 488534 12900 488540 12912
rect 337896 12872 488540 12900
rect 337896 12860 337902 12872
rect 488534 12860 488540 12872
rect 488592 12860 488598 12912
rect 337746 12792 337752 12844
rect 337804 12832 337810 12844
rect 485774 12832 485780 12844
rect 337804 12804 485780 12832
rect 337804 12792 337810 12804
rect 485774 12792 485780 12804
rect 485832 12792 485838 12844
rect 335170 12724 335176 12776
rect 335228 12764 335234 12776
rect 480254 12764 480260 12776
rect 335228 12736 480260 12764
rect 335228 12724 335234 12736
rect 480254 12724 480260 12736
rect 480312 12724 480318 12776
rect 333606 12656 333612 12708
rect 333664 12696 333670 12708
rect 477586 12696 477592 12708
rect 333664 12668 477592 12696
rect 333664 12656 333670 12668
rect 477586 12656 477592 12668
rect 477644 12656 477650 12708
rect 212258 12560 212264 12572
rect 212219 12532 212264 12560
rect 212258 12520 212264 12532
rect 212316 12520 212322 12572
rect 234706 12452 234712 12504
rect 234764 12492 234770 12504
rect 235166 12492 235172 12504
rect 234764 12464 235172 12492
rect 234764 12452 234770 12464
rect 235166 12452 235172 12464
rect 235224 12452 235230 12504
rect 285398 12492 285404 12504
rect 285324 12464 285404 12492
rect 285324 12436 285352 12464
rect 285398 12452 285404 12464
rect 285456 12452 285462 12504
rect 286686 12492 286692 12504
rect 286612 12464 286692 12492
rect 286612 12436 286640 12464
rect 286686 12452 286692 12464
rect 286744 12452 286750 12504
rect 329466 12492 329472 12504
rect 329427 12464 329472 12492
rect 329466 12452 329472 12464
rect 329524 12452 329530 12504
rect 171134 12384 171140 12436
rect 171192 12424 171198 12436
rect 171318 12424 171324 12436
rect 171192 12396 171324 12424
rect 171192 12384 171198 12396
rect 171318 12384 171324 12396
rect 171376 12384 171382 12436
rect 211890 12384 211896 12436
rect 211948 12424 211954 12436
rect 212166 12424 212172 12436
rect 211948 12396 212172 12424
rect 211948 12384 211954 12396
rect 212166 12384 212172 12396
rect 212224 12384 212230 12436
rect 265250 12384 265256 12436
rect 265308 12424 265314 12436
rect 265802 12424 265808 12436
rect 265308 12396 265808 12424
rect 265308 12384 265314 12396
rect 265802 12384 265808 12396
rect 265860 12384 265866 12436
rect 285306 12384 285312 12436
rect 285364 12384 285370 12436
rect 286594 12384 286600 12436
rect 286652 12384 286658 12436
rect 332410 12384 332416 12436
rect 332468 12424 332474 12436
rect 469214 12424 469220 12436
rect 332468 12396 469220 12424
rect 332468 12384 332474 12396
rect 469214 12384 469220 12396
rect 469272 12384 469278 12436
rect 333698 12316 333704 12368
rect 333756 12356 333762 12368
rect 473354 12356 473360 12368
rect 333756 12328 473360 12356
rect 333756 12316 333762 12328
rect 473354 12316 473360 12328
rect 473412 12316 473418 12368
rect 335262 12248 335268 12300
rect 335320 12288 335326 12300
rect 478874 12288 478880 12300
rect 335320 12260 478880 12288
rect 335320 12248 335326 12260
rect 478874 12248 478880 12260
rect 478932 12248 478938 12300
rect 336458 12180 336464 12232
rect 336516 12220 336522 12232
rect 484394 12220 484400 12232
rect 336516 12192 484400 12220
rect 336516 12180 336522 12192
rect 484394 12180 484400 12192
rect 484452 12180 484458 12232
rect 337930 12112 337936 12164
rect 337988 12152 337994 12164
rect 487154 12152 487160 12164
rect 337988 12124 487160 12152
rect 337988 12112 337994 12124
rect 487154 12112 487160 12124
rect 487212 12112 487218 12164
rect 339310 12044 339316 12096
rect 339368 12084 339374 12096
rect 491294 12084 491300 12096
rect 339368 12056 491300 12084
rect 339368 12044 339374 12056
rect 491294 12044 491300 12056
rect 491352 12044 491358 12096
rect 340598 11976 340604 12028
rect 340656 12016 340662 12028
rect 494054 12016 494060 12028
rect 340656 11988 494060 12016
rect 340656 11976 340662 11988
rect 494054 11976 494060 11988
rect 494112 11976 494118 12028
rect 342070 11908 342076 11960
rect 342128 11948 342134 11960
rect 498194 11948 498200 11960
rect 342128 11920 498200 11948
rect 342128 11908 342134 11920
rect 498194 11908 498200 11920
rect 498252 11908 498258 11960
rect 125502 11840 125508 11892
rect 125560 11880 125566 11892
rect 212718 11880 212724 11892
rect 125560 11852 212724 11880
rect 125560 11840 125566 11852
rect 212718 11840 212724 11852
rect 212776 11840 212782 11892
rect 343450 11840 343456 11892
rect 343508 11880 343514 11892
rect 502426 11880 502432 11892
rect 343508 11852 502432 11880
rect 343508 11840 343514 11852
rect 502426 11840 502432 11852
rect 502484 11840 502490 11892
rect 121362 11772 121368 11824
rect 121420 11812 121426 11824
rect 211246 11812 211252 11824
rect 121420 11784 211252 11812
rect 121420 11772 121426 11784
rect 211246 11772 211252 11784
rect 211304 11772 211310 11824
rect 344738 11772 344744 11824
rect 344796 11812 344802 11824
rect 505094 11812 505100 11824
rect 344796 11784 505100 11812
rect 344796 11772 344802 11784
rect 505094 11772 505100 11784
rect 505152 11772 505158 11824
rect 31662 11704 31668 11756
rect 31720 11744 31726 11756
rect 180978 11744 180984 11756
rect 31720 11716 180984 11744
rect 31720 11704 31726 11716
rect 180978 11704 180984 11716
rect 181036 11704 181042 11756
rect 352929 11747 352987 11753
rect 352929 11713 352941 11747
rect 352975 11744 352987 11747
rect 531314 11744 531320 11756
rect 352975 11716 531320 11744
rect 352975 11713 352987 11716
rect 352929 11707 352987 11713
rect 531314 11704 531320 11716
rect 531372 11704 531378 11756
rect 304810 11636 304816 11688
rect 304868 11676 304874 11688
rect 390554 11676 390560 11688
rect 304868 11648 390560 11676
rect 304868 11636 304874 11648
rect 390554 11636 390560 11648
rect 390612 11636 390618 11688
rect 303430 11568 303436 11620
rect 303488 11608 303494 11620
rect 387794 11608 387800 11620
rect 303488 11580 387800 11608
rect 303488 11568 303494 11580
rect 387794 11568 387800 11580
rect 387852 11568 387858 11620
rect 302050 11500 302056 11552
rect 302108 11540 302114 11552
rect 383654 11540 383660 11552
rect 302108 11512 383660 11540
rect 302108 11500 302114 11512
rect 383654 11500 383660 11512
rect 383712 11500 383718 11552
rect 300670 11432 300676 11484
rect 300728 11472 300734 11484
rect 380894 11472 380900 11484
rect 300728 11444 380900 11472
rect 300728 11432 300734 11444
rect 380894 11432 380900 11444
rect 380952 11432 380958 11484
rect 300578 11364 300584 11416
rect 300636 11404 300642 11416
rect 376754 11404 376760 11416
rect 300636 11376 376760 11404
rect 300636 11364 300642 11376
rect 376754 11364 376760 11376
rect 376812 11364 376818 11416
rect 299290 11296 299296 11348
rect 299348 11336 299354 11348
rect 374086 11336 374092 11348
rect 299348 11308 374092 11336
rect 299348 11296 299354 11308
rect 374086 11296 374092 11308
rect 374144 11296 374150 11348
rect 297818 11228 297824 11280
rect 297876 11268 297882 11280
rect 369854 11268 369860 11280
rect 297876 11240 369860 11268
rect 297876 11228 297882 11240
rect 369854 11228 369860 11240
rect 369912 11228 369918 11280
rect 366726 11024 366732 11076
rect 366784 11064 366790 11076
rect 367002 11064 367008 11076
rect 366784 11036 367008 11064
rect 366784 11024 366790 11036
rect 367002 11024 367008 11036
rect 367060 11024 367066 11076
rect 103422 10956 103428 11008
rect 103480 10996 103486 11008
rect 204346 10996 204352 11008
rect 103480 10968 204352 10996
rect 103480 10956 103486 10968
rect 204346 10956 204352 10968
rect 204404 10956 204410 11008
rect 307570 10956 307576 11008
rect 307628 10996 307634 11008
rect 397454 10996 397460 11008
rect 307628 10968 397460 10996
rect 307628 10956 307634 10968
rect 397454 10956 397460 10968
rect 397512 10956 397518 11008
rect 99282 10888 99288 10940
rect 99340 10928 99346 10940
rect 202966 10928 202972 10940
rect 99340 10900 202972 10928
rect 99340 10888 99346 10900
rect 202966 10888 202972 10900
rect 203024 10888 203030 10940
rect 308858 10888 308864 10940
rect 308916 10928 308922 10940
rect 400306 10928 400312 10940
rect 308916 10900 400312 10928
rect 308916 10888 308922 10900
rect 400306 10888 400312 10900
rect 400364 10888 400370 10940
rect 96522 10820 96528 10872
rect 96580 10860 96586 10872
rect 201678 10860 201684 10872
rect 96580 10832 201684 10860
rect 96580 10820 96586 10832
rect 201678 10820 201684 10832
rect 201736 10820 201742 10872
rect 336550 10820 336556 10872
rect 336608 10860 336614 10872
rect 483014 10860 483020 10872
rect 336608 10832 483020 10860
rect 336608 10820 336614 10832
rect 483014 10820 483020 10832
rect 483072 10820 483078 10872
rect 92382 10752 92388 10804
rect 92440 10792 92446 10804
rect 201586 10792 201592 10804
rect 92440 10764 201592 10792
rect 92440 10752 92446 10764
rect 201586 10752 201592 10764
rect 201644 10752 201650 10804
rect 338022 10752 338028 10804
rect 338080 10792 338086 10804
rect 485866 10792 485872 10804
rect 338080 10764 485872 10792
rect 338080 10752 338086 10764
rect 485866 10752 485872 10764
rect 485924 10752 485930 10804
rect 89622 10684 89628 10736
rect 89680 10724 89686 10736
rect 200206 10724 200212 10736
rect 89680 10696 200212 10724
rect 89680 10684 89686 10696
rect 200206 10684 200212 10696
rect 200264 10684 200270 10736
rect 339402 10684 339408 10736
rect 339460 10724 339466 10736
rect 489914 10724 489920 10736
rect 339460 10696 489920 10724
rect 339460 10684 339466 10696
rect 489914 10684 489920 10696
rect 489972 10684 489978 10736
rect 85482 10616 85488 10668
rect 85540 10656 85546 10668
rect 198918 10656 198924 10668
rect 85540 10628 198924 10656
rect 85540 10616 85546 10628
rect 198918 10616 198924 10628
rect 198976 10616 198982 10668
rect 340782 10616 340788 10668
rect 340840 10656 340846 10668
rect 494146 10656 494152 10668
rect 340840 10628 494152 10656
rect 340840 10616 340846 10628
rect 494146 10616 494152 10628
rect 494204 10616 494210 10668
rect 82722 10548 82728 10600
rect 82780 10588 82786 10600
rect 197446 10588 197452 10600
rect 82780 10560 197452 10588
rect 82780 10548 82786 10560
rect 197446 10548 197452 10560
rect 197504 10548 197510 10600
rect 340690 10548 340696 10600
rect 340748 10588 340754 10600
rect 496814 10588 496820 10600
rect 340748 10560 496820 10588
rect 340748 10548 340754 10560
rect 496814 10548 496820 10560
rect 496872 10548 496878 10600
rect 78582 10480 78588 10532
rect 78640 10520 78646 10532
rect 195974 10520 195980 10532
rect 78640 10492 195980 10520
rect 78640 10480 78646 10492
rect 195974 10480 195980 10492
rect 196032 10480 196038 10532
rect 342162 10480 342168 10532
rect 342220 10520 342226 10532
rect 500954 10520 500960 10532
rect 342220 10492 500960 10520
rect 342220 10480 342226 10492
rect 500954 10480 500960 10492
rect 501012 10480 501018 10532
rect 74442 10412 74448 10464
rect 74500 10452 74506 10464
rect 194870 10452 194876 10464
rect 74500 10424 194876 10452
rect 74500 10412 74506 10424
rect 194870 10412 194876 10424
rect 194928 10412 194934 10464
rect 343542 10412 343548 10464
rect 343600 10452 343606 10464
rect 503714 10452 503720 10464
rect 343600 10424 503720 10452
rect 343600 10412 343606 10424
rect 503714 10412 503720 10424
rect 503772 10412 503778 10464
rect 71682 10344 71688 10396
rect 71740 10384 71746 10396
rect 193306 10384 193312 10396
rect 71740 10356 193312 10384
rect 71740 10344 71746 10356
rect 193306 10344 193312 10356
rect 193364 10344 193370 10396
rect 344830 10344 344836 10396
rect 344888 10384 344894 10396
rect 507854 10384 507860 10396
rect 344888 10356 507860 10384
rect 344888 10344 344894 10356
rect 507854 10344 507860 10356
rect 507912 10344 507918 10396
rect 28902 10276 28908 10328
rect 28960 10316 28966 10328
rect 179598 10316 179604 10328
rect 28960 10288 179604 10316
rect 28960 10276 28966 10288
rect 179598 10276 179604 10288
rect 179656 10276 179662 10328
rect 347498 10276 347504 10328
rect 347556 10316 347562 10328
rect 513374 10316 513380 10328
rect 347556 10288 513380 10316
rect 347556 10276 347562 10288
rect 513374 10276 513380 10288
rect 513432 10276 513438 10328
rect 107562 10208 107568 10260
rect 107620 10248 107626 10260
rect 205726 10248 205732 10260
rect 107620 10220 205732 10248
rect 107620 10208 107626 10220
rect 205726 10208 205732 10220
rect 205784 10208 205790 10260
rect 306190 10208 306196 10260
rect 306248 10248 306254 10260
rect 393314 10248 393320 10260
rect 306248 10220 393320 10248
rect 306248 10208 306254 10220
rect 393314 10208 393320 10220
rect 393372 10208 393378 10260
rect 110322 10140 110328 10192
rect 110380 10180 110386 10192
rect 207106 10180 207112 10192
rect 110380 10152 207112 10180
rect 110380 10140 110386 10152
rect 207106 10140 207112 10152
rect 207164 10140 207170 10192
rect 304902 10140 304908 10192
rect 304960 10180 304966 10192
rect 390646 10180 390652 10192
rect 304960 10152 390652 10180
rect 304960 10140 304966 10152
rect 390646 10140 390652 10152
rect 390704 10140 390710 10192
rect 114462 10072 114468 10124
rect 114520 10112 114526 10124
rect 208486 10112 208492 10124
rect 114520 10084 208492 10112
rect 114520 10072 114526 10084
rect 208486 10072 208492 10084
rect 208544 10072 208550 10124
rect 303522 10072 303528 10124
rect 303580 10112 303586 10124
rect 386414 10112 386420 10124
rect 303580 10084 386420 10112
rect 303580 10072 303586 10084
rect 386414 10072 386420 10084
rect 386472 10072 386478 10124
rect 150342 10004 150348 10056
rect 150400 10044 150406 10056
rect 221090 10044 221096 10056
rect 150400 10016 221096 10044
rect 150400 10004 150406 10016
rect 221090 10004 221096 10016
rect 221148 10004 221154 10056
rect 302142 10004 302148 10056
rect 302200 10044 302206 10056
rect 382366 10044 382372 10056
rect 302200 10016 382372 10044
rect 302200 10004 302206 10016
rect 382366 10004 382372 10016
rect 382424 10004 382430 10056
rect 153102 9936 153108 9988
rect 153160 9976 153166 9988
rect 222378 9976 222384 9988
rect 153160 9948 222384 9976
rect 153160 9936 153166 9948
rect 222378 9936 222384 9948
rect 222436 9936 222442 9988
rect 300762 9936 300768 9988
rect 300820 9976 300826 9988
rect 379514 9976 379520 9988
rect 300820 9948 379520 9976
rect 300820 9936 300826 9948
rect 379514 9936 379520 9948
rect 379572 9936 379578 9988
rect 157242 9868 157248 9920
rect 157300 9908 157306 9920
rect 223850 9908 223856 9920
rect 157300 9880 223856 9908
rect 157300 9868 157306 9880
rect 223850 9868 223856 9880
rect 223908 9868 223914 9920
rect 299382 9868 299388 9920
rect 299440 9908 299446 9920
rect 375374 9908 375380 9920
rect 299440 9880 375380 9908
rect 299440 9868 299446 9880
rect 375374 9868 375380 9880
rect 375432 9868 375438 9920
rect 283929 9775 283987 9781
rect 283929 9741 283941 9775
rect 283975 9772 283987 9775
rect 284018 9772 284024 9784
rect 283975 9744 284024 9772
rect 283975 9741 283987 9744
rect 283929 9735 283987 9741
rect 284018 9732 284024 9744
rect 284076 9732 284082 9784
rect 189258 9664 189264 9716
rect 189316 9704 189322 9716
rect 189534 9704 189540 9716
rect 189316 9676 189540 9704
rect 189316 9664 189322 9676
rect 189534 9664 189540 9676
rect 189592 9664 189598 9716
rect 192110 9704 192116 9716
rect 192071 9676 192116 9704
rect 192110 9664 192116 9676
rect 192168 9664 192174 9716
rect 212258 9704 212264 9716
rect 212219 9676 212264 9704
rect 212258 9664 212264 9676
rect 212316 9664 212322 9716
rect 214282 9704 214288 9716
rect 214243 9676 214288 9704
rect 214282 9664 214288 9676
rect 214340 9664 214346 9716
rect 277121 9707 277179 9713
rect 277121 9673 277133 9707
rect 277167 9704 277179 9707
rect 277210 9704 277216 9716
rect 277167 9676 277216 9704
rect 277167 9673 277179 9676
rect 277121 9667 277179 9673
rect 277210 9664 277216 9676
rect 277268 9664 277274 9716
rect 291838 9704 291844 9716
rect 291799 9676 291844 9704
rect 291838 9664 291844 9676
rect 291896 9664 291902 9716
rect 328178 9704 328184 9716
rect 328139 9676 328184 9704
rect 328178 9664 328184 9676
rect 328236 9664 328242 9716
rect 329466 9704 329472 9716
rect 329427 9676 329472 9704
rect 329466 9664 329472 9676
rect 329524 9664 329530 9716
rect 362494 9704 362500 9716
rect 362455 9676 362500 9704
rect 362494 9664 362500 9676
rect 362552 9664 362558 9716
rect 138474 9596 138480 9648
rect 138532 9636 138538 9648
rect 138532 9608 216904 9636
rect 138532 9596 138538 9608
rect 216876 9580 216904 9608
rect 216950 9596 216956 9648
rect 217008 9596 217014 9648
rect 317046 9596 317052 9648
rect 317104 9636 317110 9648
rect 427538 9636 427544 9648
rect 317104 9608 427544 9636
rect 317104 9596 317110 9608
rect 427538 9596 427544 9608
rect 427596 9596 427602 9648
rect 137278 9528 137284 9580
rect 137336 9568 137342 9580
rect 137336 9540 215524 9568
rect 137336 9528 137342 9540
rect 134886 9460 134892 9512
rect 134944 9500 134950 9512
rect 215386 9500 215392 9512
rect 134944 9472 215392 9500
rect 134944 9460 134950 9472
rect 215386 9460 215392 9472
rect 215444 9460 215450 9512
rect 215496 9500 215524 9540
rect 216858 9528 216864 9580
rect 216916 9528 216922 9580
rect 216968 9500 216996 9596
rect 318334 9528 318340 9580
rect 318392 9568 318398 9580
rect 431126 9568 431132 9580
rect 318392 9540 431132 9568
rect 318392 9528 318398 9540
rect 431126 9528 431132 9540
rect 431184 9528 431190 9580
rect 215496 9472 216996 9500
rect 319990 9460 319996 9512
rect 320048 9500 320054 9512
rect 434622 9500 434628 9512
rect 320048 9472 434628 9500
rect 320048 9460 320054 9472
rect 434622 9460 434628 9472
rect 434680 9460 434686 9512
rect 131390 9392 131396 9444
rect 131448 9432 131454 9444
rect 214006 9432 214012 9444
rect 131448 9404 214012 9432
rect 131448 9392 131454 9404
rect 214006 9392 214012 9404
rect 214064 9392 214070 9444
rect 321370 9392 321376 9444
rect 321428 9432 321434 9444
rect 438210 9432 438216 9444
rect 321428 9404 438216 9432
rect 321428 9392 321434 9404
rect 438210 9392 438216 9404
rect 438268 9392 438274 9444
rect 133782 9324 133788 9376
rect 133840 9364 133846 9376
rect 215570 9364 215576 9376
rect 133840 9336 215576 9364
rect 133840 9324 133846 9336
rect 215570 9324 215576 9336
rect 215628 9324 215634 9376
rect 322658 9324 322664 9376
rect 322716 9364 322722 9376
rect 441798 9364 441804 9376
rect 322716 9336 441804 9364
rect 322716 9324 322722 9336
rect 441798 9324 441804 9336
rect 441856 9324 441862 9376
rect 130194 9256 130200 9308
rect 130252 9296 130258 9308
rect 214282 9296 214288 9308
rect 130252 9268 214288 9296
rect 130252 9256 130258 9268
rect 214282 9256 214288 9268
rect 214340 9256 214346 9308
rect 322750 9256 322756 9308
rect 322808 9296 322814 9308
rect 445386 9296 445392 9308
rect 322808 9268 445392 9296
rect 322808 9256 322814 9268
rect 445386 9256 445392 9268
rect 445444 9256 445450 9308
rect 126606 9188 126612 9240
rect 126664 9228 126670 9240
rect 212902 9228 212908 9240
rect 126664 9200 212908 9228
rect 126664 9188 126670 9200
rect 212902 9188 212908 9200
rect 212960 9188 212966 9240
rect 324130 9188 324136 9240
rect 324188 9228 324194 9240
rect 448974 9228 448980 9240
rect 324188 9200 448980 9228
rect 324188 9188 324194 9200
rect 448974 9188 448980 9200
rect 449032 9188 449038 9240
rect 67174 9120 67180 9172
rect 67232 9160 67238 9172
rect 192018 9160 192024 9172
rect 67232 9132 192024 9160
rect 67232 9120 67238 9132
rect 192018 9120 192024 9132
rect 192076 9120 192082 9172
rect 325510 9120 325516 9172
rect 325568 9160 325574 9172
rect 452470 9160 452476 9172
rect 325568 9132 452476 9160
rect 325568 9120 325574 9132
rect 452470 9120 452476 9132
rect 452528 9120 452534 9172
rect 23106 9052 23112 9104
rect 23164 9092 23170 9104
rect 177022 9092 177028 9104
rect 23164 9064 177028 9092
rect 23164 9052 23170 9064
rect 177022 9052 177028 9064
rect 177080 9052 177086 9104
rect 180150 9052 180156 9104
rect 180208 9092 180214 9104
rect 230934 9092 230940 9104
rect 180208 9064 230940 9092
rect 180208 9052 180214 9064
rect 230934 9052 230940 9064
rect 230992 9052 230998 9104
rect 326798 9052 326804 9104
rect 326856 9092 326862 9104
rect 456058 9092 456064 9104
rect 326856 9064 456064 9092
rect 326856 9052 326862 9064
rect 456058 9052 456064 9064
rect 456116 9052 456122 9104
rect 18322 8984 18328 9036
rect 18380 9024 18386 9036
rect 175366 9024 175372 9036
rect 18380 8996 175372 9024
rect 18380 8984 18386 8996
rect 175366 8984 175372 8996
rect 175424 8984 175430 9036
rect 177758 8984 177764 9036
rect 177816 9024 177822 9036
rect 230658 9024 230664 9036
rect 177816 8996 230664 9024
rect 177816 8984 177822 8996
rect 230658 8984 230664 8996
rect 230716 8984 230722 9036
rect 328178 8984 328184 9036
rect 328236 9024 328242 9036
rect 459646 9024 459652 9036
rect 328236 8996 459652 9024
rect 328236 8984 328242 8996
rect 459646 8984 459652 8996
rect 459704 8984 459710 9036
rect 13630 8916 13636 8968
rect 13688 8956 13694 8968
rect 173986 8956 173992 8968
rect 13688 8928 173992 8956
rect 13688 8916 13694 8928
rect 173986 8916 173992 8928
rect 174044 8916 174050 8968
rect 176562 8916 176568 8968
rect 176620 8956 176626 8968
rect 230566 8956 230572 8968
rect 176620 8928 230572 8956
rect 176620 8916 176626 8928
rect 230566 8916 230572 8928
rect 230624 8916 230630 8968
rect 329466 8916 329472 8968
rect 329524 8956 329530 8968
rect 463234 8956 463240 8968
rect 329524 8928 463240 8956
rect 329524 8916 329530 8928
rect 463234 8916 463240 8928
rect 463292 8916 463298 8968
rect 140866 8848 140872 8900
rect 140924 8888 140930 8900
rect 218146 8888 218152 8900
rect 140924 8860 218152 8888
rect 140924 8848 140930 8860
rect 218146 8848 218152 8860
rect 218204 8848 218210 8900
rect 315850 8848 315856 8900
rect 315908 8888 315914 8900
rect 423950 8888 423956 8900
rect 315908 8860 423956 8888
rect 315908 8848 315914 8860
rect 423950 8848 423956 8860
rect 424008 8848 424014 8900
rect 142062 8780 142068 8832
rect 142120 8820 142126 8832
rect 218238 8820 218244 8832
rect 142120 8792 218244 8820
rect 142120 8780 142126 8792
rect 218238 8780 218244 8792
rect 218296 8780 218302 8832
rect 314470 8780 314476 8832
rect 314528 8820 314534 8832
rect 420362 8820 420368 8832
rect 314528 8792 420368 8820
rect 314528 8780 314534 8792
rect 420362 8780 420368 8792
rect 420420 8780 420426 8832
rect 145650 8712 145656 8764
rect 145708 8752 145714 8764
rect 219618 8752 219624 8764
rect 145708 8724 219624 8752
rect 145708 8712 145714 8724
rect 219618 8712 219624 8724
rect 219676 8712 219682 8764
rect 313090 8712 313096 8764
rect 313148 8752 313154 8764
rect 416866 8752 416872 8764
rect 313148 8724 416872 8752
rect 313148 8712 313154 8724
rect 416866 8712 416872 8724
rect 416924 8712 416930 8764
rect 117130 8644 117136 8696
rect 117188 8684 117194 8696
rect 179966 8684 179972 8696
rect 117188 8656 179972 8684
rect 117188 8644 117194 8656
rect 179966 8644 179972 8656
rect 180024 8644 180030 8696
rect 311710 8644 311716 8696
rect 311768 8684 311774 8696
rect 413278 8684 413284 8696
rect 311768 8656 413284 8684
rect 311768 8644 311774 8656
rect 413278 8644 413284 8656
rect 413336 8644 413342 8696
rect 162302 8576 162308 8628
rect 162360 8616 162366 8628
rect 225230 8616 225236 8628
rect 162360 8588 225236 8616
rect 162360 8576 162366 8588
rect 225230 8576 225236 8588
rect 225288 8576 225294 8628
rect 311618 8576 311624 8628
rect 311676 8616 311682 8628
rect 409690 8616 409696 8628
rect 311676 8588 409696 8616
rect 311676 8576 311682 8588
rect 409690 8576 409696 8588
rect 409748 8576 409754 8628
rect 165890 8508 165896 8560
rect 165948 8548 165954 8560
rect 226610 8548 226616 8560
rect 165948 8520 226616 8548
rect 165948 8508 165954 8520
rect 226610 8508 226616 8520
rect 226668 8508 226674 8560
rect 310330 8508 310336 8560
rect 310388 8548 310394 8560
rect 406102 8548 406108 8560
rect 310388 8520 406108 8548
rect 310388 8508 310394 8520
rect 406102 8508 406108 8520
rect 406160 8508 406166 8560
rect 169386 8440 169392 8492
rect 169444 8480 169450 8492
rect 227990 8480 227996 8492
rect 169444 8452 227996 8480
rect 169444 8440 169450 8452
rect 227990 8440 227996 8452
rect 228048 8440 228054 8492
rect 308950 8440 308956 8492
rect 309008 8480 309014 8492
rect 402514 8480 402520 8492
rect 309008 8452 402520 8480
rect 309008 8440 309014 8452
rect 402514 8440 402520 8452
rect 402572 8440 402578 8492
rect 172974 8372 172980 8424
rect 173032 8412 173038 8424
rect 229370 8412 229376 8424
rect 173032 8384 229376 8412
rect 173032 8372 173038 8384
rect 229370 8372 229376 8384
rect 229428 8372 229434 8424
rect 307662 8372 307668 8424
rect 307720 8412 307726 8424
rect 399018 8412 399024 8424
rect 307720 8384 399024 8412
rect 307720 8372 307726 8384
rect 399018 8372 399024 8384
rect 399076 8372 399082 8424
rect 181070 8304 181076 8356
rect 181128 8344 181134 8356
rect 181254 8344 181260 8356
rect 181128 8316 181260 8344
rect 181128 8304 181134 8316
rect 181254 8304 181260 8316
rect 181312 8304 181318 8356
rect 182174 8304 182180 8356
rect 182232 8344 182238 8356
rect 182450 8344 182456 8356
rect 182232 8316 182456 8344
rect 182232 8304 182238 8316
rect 182450 8304 182456 8316
rect 182508 8304 182514 8356
rect 283926 8344 283932 8356
rect 283887 8316 283932 8344
rect 283926 8304 283932 8316
rect 283984 8304 283990 8356
rect 306282 8304 306288 8356
rect 306340 8344 306346 8356
rect 395430 8344 395436 8356
rect 306340 8316 395436 8344
rect 306340 8304 306346 8316
rect 395430 8304 395436 8316
rect 395488 8304 395494 8356
rect 101582 8236 101588 8288
rect 101640 8276 101646 8288
rect 204530 8276 204536 8288
rect 101640 8248 204536 8276
rect 101640 8236 101646 8248
rect 204530 8236 204536 8248
rect 204588 8236 204594 8288
rect 355778 8236 355784 8288
rect 355836 8276 355842 8288
rect 541710 8276 541716 8288
rect 355836 8248 541716 8276
rect 355836 8236 355842 8248
rect 541710 8236 541716 8248
rect 541768 8236 541774 8288
rect 98086 8168 98092 8220
rect 98144 8208 98150 8220
rect 203150 8208 203156 8220
rect 98144 8180 203156 8208
rect 98144 8168 98150 8180
rect 203150 8168 203156 8180
rect 203208 8168 203214 8220
rect 357250 8168 357256 8220
rect 357308 8208 357314 8220
rect 545298 8208 545304 8220
rect 357308 8180 545304 8208
rect 357308 8168 357314 8180
rect 545298 8168 545304 8180
rect 545356 8168 545362 8220
rect 94498 8100 94504 8152
rect 94556 8140 94562 8152
rect 201862 8140 201868 8152
rect 94556 8112 201868 8140
rect 94556 8100 94562 8112
rect 201862 8100 201868 8112
rect 201920 8100 201926 8152
rect 358630 8100 358636 8152
rect 358688 8140 358694 8152
rect 548886 8140 548892 8152
rect 358688 8112 548892 8140
rect 358688 8100 358694 8112
rect 548886 8100 548892 8112
rect 548944 8100 548950 8152
rect 90910 8032 90916 8084
rect 90968 8072 90974 8084
rect 200390 8072 200396 8084
rect 90968 8044 200396 8072
rect 90968 8032 90974 8044
rect 200390 8032 200396 8044
rect 200448 8032 200454 8084
rect 289265 8075 289323 8081
rect 289265 8041 289277 8075
rect 289311 8072 289323 8075
rect 346670 8072 346676 8084
rect 289311 8044 346676 8072
rect 289311 8041 289323 8044
rect 289265 8035 289323 8041
rect 346670 8032 346676 8044
rect 346728 8032 346734 8084
rect 359918 8032 359924 8084
rect 359976 8072 359982 8084
rect 552382 8072 552388 8084
rect 359976 8044 552388 8072
rect 359976 8032 359982 8044
rect 552382 8032 552388 8044
rect 552440 8032 552446 8084
rect 87322 7964 87328 8016
rect 87380 8004 87386 8016
rect 198826 8004 198832 8016
rect 87380 7976 198832 8004
rect 87380 7964 87386 7976
rect 198826 7964 198832 7976
rect 198884 7964 198890 8016
rect 289538 7964 289544 8016
rect 289596 8004 289602 8016
rect 349062 8004 349068 8016
rect 289596 7976 349068 8004
rect 289596 7964 289602 7976
rect 349062 7964 349068 7976
rect 349120 7964 349126 8016
rect 361298 7964 361304 8016
rect 361356 8004 361362 8016
rect 555970 8004 555976 8016
rect 361356 7976 555976 8004
rect 361356 7964 361362 7976
rect 555970 7964 555976 7976
rect 556028 7964 556034 8016
rect 83826 7896 83832 7948
rect 83884 7936 83890 7948
rect 198734 7936 198740 7948
rect 83884 7908 198740 7936
rect 83884 7896 83890 7908
rect 198734 7896 198740 7908
rect 198792 7896 198798 7948
rect 290918 7896 290924 7948
rect 290976 7936 290982 7948
rect 352558 7936 352564 7948
rect 290976 7908 352564 7936
rect 290976 7896 290982 7908
rect 352558 7896 352564 7908
rect 352616 7896 352622 7948
rect 363598 7896 363604 7948
rect 363656 7936 363662 7948
rect 559558 7936 559564 7948
rect 363656 7908 559564 7936
rect 363656 7896 363662 7908
rect 559558 7896 559564 7908
rect 559616 7896 559622 7948
rect 80238 7828 80244 7880
rect 80296 7868 80302 7880
rect 197538 7868 197544 7880
rect 80296 7840 197544 7868
rect 80296 7828 80302 7840
rect 197538 7828 197544 7840
rect 197596 7828 197602 7880
rect 292298 7828 292304 7880
rect 292356 7868 292362 7880
rect 356146 7868 356152 7880
rect 292356 7840 356152 7868
rect 292356 7828 292362 7840
rect 356146 7828 356152 7840
rect 356204 7828 356210 7880
rect 364150 7828 364156 7880
rect 364208 7868 364214 7880
rect 563146 7868 563152 7880
rect 364208 7840 563152 7868
rect 364208 7828 364214 7840
rect 563146 7828 563152 7840
rect 563204 7828 563210 7880
rect 76650 7760 76656 7812
rect 76708 7800 76714 7812
rect 196158 7800 196164 7812
rect 76708 7772 196164 7800
rect 76708 7760 76714 7772
rect 196158 7760 196164 7772
rect 196216 7760 196222 7812
rect 293678 7760 293684 7812
rect 293736 7800 293742 7812
rect 359734 7800 359740 7812
rect 293736 7772 359740 7800
rect 293736 7760 293742 7772
rect 359734 7760 359740 7772
rect 359792 7760 359798 7812
rect 365438 7760 365444 7812
rect 365496 7800 365502 7812
rect 566734 7800 566740 7812
rect 365496 7772 566740 7800
rect 365496 7760 365502 7772
rect 566734 7760 566740 7772
rect 566792 7760 566798 7812
rect 63586 7692 63592 7744
rect 63644 7732 63650 7744
rect 191926 7732 191932 7744
rect 63644 7704 191932 7732
rect 63644 7692 63650 7704
rect 191926 7692 191932 7704
rect 191984 7692 191990 7744
rect 294966 7692 294972 7744
rect 295024 7732 295030 7744
rect 363322 7732 363328 7744
rect 295024 7704 363328 7732
rect 295024 7692 295030 7704
rect 363322 7692 363328 7704
rect 363380 7692 363386 7744
rect 366818 7692 366824 7744
rect 366876 7732 366882 7744
rect 570230 7732 570236 7744
rect 366876 7704 570236 7732
rect 366876 7692 366882 7704
rect 570230 7692 570236 7704
rect 570288 7692 570294 7744
rect 59998 7624 60004 7676
rect 60056 7664 60062 7676
rect 190546 7664 190552 7676
rect 60056 7636 190552 7664
rect 60056 7624 60062 7636
rect 190546 7624 190552 7636
rect 190604 7624 190610 7676
rect 296530 7624 296536 7676
rect 296588 7664 296594 7676
rect 366910 7664 366916 7676
rect 296588 7636 366916 7664
rect 296588 7624 296594 7636
rect 366910 7624 366916 7636
rect 366968 7624 366974 7676
rect 367002 7624 367008 7676
rect 367060 7664 367066 7676
rect 573818 7664 573824 7676
rect 367060 7636 573824 7664
rect 367060 7624 367066 7636
rect 573818 7624 573824 7636
rect 573876 7624 573882 7676
rect 56410 7556 56416 7608
rect 56468 7596 56474 7608
rect 189166 7596 189172 7608
rect 56468 7568 189172 7596
rect 56468 7556 56474 7568
rect 189166 7556 189172 7568
rect 189224 7556 189230 7608
rect 295150 7556 295156 7608
rect 295208 7596 295214 7608
rect 364518 7596 364524 7608
rect 295208 7568 364524 7596
rect 295208 7556 295214 7568
rect 364518 7556 364524 7568
rect 364576 7556 364582 7608
rect 368198 7556 368204 7608
rect 368256 7596 368262 7608
rect 577406 7596 577412 7608
rect 368256 7568 577412 7596
rect 368256 7556 368262 7568
rect 577406 7556 577412 7568
rect 577464 7556 577470 7608
rect 105170 7488 105176 7540
rect 105228 7528 105234 7540
rect 205818 7528 205824 7540
rect 105228 7500 205824 7528
rect 105228 7488 105234 7500
rect 205818 7488 205824 7500
rect 205876 7488 205882 7540
rect 355870 7488 355876 7540
rect 355928 7528 355934 7540
rect 538122 7528 538128 7540
rect 355928 7500 538128 7528
rect 355928 7488 355934 7500
rect 538122 7488 538128 7500
rect 538180 7488 538186 7540
rect 108758 7420 108764 7472
rect 108816 7460 108822 7472
rect 207198 7460 207204 7472
rect 108816 7432 207204 7460
rect 108816 7420 108822 7432
rect 207198 7420 207204 7432
rect 207256 7420 207262 7472
rect 354490 7420 354496 7472
rect 354548 7460 354554 7472
rect 534534 7460 534540 7472
rect 354548 7432 534540 7460
rect 354548 7420 354554 7432
rect 534534 7420 534540 7432
rect 534592 7420 534598 7472
rect 112346 7352 112352 7404
rect 112404 7392 112410 7404
rect 208578 7392 208584 7404
rect 112404 7364 208584 7392
rect 112404 7352 112410 7364
rect 208578 7352 208584 7364
rect 208636 7352 208642 7404
rect 353110 7352 353116 7404
rect 353168 7392 353174 7404
rect 531038 7392 531044 7404
rect 353168 7364 531044 7392
rect 353168 7352 353174 7364
rect 531038 7352 531044 7364
rect 531096 7352 531102 7404
rect 115934 7284 115940 7336
rect 115992 7324 115998 7336
rect 209774 7324 209780 7336
rect 115992 7296 209780 7324
rect 115992 7284 115998 7296
rect 209774 7284 209780 7296
rect 209832 7284 209838 7336
rect 351638 7284 351644 7336
rect 351696 7324 351702 7336
rect 527450 7324 527456 7336
rect 351696 7296 527456 7324
rect 351696 7284 351702 7296
rect 527450 7284 527456 7296
rect 527508 7284 527514 7336
rect 119430 7216 119436 7268
rect 119488 7256 119494 7268
rect 209866 7256 209872 7268
rect 119488 7228 209872 7256
rect 119488 7216 119494 7228
rect 209866 7216 209872 7228
rect 209924 7216 209930 7268
rect 350350 7216 350356 7268
rect 350408 7256 350414 7268
rect 523862 7256 523868 7268
rect 350408 7228 523868 7256
rect 350408 7216 350414 7228
rect 523862 7216 523868 7228
rect 523920 7216 523926 7268
rect 123018 7148 123024 7200
rect 123076 7188 123082 7200
rect 211338 7188 211344 7200
rect 123076 7160 211344 7188
rect 123076 7148 123082 7160
rect 211338 7148 211344 7160
rect 211396 7148 211402 7200
rect 348786 7148 348792 7200
rect 348844 7188 348850 7200
rect 520366 7188 520372 7200
rect 348844 7160 520372 7188
rect 348844 7148 348850 7160
rect 520366 7148 520372 7160
rect 520424 7148 520430 7200
rect 153930 7080 153936 7132
rect 153988 7120 153994 7132
rect 222286 7120 222292 7132
rect 153988 7092 222292 7120
rect 153988 7080 153994 7092
rect 222286 7080 222292 7092
rect 222344 7080 222350 7132
rect 347590 7080 347596 7132
rect 347648 7120 347654 7132
rect 516778 7120 516784 7132
rect 347648 7092 516784 7120
rect 347648 7080 347654 7092
rect 516778 7080 516784 7092
rect 516836 7080 516842 7132
rect 157518 7012 157524 7064
rect 157576 7052 157582 7064
rect 223758 7052 223764 7064
rect 157576 7024 223764 7052
rect 157576 7012 157582 7024
rect 223758 7012 223764 7024
rect 223816 7012 223822 7064
rect 346210 7012 346216 7064
rect 346268 7052 346274 7064
rect 513190 7052 513196 7064
rect 346268 7024 513196 7052
rect 346268 7012 346274 7024
rect 513190 7012 513196 7024
rect 513248 7012 513254 7064
rect 161106 6944 161112 6996
rect 161164 6984 161170 6996
rect 225046 6984 225052 6996
rect 161164 6956 225052 6984
rect 161164 6944 161170 6956
rect 225046 6944 225052 6956
rect 225104 6944 225110 6996
rect 344922 6944 344928 6996
rect 344980 6984 344986 6996
rect 509602 6984 509608 6996
rect 344980 6956 509608 6984
rect 344980 6944 344986 6956
rect 509602 6944 509608 6956
rect 509660 6944 509666 6996
rect 128998 6808 129004 6860
rect 129056 6848 129062 6860
rect 213914 6848 213920 6860
rect 129056 6820 213920 6848
rect 129056 6808 129062 6820
rect 213914 6808 213920 6820
rect 213972 6808 213978 6860
rect 320082 6808 320088 6860
rect 320140 6848 320146 6860
rect 437014 6848 437020 6860
rect 320140 6820 437020 6848
rect 320140 6808 320146 6820
rect 437014 6808 437020 6820
rect 437072 6808 437078 6860
rect 73062 6740 73068 6792
rect 73120 6780 73126 6792
rect 194778 6780 194784 6792
rect 73120 6752 194784 6780
rect 73120 6740 73126 6752
rect 194778 6740 194784 6752
rect 194836 6740 194842 6792
rect 321462 6740 321468 6792
rect 321520 6780 321526 6792
rect 440602 6780 440608 6792
rect 321520 6752 440608 6780
rect 321520 6740 321526 6752
rect 440602 6740 440608 6752
rect 440660 6740 440666 6792
rect 49326 6672 49332 6724
rect 49384 6712 49390 6724
rect 186406 6712 186412 6724
rect 49384 6684 186412 6712
rect 49384 6672 49390 6684
rect 186406 6672 186412 6684
rect 186464 6672 186470 6724
rect 322842 6672 322848 6724
rect 322900 6712 322906 6724
rect 444190 6712 444196 6724
rect 322900 6684 444196 6712
rect 322900 6672 322906 6684
rect 444190 6672 444196 6684
rect 444248 6672 444254 6724
rect 44542 6604 44548 6656
rect 44600 6644 44606 6656
rect 185118 6644 185124 6656
rect 44600 6616 185124 6644
rect 44600 6604 44606 6616
rect 185118 6604 185124 6616
rect 185176 6604 185182 6656
rect 324222 6604 324228 6656
rect 324280 6644 324286 6656
rect 447778 6644 447784 6656
rect 324280 6616 447784 6644
rect 324280 6604 324286 6616
rect 447778 6604 447784 6616
rect 447836 6604 447842 6656
rect 40954 6536 40960 6588
rect 41012 6576 41018 6588
rect 183738 6576 183744 6588
rect 41012 6548 183744 6576
rect 41012 6536 41018 6548
rect 183738 6536 183744 6548
rect 183796 6536 183802 6588
rect 325602 6536 325608 6588
rect 325660 6576 325666 6588
rect 451274 6576 451280 6588
rect 325660 6548 451280 6576
rect 325660 6536 325666 6548
rect 451274 6536 451280 6548
rect 451332 6536 451338 6588
rect 37366 6468 37372 6520
rect 37424 6508 37430 6520
rect 182266 6508 182272 6520
rect 37424 6480 182272 6508
rect 37424 6468 37430 6480
rect 182266 6468 182272 6480
rect 182324 6468 182330 6520
rect 326982 6468 326988 6520
rect 327040 6508 327046 6520
rect 454862 6508 454868 6520
rect 327040 6480 454868 6508
rect 327040 6468 327046 6480
rect 454862 6468 454868 6480
rect 454920 6468 454926 6520
rect 33870 6400 33876 6452
rect 33928 6440 33934 6452
rect 180886 6440 180892 6452
rect 33928 6412 180892 6440
rect 33928 6400 33934 6412
rect 180886 6400 180892 6412
rect 180944 6400 180950 6452
rect 186038 6400 186044 6452
rect 186096 6440 186102 6452
rect 233510 6440 233516 6452
rect 186096 6412 233516 6440
rect 186096 6400 186102 6412
rect 233510 6400 233516 6412
rect 233568 6400 233574 6452
rect 328362 6400 328368 6452
rect 328420 6440 328426 6452
rect 458450 6440 458456 6452
rect 328420 6412 458456 6440
rect 328420 6400 328426 6412
rect 458450 6400 458456 6412
rect 458508 6400 458514 6452
rect 30282 6332 30288 6384
rect 30340 6372 30346 6384
rect 179506 6372 179512 6384
rect 30340 6344 179512 6372
rect 30340 6332 30346 6344
rect 179506 6332 179512 6344
rect 179564 6332 179570 6384
rect 182542 6332 182548 6384
rect 182600 6372 182606 6384
rect 232130 6372 232136 6384
rect 182600 6344 232136 6372
rect 182600 6332 182606 6344
rect 232130 6332 232136 6344
rect 232188 6332 232194 6384
rect 329650 6332 329656 6384
rect 329708 6372 329714 6384
rect 462038 6372 462044 6384
rect 329708 6344 462044 6372
rect 329708 6332 329714 6344
rect 462038 6332 462044 6344
rect 462096 6332 462102 6384
rect 26694 6264 26700 6316
rect 26752 6304 26758 6316
rect 178126 6304 178132 6316
rect 26752 6276 178132 6304
rect 26752 6264 26758 6276
rect 178126 6264 178132 6276
rect 178184 6264 178190 6316
rect 178954 6264 178960 6316
rect 179012 6304 179018 6316
rect 230474 6304 230480 6316
rect 179012 6276 230480 6304
rect 179012 6264 179018 6276
rect 230474 6264 230480 6276
rect 230532 6264 230538 6316
rect 329742 6264 329748 6316
rect 329800 6304 329806 6316
rect 465626 6304 465632 6316
rect 329800 6276 465632 6304
rect 329800 6264 329806 6276
rect 465626 6264 465632 6276
rect 465684 6264 465690 6316
rect 8846 6196 8852 6248
rect 8904 6236 8910 6248
rect 172790 6236 172796 6248
rect 8904 6208 172796 6236
rect 8904 6196 8910 6208
rect 172790 6196 172796 6208
rect 172848 6196 172854 6248
rect 175366 6196 175372 6248
rect 175424 6236 175430 6248
rect 229186 6236 229192 6248
rect 175424 6208 229192 6236
rect 175424 6196 175430 6208
rect 229186 6196 229192 6208
rect 229244 6196 229250 6248
rect 331122 6196 331128 6248
rect 331180 6236 331186 6248
rect 469122 6236 469128 6248
rect 331180 6208 469128 6236
rect 331180 6196 331186 6208
rect 469122 6196 469128 6208
rect 469180 6196 469186 6248
rect 4062 6128 4068 6180
rect 4120 6168 4126 6180
rect 171226 6168 171232 6180
rect 4120 6140 171232 6168
rect 4120 6128 4126 6140
rect 171226 6128 171232 6140
rect 171284 6128 171290 6180
rect 171778 6128 171784 6180
rect 171836 6168 171842 6180
rect 227898 6168 227904 6180
rect 171836 6140 227904 6168
rect 171836 6128 171842 6140
rect 227898 6128 227904 6140
rect 227956 6128 227962 6180
rect 332502 6128 332508 6180
rect 332560 6168 332566 6180
rect 472710 6168 472716 6180
rect 332560 6140 472716 6168
rect 332560 6128 332566 6140
rect 472710 6128 472716 6140
rect 472768 6128 472774 6180
rect 132586 6060 132592 6112
rect 132644 6100 132650 6112
rect 215294 6100 215300 6112
rect 132644 6072 215300 6100
rect 132644 6060 132650 6072
rect 215294 6060 215300 6072
rect 215352 6060 215358 6112
rect 318702 6060 318708 6112
rect 318760 6100 318766 6112
rect 433518 6100 433524 6112
rect 318760 6072 433524 6100
rect 318760 6060 318766 6072
rect 433518 6060 433524 6072
rect 433576 6060 433582 6112
rect 136082 5992 136088 6044
rect 136140 6032 136146 6044
rect 216766 6032 216772 6044
rect 136140 6004 216772 6032
rect 136140 5992 136146 6004
rect 216766 5992 216772 6004
rect 216824 5992 216830 6044
rect 318610 5992 318616 6044
rect 318668 6032 318674 6044
rect 429930 6032 429936 6044
rect 318668 6004 429936 6032
rect 318668 5992 318674 6004
rect 429930 5992 429936 6004
rect 429988 5992 429994 6044
rect 139670 5924 139676 5976
rect 139728 5964 139734 5976
rect 217134 5964 217140 5976
rect 139728 5936 217140 5964
rect 139728 5924 139734 5936
rect 217134 5924 217140 5936
rect 217192 5924 217198 5976
rect 317322 5924 317328 5976
rect 317380 5964 317386 5976
rect 426342 5964 426348 5976
rect 317380 5936 426348 5964
rect 317380 5924 317386 5936
rect 426342 5924 426348 5936
rect 426400 5924 426406 5976
rect 143258 5856 143264 5908
rect 143316 5896 143322 5908
rect 218054 5896 218060 5908
rect 143316 5868 218060 5896
rect 143316 5856 143322 5868
rect 218054 5856 218060 5868
rect 218112 5856 218118 5908
rect 315942 5856 315948 5908
rect 316000 5896 316006 5908
rect 422754 5896 422760 5908
rect 316000 5868 422760 5896
rect 316000 5856 316006 5868
rect 422754 5856 422760 5868
rect 422812 5856 422818 5908
rect 146846 5788 146852 5840
rect 146904 5828 146910 5840
rect 219802 5828 219808 5840
rect 146904 5800 219808 5828
rect 146904 5788 146910 5800
rect 219802 5788 219808 5800
rect 219860 5788 219866 5840
rect 314562 5788 314568 5840
rect 314620 5828 314626 5840
rect 419166 5828 419172 5840
rect 314620 5800 419172 5828
rect 314620 5788 314626 5800
rect 419166 5788 419172 5800
rect 419224 5788 419230 5840
rect 150434 5720 150440 5772
rect 150492 5760 150498 5772
rect 220998 5760 221004 5772
rect 150492 5732 221004 5760
rect 150492 5720 150498 5732
rect 220998 5720 221004 5732
rect 221056 5720 221062 5772
rect 313182 5720 313188 5772
rect 313240 5760 313246 5772
rect 415670 5760 415676 5772
rect 313240 5732 415676 5760
rect 313240 5720 313246 5732
rect 415670 5720 415676 5732
rect 415728 5720 415734 5772
rect 159910 5652 159916 5704
rect 159968 5692 159974 5704
rect 224034 5692 224040 5704
rect 159968 5664 224040 5692
rect 159968 5652 159974 5664
rect 224034 5652 224040 5664
rect 224092 5652 224098 5704
rect 311802 5652 311808 5704
rect 311860 5692 311866 5704
rect 412082 5692 412088 5704
rect 311860 5664 412088 5692
rect 311860 5652 311866 5664
rect 412082 5652 412088 5664
rect 412140 5652 412146 5704
rect 164694 5584 164700 5636
rect 164752 5624 164758 5636
rect 226426 5624 226432 5636
rect 164752 5596 226432 5624
rect 164752 5584 164758 5596
rect 226426 5584 226432 5596
rect 226484 5584 226490 5636
rect 310422 5584 310428 5636
rect 310480 5624 310486 5636
rect 408494 5624 408500 5636
rect 310480 5596 408500 5624
rect 310480 5584 310486 5596
rect 408494 5584 408500 5596
rect 408552 5584 408558 5636
rect 168190 5516 168196 5568
rect 168248 5556 168254 5568
rect 227806 5556 227812 5568
rect 168248 5528 227812 5556
rect 168248 5516 168254 5528
rect 227806 5516 227812 5528
rect 227864 5516 227870 5568
rect 309042 5516 309048 5568
rect 309100 5556 309106 5568
rect 404906 5556 404912 5568
rect 309100 5528 404912 5556
rect 309100 5516 309106 5528
rect 404906 5516 404912 5528
rect 404964 5516 404970 5568
rect 65978 5448 65984 5500
rect 66036 5488 66042 5500
rect 192110 5488 192116 5500
rect 66036 5460 192116 5488
rect 66036 5448 66042 5460
rect 192110 5448 192116 5460
rect 192168 5448 192174 5500
rect 288250 5448 288256 5500
rect 288308 5488 288314 5500
rect 341886 5488 341892 5500
rect 288308 5460 341892 5488
rect 288308 5448 288314 5460
rect 341886 5448 341892 5460
rect 341944 5448 341950 5500
rect 357342 5448 357348 5500
rect 357400 5488 357406 5500
rect 544102 5488 544108 5500
rect 357400 5460 544108 5488
rect 357400 5448 357406 5460
rect 544102 5448 544108 5460
rect 544160 5448 544166 5500
rect 62390 5380 62396 5432
rect 62448 5420 62454 5432
rect 190638 5420 190644 5432
rect 62448 5392 190644 5420
rect 62448 5380 62454 5392
rect 190638 5380 190644 5392
rect 190696 5380 190702 5432
rect 286778 5380 286784 5432
rect 286836 5420 286842 5432
rect 340690 5420 340696 5432
rect 286836 5392 340696 5420
rect 286836 5380 286842 5392
rect 340690 5380 340696 5392
rect 340748 5380 340754 5432
rect 358722 5380 358728 5432
rect 358780 5420 358786 5432
rect 547690 5420 547696 5432
rect 358780 5392 547696 5420
rect 358780 5380 358786 5392
rect 547690 5380 547696 5392
rect 547748 5380 547754 5432
rect 58802 5312 58808 5364
rect 58860 5352 58866 5364
rect 189350 5352 189356 5364
rect 58860 5324 189356 5352
rect 58860 5312 58866 5324
rect 189350 5312 189356 5324
rect 189408 5312 189414 5364
rect 208670 5312 208676 5364
rect 208728 5352 208734 5364
rect 241698 5352 241704 5364
rect 208728 5324 241704 5352
rect 208728 5312 208734 5324
rect 241698 5312 241704 5324
rect 241756 5312 241762 5364
rect 289630 5312 289636 5364
rect 289688 5352 289694 5364
rect 345474 5352 345480 5364
rect 289688 5324 345480 5352
rect 289688 5312 289694 5324
rect 345474 5312 345480 5324
rect 345532 5312 345538 5364
rect 360010 5312 360016 5364
rect 360068 5352 360074 5364
rect 551186 5352 551192 5364
rect 360068 5324 551192 5352
rect 360068 5312 360074 5324
rect 551186 5312 551192 5324
rect 551244 5312 551250 5364
rect 55214 5244 55220 5296
rect 55272 5284 55278 5296
rect 187970 5284 187976 5296
rect 55272 5256 187976 5284
rect 55272 5244 55278 5256
rect 187970 5244 187976 5256
rect 188028 5244 188034 5296
rect 205082 5244 205088 5296
rect 205140 5284 205146 5296
rect 240318 5284 240324 5296
rect 205140 5256 240324 5284
rect 205140 5244 205146 5256
rect 240318 5244 240324 5256
rect 240376 5244 240382 5296
rect 288158 5244 288164 5296
rect 288216 5284 288222 5296
rect 344278 5284 344284 5296
rect 288216 5256 344284 5284
rect 288216 5244 288222 5256
rect 344278 5244 344284 5256
rect 344336 5244 344342 5296
rect 361482 5244 361488 5296
rect 361540 5284 361546 5296
rect 554774 5284 554780 5296
rect 361540 5256 554780 5284
rect 361540 5244 361546 5256
rect 554774 5244 554780 5256
rect 554832 5244 554838 5296
rect 51626 5176 51632 5228
rect 51684 5216 51690 5228
rect 187786 5216 187792 5228
rect 51684 5188 187792 5216
rect 51684 5176 51690 5188
rect 187786 5176 187792 5188
rect 187844 5176 187850 5228
rect 201494 5176 201500 5228
rect 201552 5216 201558 5228
rect 238938 5216 238944 5228
rect 201552 5188 238944 5216
rect 201552 5176 201558 5188
rect 238938 5176 238944 5188
rect 238996 5176 239002 5228
rect 289722 5176 289728 5228
rect 289780 5216 289786 5228
rect 347866 5216 347872 5228
rect 289780 5188 347872 5216
rect 289780 5176 289786 5188
rect 347866 5176 347872 5188
rect 347924 5176 347930 5228
rect 362770 5176 362776 5228
rect 362828 5216 362834 5228
rect 558362 5216 558368 5228
rect 362828 5188 558368 5216
rect 362828 5176 362834 5188
rect 558362 5176 558368 5188
rect 558420 5176 558426 5228
rect 48130 5108 48136 5160
rect 48188 5148 48194 5160
rect 186498 5148 186504 5160
rect 48188 5120 186504 5148
rect 48188 5108 48194 5120
rect 186498 5108 186504 5120
rect 186556 5108 186562 5160
rect 197998 5108 198004 5160
rect 198056 5148 198062 5160
rect 237650 5148 237656 5160
rect 198056 5120 237656 5148
rect 198056 5108 198062 5120
rect 237650 5108 237656 5120
rect 237708 5108 237714 5160
rect 291010 5108 291016 5160
rect 291068 5148 291074 5160
rect 351362 5148 351368 5160
rect 291068 5120 351368 5148
rect 291068 5108 291074 5120
rect 351362 5108 351368 5120
rect 351420 5108 351426 5160
rect 362678 5108 362684 5160
rect 362736 5148 362742 5160
rect 561950 5148 561956 5160
rect 362736 5120 561956 5148
rect 362736 5108 362742 5120
rect 561950 5108 561956 5120
rect 562008 5108 562014 5160
rect 17310 5040 17316 5092
rect 17368 5080 17374 5092
rect 175550 5080 175556 5092
rect 17368 5052 175556 5080
rect 17368 5040 17374 5052
rect 175550 5040 175556 5052
rect 175608 5040 175614 5092
rect 194410 5040 194416 5092
rect 194468 5080 194474 5092
rect 236362 5080 236368 5092
rect 194468 5052 236368 5080
rect 194468 5040 194474 5052
rect 236362 5040 236368 5052
rect 236420 5040 236426 5092
rect 292390 5040 292396 5092
rect 292448 5080 292454 5092
rect 354950 5080 354956 5092
rect 292448 5052 354956 5080
rect 292448 5040 292454 5052
rect 354950 5040 354956 5052
rect 355008 5040 355014 5092
rect 364242 5040 364248 5092
rect 364300 5080 364306 5092
rect 565538 5080 565544 5092
rect 364300 5052 565544 5080
rect 364300 5040 364306 5052
rect 565538 5040 565544 5052
rect 565596 5040 565602 5092
rect 12434 4972 12440 5024
rect 12492 5012 12498 5024
rect 174078 5012 174084 5024
rect 12492 4984 174084 5012
rect 12492 4972 12498 4984
rect 174078 4972 174084 4984
rect 174136 4972 174142 5024
rect 190822 4972 190828 5024
rect 190880 5012 190886 5024
rect 234890 5012 234896 5024
rect 190880 4984 234896 5012
rect 190880 4972 190886 4984
rect 234890 4972 234896 4984
rect 234948 4972 234954 5024
rect 293770 4972 293776 5024
rect 293828 5012 293834 5024
rect 358538 5012 358544 5024
rect 293828 4984 358544 5012
rect 293828 4972 293834 4984
rect 358538 4972 358544 4984
rect 358596 4972 358602 5024
rect 365530 4972 365536 5024
rect 365588 5012 365594 5024
rect 569034 5012 569040 5024
rect 365588 4984 569040 5012
rect 365588 4972 365594 4984
rect 569034 4972 569040 4984
rect 569092 4972 569098 5024
rect 7650 4904 7656 4956
rect 7708 4944 7714 4956
rect 172698 4944 172704 4956
rect 7708 4916 172704 4944
rect 7708 4904 7714 4916
rect 172698 4904 172704 4916
rect 172756 4904 172762 4956
rect 187234 4904 187240 4956
rect 187292 4944 187298 4956
rect 233326 4944 233332 4956
rect 187292 4916 233332 4944
rect 187292 4904 187298 4916
rect 233326 4904 233332 4916
rect 233384 4904 233390 4956
rect 295242 4904 295248 4956
rect 295300 4944 295306 4956
rect 362126 4944 362132 4956
rect 295300 4916 362132 4944
rect 295300 4904 295306 4916
rect 362126 4904 362132 4916
rect 362184 4904 362190 4956
rect 366726 4904 366732 4956
rect 366784 4944 366790 4956
rect 572622 4944 572628 4956
rect 366784 4916 572628 4944
rect 366784 4904 366790 4916
rect 572622 4904 572628 4916
rect 572680 4904 572686 4956
rect 2866 4836 2872 4888
rect 2924 4876 2930 4888
rect 169938 4876 169944 4888
rect 2924 4848 169944 4876
rect 2924 4836 2930 4848
rect 169938 4836 169944 4848
rect 169996 4836 170002 4888
rect 174170 4836 174176 4888
rect 174228 4876 174234 4888
rect 229094 4876 229100 4888
rect 174228 4848 229100 4876
rect 174228 4836 174234 4848
rect 229094 4836 229100 4848
rect 229152 4836 229158 4888
rect 296622 4836 296628 4888
rect 296680 4876 296686 4888
rect 365714 4876 365720 4888
rect 296680 4848 365720 4876
rect 296680 4836 296686 4848
rect 365714 4836 365720 4848
rect 365772 4836 365778 4888
rect 368290 4836 368296 4888
rect 368348 4876 368354 4888
rect 576210 4876 576216 4888
rect 368348 4848 576216 4876
rect 368348 4836 368354 4848
rect 576210 4836 576216 4848
rect 576268 4836 576274 4888
rect 1670 4768 1676 4820
rect 1728 4808 1734 4820
rect 169846 4808 169852 4820
rect 1728 4780 169852 4808
rect 1728 4768 1734 4780
rect 169846 4768 169852 4780
rect 169904 4768 169910 4820
rect 170582 4768 170588 4820
rect 170640 4808 170646 4820
rect 228174 4808 228180 4820
rect 170640 4780 228180 4808
rect 170640 4768 170646 4780
rect 228174 4768 228180 4780
rect 228232 4768 228238 4820
rect 298002 4768 298008 4820
rect 298060 4808 298066 4820
rect 369210 4808 369216 4820
rect 298060 4780 369216 4808
rect 298060 4768 298066 4780
rect 369210 4768 369216 4780
rect 369268 4768 369274 4820
rect 369670 4768 369676 4820
rect 369728 4808 369734 4820
rect 579798 4808 579804 4820
rect 369728 4780 579804 4808
rect 369728 4768 369734 4780
rect 579798 4768 579804 4780
rect 579856 4768 579862 4820
rect 69474 4700 69480 4752
rect 69532 4740 69538 4752
rect 193490 4740 193496 4752
rect 69532 4712 193496 4740
rect 69532 4700 69538 4712
rect 193490 4700 193496 4712
rect 193548 4700 193554 4752
rect 286594 4700 286600 4752
rect 286652 4740 286658 4752
rect 338298 4740 338304 4752
rect 286652 4712 338304 4740
rect 286652 4700 286658 4712
rect 338298 4700 338304 4712
rect 338356 4700 338362 4752
rect 355962 4700 355968 4752
rect 356020 4740 356026 4752
rect 540514 4740 540520 4752
rect 356020 4712 540520 4740
rect 356020 4700 356026 4712
rect 540514 4700 540520 4712
rect 540572 4700 540578 4752
rect 127802 4632 127808 4684
rect 127860 4672 127866 4684
rect 212810 4672 212816 4684
rect 127860 4644 212816 4672
rect 127860 4632 127866 4644
rect 212810 4632 212816 4644
rect 212868 4632 212874 4684
rect 286870 4632 286876 4684
rect 286928 4672 286934 4684
rect 337102 4672 337108 4684
rect 286928 4644 337108 4672
rect 286928 4632 286934 4644
rect 337102 4632 337108 4644
rect 337160 4632 337166 4684
rect 354582 4632 354588 4684
rect 354640 4672 354646 4684
rect 536926 4672 536932 4684
rect 354640 4644 536932 4672
rect 354640 4632 354646 4644
rect 536926 4632 536932 4644
rect 536984 4632 536990 4684
rect 144454 4564 144460 4616
rect 144512 4604 144518 4616
rect 219434 4604 219440 4616
rect 144512 4576 219440 4604
rect 144512 4564 144518 4576
rect 219434 4564 219440 4576
rect 219492 4564 219498 4616
rect 285306 4564 285312 4616
rect 285364 4604 285370 4616
rect 334710 4604 334716 4616
rect 285364 4576 334716 4604
rect 285364 4564 285370 4576
rect 334710 4564 334716 4576
rect 334768 4564 334774 4616
rect 353202 4564 353208 4616
rect 353260 4604 353266 4616
rect 533430 4604 533436 4616
rect 353260 4576 533436 4604
rect 353260 4564 353266 4576
rect 533430 4564 533436 4576
rect 533488 4564 533494 4616
rect 148042 4496 148048 4548
rect 148100 4536 148106 4548
rect 220814 4536 220820 4548
rect 148100 4508 220820 4536
rect 148100 4496 148106 4508
rect 220814 4496 220820 4508
rect 220872 4496 220878 4548
rect 283926 4496 283932 4548
rect 283984 4536 283990 4548
rect 331214 4536 331220 4548
rect 283984 4508 331220 4536
rect 283984 4496 283990 4508
rect 331214 4496 331220 4508
rect 331272 4496 331278 4548
rect 351730 4496 351736 4548
rect 351788 4536 351794 4548
rect 529842 4536 529848 4548
rect 351788 4508 529848 4536
rect 351788 4496 351794 4508
rect 529842 4496 529848 4508
rect 529900 4496 529906 4548
rect 151538 4428 151544 4480
rect 151596 4468 151602 4480
rect 220906 4468 220912 4480
rect 151596 4440 220912 4468
rect 151596 4428 151602 4440
rect 220906 4428 220912 4440
rect 220964 4428 220970 4480
rect 285490 4428 285496 4480
rect 285548 4468 285554 4480
rect 333606 4468 333612 4480
rect 285548 4440 333612 4468
rect 285548 4428 285554 4440
rect 333606 4428 333612 4440
rect 333664 4428 333670 4480
rect 351822 4428 351828 4480
rect 351880 4468 351886 4480
rect 526254 4468 526260 4480
rect 351880 4440 526260 4468
rect 351880 4428 351886 4440
rect 526254 4428 526260 4440
rect 526312 4428 526318 4480
rect 155126 4360 155132 4412
rect 155184 4400 155190 4412
rect 222194 4400 222200 4412
rect 155184 4372 222200 4400
rect 155184 4360 155190 4372
rect 222194 4360 222200 4372
rect 222252 4360 222258 4412
rect 284110 4360 284116 4412
rect 284168 4400 284174 4412
rect 330018 4400 330024 4412
rect 284168 4372 330024 4400
rect 284168 4360 284174 4372
rect 330018 4360 330024 4372
rect 330076 4360 330082 4412
rect 350442 4360 350448 4412
rect 350500 4400 350506 4412
rect 522666 4400 522672 4412
rect 350500 4372 522672 4400
rect 350500 4360 350506 4372
rect 522666 4360 522672 4372
rect 522724 4360 522730 4412
rect 158714 4292 158720 4344
rect 158772 4332 158778 4344
rect 223574 4332 223580 4344
rect 158772 4304 223580 4332
rect 158772 4292 158778 4304
rect 223574 4292 223580 4304
rect 223632 4292 223638 4344
rect 282730 4292 282736 4344
rect 282788 4332 282794 4344
rect 327626 4332 327632 4344
rect 282788 4304 327632 4332
rect 282788 4292 282794 4304
rect 327626 4292 327632 4304
rect 327684 4292 327690 4344
rect 348970 4292 348976 4344
rect 349028 4332 349034 4344
rect 519078 4332 519084 4344
rect 349028 4304 519084 4332
rect 349028 4292 349034 4304
rect 519078 4292 519084 4304
rect 519136 4292 519142 4344
rect 163498 4224 163504 4276
rect 163556 4264 163562 4276
rect 224954 4264 224960 4276
rect 163556 4236 224960 4264
rect 163556 4224 163562 4236
rect 224954 4224 224960 4236
rect 225012 4224 225018 4276
rect 281350 4224 281356 4276
rect 281408 4264 281414 4276
rect 324038 4264 324044 4276
rect 281408 4236 324044 4264
rect 281408 4224 281414 4236
rect 324038 4224 324044 4236
rect 324096 4224 324102 4276
rect 347682 4224 347688 4276
rect 347740 4264 347746 4276
rect 515582 4264 515588 4276
rect 347740 4236 515588 4264
rect 347740 4224 347746 4236
rect 515582 4224 515588 4236
rect 515640 4224 515646 4276
rect 167086 4156 167092 4208
rect 167144 4196 167150 4208
rect 226334 4196 226340 4208
rect 167144 4168 226340 4196
rect 167144 4156 167150 4168
rect 226334 4156 226340 4168
rect 226392 4156 226398 4208
rect 277210 4156 277216 4208
rect 277268 4196 277274 4208
rect 277268 4168 277808 4196
rect 277268 4156 277274 4168
rect 61194 4088 61200 4140
rect 61252 4128 61258 4140
rect 186958 4128 186964 4140
rect 61252 4100 186964 4128
rect 61252 4088 61258 4100
rect 186958 4088 186964 4100
rect 187016 4088 187022 4140
rect 199194 4088 199200 4140
rect 199252 4128 199258 4140
rect 203518 4128 203524 4140
rect 199252 4100 203524 4128
rect 199252 4088 199258 4100
rect 203518 4088 203524 4100
rect 203576 4088 203582 4140
rect 211062 4088 211068 4140
rect 211120 4128 211126 4140
rect 211798 4128 211804 4140
rect 211120 4100 211804 4128
rect 211120 4088 211126 4100
rect 211798 4088 211804 4100
rect 211856 4088 211862 4140
rect 214650 4088 214656 4140
rect 214708 4128 214714 4140
rect 215202 4128 215208 4140
rect 214708 4100 215208 4128
rect 214708 4088 214714 4100
rect 215202 4088 215208 4100
rect 215260 4088 215266 4140
rect 217042 4088 217048 4140
rect 217100 4128 217106 4140
rect 218698 4128 218704 4140
rect 217100 4100 218704 4128
rect 217100 4088 217106 4100
rect 218698 4088 218704 4100
rect 218756 4088 218762 4140
rect 221734 4088 221740 4140
rect 221792 4128 221798 4140
rect 245010 4128 245016 4140
rect 221792 4100 245016 4128
rect 221792 4088 221798 4100
rect 245010 4088 245016 4100
rect 245068 4088 245074 4140
rect 257430 4088 257436 4140
rect 257488 4128 257494 4140
rect 257982 4128 257988 4140
rect 257488 4100 257988 4128
rect 257488 4088 257494 4100
rect 257982 4088 257988 4100
rect 258040 4088 258046 4140
rect 258166 4088 258172 4140
rect 258224 4128 258230 4140
rect 258626 4128 258632 4140
rect 258224 4100 258632 4128
rect 258224 4088 258230 4100
rect 258626 4088 258632 4100
rect 258684 4088 258690 4140
rect 259362 4088 259368 4140
rect 259420 4128 259426 4140
rect 259822 4128 259828 4140
rect 259420 4100 259828 4128
rect 259420 4088 259426 4100
rect 259822 4088 259828 4100
rect 259880 4088 259886 4140
rect 261478 4088 261484 4140
rect 261536 4128 261542 4140
rect 262214 4128 262220 4140
rect 261536 4100 262220 4128
rect 261536 4088 261542 4100
rect 262214 4088 262220 4100
rect 262272 4088 262278 4140
rect 264606 4128 264612 4140
rect 262416 4100 264612 4128
rect 54018 4020 54024 4072
rect 54076 4060 54082 4072
rect 185578 4060 185584 4072
rect 54076 4032 185584 4060
rect 54076 4020 54082 4032
rect 185578 4020 185584 4032
rect 185636 4020 185642 4072
rect 206278 4020 206284 4072
rect 206336 4060 206342 4072
rect 211890 4060 211896 4072
rect 206336 4032 211896 4060
rect 206336 4020 206342 4032
rect 211890 4020 211896 4032
rect 211948 4020 211954 4072
rect 215846 4020 215852 4072
rect 215904 4060 215910 4072
rect 238757 4063 238815 4069
rect 238757 4060 238769 4063
rect 215904 4032 238769 4060
rect 215904 4020 215910 4032
rect 238757 4029 238769 4032
rect 238803 4029 238815 4063
rect 238757 4023 238815 4029
rect 240778 4020 240784 4072
rect 240836 4060 240842 4072
rect 241422 4060 241428 4072
rect 240836 4032 241428 4060
rect 240836 4020 240842 4032
rect 241422 4020 241428 4032
rect 241480 4020 241486 4072
rect 261570 4020 261576 4072
rect 261628 4060 261634 4072
rect 262416 4060 262444 4100
rect 264606 4088 264612 4100
rect 264664 4088 264670 4140
rect 269758 4088 269764 4140
rect 269816 4128 269822 4140
rect 272886 4128 272892 4140
rect 269816 4100 272892 4128
rect 269816 4088 269822 4100
rect 272886 4088 272892 4100
rect 272944 4088 272950 4140
rect 272996 4100 276612 4128
rect 261628 4032 262444 4060
rect 261628 4020 261634 4032
rect 263502 4020 263508 4072
rect 263560 4060 263566 4072
rect 270494 4060 270500 4072
rect 263560 4032 270500 4060
rect 263560 4020 263566 4032
rect 270494 4020 270500 4032
rect 270552 4020 270558 4072
rect 272996 4060 273024 4100
rect 270604 4032 273024 4060
rect 273073 4063 273131 4069
rect 14826 3952 14832 4004
rect 14884 3992 14890 4004
rect 17218 3992 17224 4004
rect 14884 3964 17224 3992
rect 14884 3952 14890 3964
rect 17218 3952 17224 3964
rect 17276 3952 17282 4004
rect 43346 3952 43352 4004
rect 43404 3992 43410 4004
rect 183830 3992 183836 4004
rect 43404 3964 183836 3992
rect 43404 3952 43410 3964
rect 183830 3952 183836 3964
rect 183888 3952 183894 4004
rect 213454 3952 213460 4004
rect 213512 3992 213518 4004
rect 234709 3995 234767 4001
rect 234709 3992 234721 3995
rect 213512 3964 234721 3992
rect 213512 3952 213518 3964
rect 234709 3961 234721 3964
rect 234755 3961 234767 3995
rect 234709 3955 234767 3961
rect 234798 3952 234804 4004
rect 234856 3992 234862 4004
rect 247770 3992 247776 4004
rect 234856 3964 247776 3992
rect 234856 3952 234862 3964
rect 247770 3952 247776 3964
rect 247828 3952 247834 4004
rect 267550 3952 267556 4004
rect 267608 3992 267614 4004
rect 270604 3992 270632 4032
rect 273073 4029 273085 4063
rect 273119 4060 273131 4063
rect 276474 4060 276480 4072
rect 273119 4032 276480 4060
rect 273119 4029 273131 4032
rect 273073 4023 273131 4029
rect 276474 4020 276480 4032
rect 276532 4020 276538 4072
rect 276584 4060 276612 4100
rect 276658 4088 276664 4140
rect 276716 4128 276722 4140
rect 277670 4128 277676 4140
rect 276716 4100 277676 4128
rect 276716 4088 276722 4100
rect 277670 4088 277676 4100
rect 277728 4088 277734 4140
rect 277780 4128 277808 4168
rect 279970 4156 279976 4208
rect 280028 4196 280034 4208
rect 320450 4196 320456 4208
rect 280028 4168 320456 4196
rect 280028 4156 280034 4168
rect 320450 4156 320456 4168
rect 320508 4156 320514 4208
rect 346302 4156 346308 4208
rect 346360 4196 346366 4208
rect 511994 4196 512000 4208
rect 346360 4168 512000 4196
rect 346360 4156 346366 4168
rect 511994 4156 512000 4168
rect 512052 4156 512058 4208
rect 277780 4100 278268 4128
rect 278133 4063 278191 4069
rect 278133 4060 278145 4063
rect 276584 4032 278145 4060
rect 278133 4029 278145 4032
rect 278179 4029 278191 4063
rect 278240 4060 278268 4100
rect 279418 4088 279424 4140
rect 279476 4128 279482 4140
rect 282454 4128 282460 4140
rect 279476 4100 282460 4128
rect 279476 4088 279482 4100
rect 282454 4088 282460 4100
rect 282512 4088 282518 4140
rect 283650 4088 283656 4140
rect 283708 4128 283714 4140
rect 283708 4100 286180 4128
rect 283708 4088 283714 4100
rect 286045 4063 286103 4069
rect 286045 4060 286057 4063
rect 278240 4032 286057 4060
rect 278133 4023 278191 4029
rect 286045 4029 286057 4032
rect 286091 4029 286103 4063
rect 286045 4023 286103 4029
rect 267608 3964 270632 3992
rect 267608 3952 267614 3964
rect 272794 3952 272800 4004
rect 272852 3992 272858 4004
rect 277949 3995 278007 4001
rect 277949 3992 277961 3995
rect 272852 3964 277961 3992
rect 272852 3952 272858 3964
rect 277949 3961 277961 3964
rect 277995 3961 278007 3995
rect 285950 3992 285956 4004
rect 277949 3955 278007 3961
rect 278056 3964 285956 3992
rect 42150 3884 42156 3936
rect 42208 3924 42214 3936
rect 183922 3924 183928 3936
rect 42208 3896 183928 3924
rect 42208 3884 42214 3896
rect 183922 3884 183928 3896
rect 183980 3884 183986 3936
rect 195606 3884 195612 3936
rect 195664 3924 195670 3936
rect 225233 3927 225291 3933
rect 225233 3924 225245 3927
rect 195664 3896 225245 3924
rect 195664 3884 195670 3896
rect 225233 3893 225245 3896
rect 225279 3893 225291 3927
rect 225233 3887 225291 3893
rect 225322 3884 225328 3936
rect 225380 3924 225386 3936
rect 226242 3924 226248 3936
rect 225380 3896 226248 3924
rect 225380 3884 225386 3896
rect 226242 3884 226248 3896
rect 226300 3884 226306 3936
rect 226337 3927 226395 3933
rect 226337 3893 226349 3927
rect 226383 3924 226395 3927
rect 233234 3924 233240 3936
rect 226383 3896 233240 3924
rect 226383 3893 226395 3896
rect 226337 3887 226395 3893
rect 233234 3884 233240 3896
rect 233292 3884 233298 3936
rect 233694 3884 233700 3936
rect 233752 3924 233758 3936
rect 240686 3924 240692 3936
rect 233752 3896 240692 3924
rect 233752 3884 233758 3896
rect 240686 3884 240692 3896
rect 240744 3884 240750 3936
rect 241974 3884 241980 3936
rect 242032 3924 242038 3936
rect 249150 3924 249156 3936
rect 242032 3896 249156 3924
rect 242032 3884 242038 3896
rect 249150 3884 249156 3896
rect 249208 3884 249214 3936
rect 268746 3884 268752 3936
rect 268804 3924 268810 3936
rect 278056 3924 278084 3964
rect 285950 3952 285956 3964
rect 286008 3952 286014 4004
rect 286152 3992 286180 4100
rect 286962 4088 286968 4140
rect 287020 4128 287026 4140
rect 287885 4131 287943 4137
rect 287885 4128 287897 4131
rect 287020 4100 287897 4128
rect 287020 4088 287026 4100
rect 287885 4097 287897 4100
rect 287931 4097 287943 4131
rect 287885 4091 287943 4097
rect 287977 4131 288035 4137
rect 287977 4097 287989 4131
rect 288023 4128 288035 4131
rect 306374 4128 306380 4140
rect 288023 4100 306380 4128
rect 288023 4097 288035 4100
rect 287977 4091 288035 4097
rect 306374 4088 306380 4100
rect 306432 4088 306438 4140
rect 352466 4088 352472 4140
rect 352524 4128 352530 4140
rect 460842 4128 460848 4140
rect 352524 4100 460848 4128
rect 352524 4088 352530 4100
rect 460842 4088 460848 4100
rect 460900 4088 460906 4140
rect 469858 4088 469864 4140
rect 469916 4128 469922 4140
rect 550082 4128 550088 4140
rect 469916 4100 550088 4128
rect 469916 4088 469922 4100
rect 550082 4088 550088 4100
rect 550140 4088 550146 4140
rect 286229 4063 286287 4069
rect 286229 4029 286241 4063
rect 286275 4060 286287 4063
rect 310974 4060 310980 4072
rect 286275 4032 310980 4060
rect 286275 4029 286287 4032
rect 286229 4023 286287 4029
rect 310974 4020 310980 4032
rect 311032 4020 311038 4072
rect 311066 4020 311072 4072
rect 311124 4060 311130 4072
rect 316954 4060 316960 4072
rect 311124 4032 316960 4060
rect 311124 4020 311130 4032
rect 316954 4020 316960 4032
rect 317012 4020 317018 4072
rect 345658 4020 345664 4072
rect 345716 4060 345722 4072
rect 453666 4060 453672 4072
rect 345716 4032 453672 4060
rect 345716 4020 345722 4032
rect 453666 4020 453672 4032
rect 453724 4020 453730 4072
rect 473998 4020 474004 4072
rect 474056 4060 474062 4072
rect 557166 4060 557172 4072
rect 474056 4032 557172 4060
rect 474056 4020 474062 4032
rect 557166 4020 557172 4032
rect 557224 4020 557230 4072
rect 287517 3995 287575 4001
rect 287517 3992 287529 3995
rect 286152 3964 287529 3992
rect 287517 3961 287529 3964
rect 287563 3961 287575 3995
rect 287517 3955 287575 3961
rect 287701 3995 287759 4001
rect 287701 3961 287713 3995
rect 287747 3992 287759 3995
rect 314562 3992 314568 4004
rect 287747 3964 314568 3992
rect 287747 3961 287759 3964
rect 287701 3955 287759 3961
rect 314562 3952 314568 3964
rect 314620 3952 314626 4004
rect 316678 3952 316684 4004
rect 316736 3992 316742 4004
rect 328822 3992 328828 4004
rect 316736 3964 328828 3992
rect 316736 3952 316742 3964
rect 328822 3952 328828 3964
rect 328880 3952 328886 4004
rect 330478 3952 330484 4004
rect 330536 3992 330542 4004
rect 439406 3992 439412 4004
rect 330536 3964 439412 3992
rect 330536 3952 330542 3964
rect 439406 3952 439412 3964
rect 439464 3952 439470 4004
rect 475378 3952 475384 4004
rect 475436 3992 475442 4004
rect 564342 3992 564348 4004
rect 475436 3964 564348 3992
rect 475436 3952 475442 3964
rect 564342 3952 564348 3964
rect 564400 3952 564406 4004
rect 268804 3896 278084 3924
rect 278133 3927 278191 3933
rect 268804 3884 268810 3896
rect 278133 3893 278145 3927
rect 278179 3924 278191 3927
rect 283650 3924 283656 3936
rect 278179 3896 283656 3924
rect 278179 3893 278191 3896
rect 278133 3887 278191 3893
rect 283650 3884 283656 3896
rect 283708 3884 283714 3936
rect 285582 3884 285588 3936
rect 285640 3924 285646 3936
rect 287606 3924 287612 3936
rect 285640 3896 287612 3924
rect 285640 3884 285646 3896
rect 287606 3884 287612 3896
rect 287664 3884 287670 3936
rect 318058 3924 318064 3936
rect 287716 3896 318064 3924
rect 24302 3816 24308 3868
rect 24360 3856 24366 3868
rect 31018 3856 31024 3868
rect 24360 3828 31024 3856
rect 24360 3816 24366 3828
rect 31018 3816 31024 3828
rect 31076 3816 31082 3868
rect 36170 3816 36176 3868
rect 36228 3856 36234 3868
rect 182358 3856 182364 3868
rect 36228 3828 182364 3856
rect 36228 3816 36234 3828
rect 182358 3816 182364 3828
rect 182416 3816 182422 3868
rect 192018 3816 192024 3868
rect 192076 3856 192082 3868
rect 235258 3856 235264 3868
rect 192076 3828 235264 3856
rect 192076 3816 192082 3828
rect 235258 3816 235264 3828
rect 235316 3816 235322 3868
rect 238757 3859 238815 3865
rect 238757 3825 238769 3859
rect 238803 3856 238815 3859
rect 242986 3856 242992 3868
rect 238803 3828 242992 3856
rect 238803 3825 238815 3828
rect 238757 3819 238815 3825
rect 242986 3816 242992 3828
rect 243044 3816 243050 3868
rect 265618 3816 265624 3868
rect 265676 3856 265682 3868
rect 273073 3859 273131 3865
rect 273073 3856 273085 3859
rect 265676 3828 273085 3856
rect 265676 3816 265682 3828
rect 273073 3825 273085 3828
rect 273119 3825 273131 3859
rect 273073 3819 273131 3825
rect 273165 3859 273223 3865
rect 273165 3825 273177 3859
rect 273211 3856 273223 3859
rect 274361 3859 274419 3865
rect 273211 3828 274312 3856
rect 273211 3825 273223 3828
rect 273165 3819 273223 3825
rect 25498 3748 25504 3800
rect 25556 3788 25562 3800
rect 32398 3788 32404 3800
rect 25556 3760 32404 3788
rect 25556 3748 25562 3760
rect 32398 3748 32404 3760
rect 32456 3748 32462 3800
rect 34974 3748 34980 3800
rect 35032 3788 35038 3800
rect 181070 3788 181076 3800
rect 35032 3760 181076 3788
rect 35032 3748 35038 3760
rect 181070 3748 181076 3760
rect 181128 3748 181134 3800
rect 193214 3748 193220 3800
rect 193272 3788 193278 3800
rect 225141 3791 225199 3797
rect 225141 3788 225153 3791
rect 193272 3760 225153 3788
rect 193272 3748 193278 3760
rect 225141 3757 225153 3760
rect 225187 3757 225199 3791
rect 225141 3751 225199 3757
rect 225233 3791 225291 3797
rect 225233 3757 225245 3791
rect 225279 3788 225291 3791
rect 235994 3788 236000 3800
rect 225279 3760 236000 3788
rect 225279 3757 225291 3760
rect 225233 3751 225291 3757
rect 235994 3748 236000 3760
rect 236052 3748 236058 3800
rect 246758 3748 246764 3800
rect 246816 3788 246822 3800
rect 254118 3788 254124 3800
rect 246816 3760 254124 3788
rect 246816 3748 246822 3760
rect 254118 3748 254124 3760
rect 254176 3748 254182 3800
rect 267642 3748 267648 3800
rect 267700 3788 267706 3800
rect 274177 3791 274235 3797
rect 274177 3788 274189 3791
rect 267700 3760 274189 3788
rect 267700 3748 267706 3760
rect 274177 3757 274189 3760
rect 274223 3757 274235 3791
rect 274284 3788 274312 3828
rect 274361 3825 274373 3859
rect 274407 3856 274419 3859
rect 287146 3856 287152 3868
rect 274407 3828 287152 3856
rect 274407 3825 274419 3828
rect 274361 3819 274419 3825
rect 287146 3816 287152 3828
rect 287204 3816 287210 3868
rect 278866 3788 278872 3800
rect 274284 3760 278872 3788
rect 274177 3751 274235 3757
rect 278866 3748 278872 3760
rect 278924 3748 278930 3800
rect 280062 3748 280068 3800
rect 280120 3788 280126 3800
rect 287716 3788 287744 3896
rect 318058 3884 318064 3896
rect 318116 3884 318122 3936
rect 337378 3884 337384 3936
rect 337436 3924 337442 3936
rect 467926 3924 467932 3936
rect 337436 3896 467932 3924
rect 337436 3884 337442 3896
rect 467926 3884 467932 3896
rect 467984 3884 467990 3936
rect 478138 3884 478144 3936
rect 478196 3924 478202 3936
rect 571426 3924 571432 3936
rect 478196 3896 571432 3924
rect 478196 3884 478202 3896
rect 571426 3884 571432 3896
rect 571484 3884 571490 3936
rect 321646 3856 321652 3868
rect 280120 3760 287744 3788
rect 287808 3828 321652 3856
rect 280120 3748 280126 3760
rect 16022 3680 16028 3732
rect 16080 3720 16086 3732
rect 24118 3720 24124 3732
rect 16080 3692 24124 3720
rect 16080 3680 16086 3692
rect 24118 3680 24124 3692
rect 24176 3680 24182 3732
rect 29086 3680 29092 3732
rect 29144 3720 29150 3732
rect 179414 3720 179420 3732
rect 29144 3692 179420 3720
rect 29144 3680 29150 3692
rect 179414 3680 179420 3692
rect 179472 3680 179478 3732
rect 189626 3680 189632 3732
rect 189684 3720 189690 3732
rect 234614 3720 234620 3732
rect 189684 3692 234620 3720
rect 189684 3680 189690 3692
rect 234614 3680 234620 3692
rect 234672 3680 234678 3732
rect 234801 3723 234859 3729
rect 234801 3689 234813 3723
rect 234847 3720 234859 3723
rect 243078 3720 243084 3732
rect 234847 3692 243084 3720
rect 234847 3689 234859 3692
rect 234801 3683 234859 3689
rect 243078 3680 243084 3692
rect 243136 3680 243142 3732
rect 243170 3680 243176 3732
rect 243228 3720 243234 3732
rect 251818 3720 251824 3732
rect 243228 3692 251824 3720
rect 243228 3680 243234 3692
rect 251818 3680 251824 3692
rect 251876 3680 251882 3732
rect 262122 3680 262128 3732
rect 262180 3720 262186 3732
rect 268102 3720 268108 3732
rect 262180 3692 268108 3720
rect 262180 3680 262186 3692
rect 268102 3680 268108 3692
rect 268160 3680 268166 3732
rect 270402 3680 270408 3732
rect 270460 3720 270466 3732
rect 278041 3723 278099 3729
rect 278041 3720 278053 3723
rect 270460 3692 278053 3720
rect 270460 3680 270466 3692
rect 278041 3689 278053 3692
rect 278087 3689 278099 3723
rect 278041 3683 278099 3689
rect 278682 3680 278688 3732
rect 278740 3720 278746 3732
rect 287701 3723 287759 3729
rect 287701 3720 287713 3723
rect 278740 3692 287713 3720
rect 278740 3680 278746 3692
rect 287701 3689 287713 3692
rect 287747 3689 287759 3723
rect 287701 3683 287759 3689
rect 20714 3612 20720 3664
rect 20772 3652 20778 3664
rect 176746 3652 176752 3664
rect 20772 3624 176752 3652
rect 20772 3612 20778 3624
rect 176746 3612 176752 3624
rect 176804 3612 176810 3664
rect 188430 3612 188436 3664
rect 188488 3652 188494 3664
rect 234706 3652 234712 3664
rect 188488 3624 234712 3652
rect 188488 3612 188494 3624
rect 234706 3612 234712 3624
rect 234764 3612 234770 3664
rect 239582 3612 239588 3664
rect 239640 3652 239646 3664
rect 250438 3652 250444 3664
rect 239640 3624 250444 3652
rect 239640 3612 239646 3624
rect 250438 3612 250444 3624
rect 250496 3612 250502 3664
rect 266170 3612 266176 3664
rect 266228 3652 266234 3664
rect 273165 3655 273223 3661
rect 273165 3652 273177 3655
rect 266228 3624 273177 3652
rect 266228 3612 266234 3624
rect 273165 3621 273177 3624
rect 273211 3621 273223 3655
rect 273165 3615 273223 3621
rect 274177 3655 274235 3661
rect 274177 3621 274189 3655
rect 274223 3652 274235 3655
rect 281258 3652 281264 3664
rect 274223 3624 281264 3652
rect 274223 3621 274235 3624
rect 274177 3615 274235 3621
rect 281258 3612 281264 3624
rect 281316 3612 281322 3664
rect 281442 3612 281448 3664
rect 281500 3652 281506 3664
rect 287808 3652 287836 3828
rect 321646 3816 321652 3828
rect 321704 3816 321710 3868
rect 333882 3816 333888 3868
rect 333940 3856 333946 3868
rect 475102 3856 475108 3868
rect 333940 3828 475108 3856
rect 333940 3816 333946 3828
rect 475102 3816 475108 3828
rect 475160 3816 475166 3868
rect 477494 3816 477500 3868
rect 477552 3856 477558 3868
rect 478690 3856 478696 3868
rect 477552 3828 478696 3856
rect 477552 3816 477558 3828
rect 478690 3816 478696 3828
rect 478748 3816 478754 3868
rect 480898 3816 480904 3868
rect 480956 3856 480962 3868
rect 578602 3856 578608 3868
rect 480956 3828 578608 3856
rect 480956 3816 480962 3828
rect 578602 3816 578608 3828
rect 578660 3816 578666 3868
rect 287974 3748 287980 3800
rect 288032 3788 288038 3800
rect 335906 3788 335912 3800
rect 288032 3760 335912 3788
rect 288032 3748 288038 3760
rect 335906 3748 335912 3760
rect 335964 3748 335970 3800
rect 336642 3748 336648 3800
rect 336700 3788 336706 3800
rect 482278 3788 482284 3800
rect 336700 3760 482284 3788
rect 336700 3748 336706 3760
rect 482278 3748 482284 3760
rect 482336 3748 482342 3800
rect 520274 3748 520280 3800
rect 520332 3788 520338 3800
rect 521470 3788 521476 3800
rect 520332 3760 521476 3788
rect 520332 3748 520338 3760
rect 521470 3748 521476 3760
rect 521528 3748 521534 3800
rect 287885 3723 287943 3729
rect 287885 3689 287897 3723
rect 287931 3720 287943 3723
rect 339494 3720 339500 3732
rect 287931 3692 339500 3720
rect 287931 3689 287943 3692
rect 287885 3683 287943 3689
rect 339494 3680 339500 3692
rect 339552 3680 339558 3732
rect 360102 3680 360108 3732
rect 360160 3720 360166 3732
rect 553578 3720 553584 3732
rect 360160 3692 553584 3720
rect 360160 3680 360166 3692
rect 553578 3680 553584 3692
rect 553636 3680 553642 3732
rect 281500 3624 287836 3652
rect 281500 3612 281506 3624
rect 288342 3612 288348 3664
rect 288400 3652 288406 3664
rect 343082 3652 343088 3664
rect 288400 3624 343088 3652
rect 288400 3612 288406 3624
rect 343082 3612 343088 3624
rect 343140 3612 343146 3664
rect 362862 3612 362868 3664
rect 362920 3652 362926 3664
rect 560754 3652 560760 3664
rect 362920 3624 560760 3652
rect 362920 3612 362926 3624
rect 560754 3612 560760 3624
rect 560812 3612 560818 3664
rect 19518 3544 19524 3596
rect 19576 3584 19582 3596
rect 176654 3584 176660 3596
rect 19576 3556 176660 3584
rect 19576 3544 19582 3556
rect 176654 3544 176660 3556
rect 176712 3544 176718 3596
rect 183738 3544 183744 3596
rect 183796 3584 183802 3596
rect 231854 3584 231860 3596
rect 183796 3556 231860 3584
rect 183796 3544 183802 3556
rect 231854 3544 231860 3556
rect 231912 3544 231918 3596
rect 236086 3584 236092 3596
rect 235368 3556 236092 3584
rect 6454 3476 6460 3528
rect 6512 3516 6518 3528
rect 10318 3516 10324 3528
rect 6512 3488 10324 3516
rect 6512 3476 6518 3488
rect 10318 3476 10324 3488
rect 10376 3476 10382 3528
rect 11238 3476 11244 3528
rect 11296 3516 11302 3528
rect 173158 3516 173164 3528
rect 11296 3488 173164 3516
rect 11296 3476 11302 3488
rect 173158 3476 173164 3488
rect 173216 3476 173222 3528
rect 184842 3476 184848 3528
rect 184900 3516 184906 3528
rect 225049 3519 225107 3525
rect 225049 3516 225061 3519
rect 184900 3488 225061 3516
rect 184900 3476 184906 3488
rect 225049 3485 225061 3488
rect 225095 3485 225107 3519
rect 225049 3479 225107 3485
rect 225141 3519 225199 3525
rect 225141 3485 225153 3519
rect 225187 3516 225199 3519
rect 235368 3516 235396 3556
rect 236086 3544 236092 3556
rect 236144 3544 236150 3596
rect 244366 3544 244372 3596
rect 244424 3584 244430 3596
rect 245562 3584 245568 3596
rect 244424 3556 245568 3584
rect 244424 3544 244430 3556
rect 245562 3544 245568 3556
rect 245620 3544 245626 3596
rect 263410 3544 263416 3596
rect 263468 3584 263474 3596
rect 269298 3584 269304 3596
rect 263468 3556 269304 3584
rect 263468 3544 263474 3556
rect 269298 3544 269304 3556
rect 269356 3544 269362 3596
rect 270126 3544 270132 3596
rect 270184 3584 270190 3596
rect 290734 3584 290740 3596
rect 270184 3556 290740 3584
rect 270184 3544 270190 3556
rect 290734 3544 290740 3556
rect 290792 3544 290798 3596
rect 291102 3544 291108 3596
rect 291160 3584 291166 3596
rect 350258 3584 350264 3596
rect 291160 3556 350264 3584
rect 291160 3544 291166 3556
rect 350258 3544 350264 3556
rect 350316 3544 350322 3596
rect 365622 3544 365628 3596
rect 365680 3584 365686 3596
rect 567838 3584 567844 3596
rect 365680 3556 567844 3584
rect 365680 3544 365686 3556
rect 567838 3544 567844 3556
rect 567896 3544 567902 3596
rect 225187 3488 235396 3516
rect 225187 3485 225199 3488
rect 225141 3479 225199 3485
rect 235994 3476 236000 3528
rect 236052 3516 236058 3528
rect 249978 3516 249984 3528
rect 236052 3488 249984 3516
rect 236052 3476 236058 3488
rect 249978 3476 249984 3488
rect 250036 3476 250042 3528
rect 251450 3476 251456 3528
rect 251508 3516 251514 3528
rect 252462 3516 252468 3528
rect 251508 3488 252468 3516
rect 251508 3476 251514 3488
rect 252462 3476 252468 3488
rect 252520 3476 252526 3528
rect 266262 3476 266268 3528
rect 266320 3516 266326 3528
rect 266320 3488 271828 3516
rect 266320 3476 266326 3488
rect 10042 3408 10048 3460
rect 10100 3448 10106 3460
rect 172882 3448 172888 3460
rect 10100 3420 172888 3448
rect 10100 3408 10106 3420
rect 172882 3408 172888 3420
rect 172940 3408 172946 3460
rect 181346 3408 181352 3460
rect 181404 3448 181410 3460
rect 181404 3420 226472 3448
rect 181404 3408 181410 3420
rect 27890 3340 27896 3392
rect 27948 3380 27954 3392
rect 28902 3380 28908 3392
rect 27948 3352 28908 3380
rect 27948 3340 27954 3352
rect 28902 3340 28908 3352
rect 28960 3340 28966 3392
rect 32674 3340 32680 3392
rect 32732 3380 32738 3392
rect 35158 3380 35164 3392
rect 32732 3352 35164 3380
rect 32732 3340 32738 3352
rect 35158 3340 35164 3352
rect 35216 3340 35222 3392
rect 39758 3340 39764 3392
rect 39816 3380 39822 3392
rect 42058 3380 42064 3392
rect 39816 3352 42064 3380
rect 39816 3340 39822 3352
rect 42058 3340 42064 3352
rect 42116 3340 42122 3392
rect 70670 3340 70676 3392
rect 70728 3380 70734 3392
rect 71682 3380 71688 3392
rect 70728 3352 71688 3380
rect 70728 3340 70734 3352
rect 71682 3340 71688 3352
rect 71740 3340 71746 3392
rect 188338 3380 188344 3392
rect 71792 3352 188344 3380
rect 38562 3272 38568 3324
rect 38620 3312 38626 3324
rect 67913 3315 67971 3321
rect 67913 3312 67925 3315
rect 38620 3284 67925 3312
rect 38620 3272 38626 3284
rect 67913 3281 67925 3284
rect 67959 3281 67971 3315
rect 67913 3275 67971 3281
rect 68278 3272 68284 3324
rect 68336 3312 68342 3324
rect 71792 3312 71820 3352
rect 188338 3340 188344 3352
rect 188396 3340 188402 3392
rect 224957 3383 225015 3389
rect 224957 3380 224969 3383
rect 224880 3352 224969 3380
rect 68336 3284 71820 3312
rect 74537 3315 74595 3321
rect 68336 3272 68342 3284
rect 74537 3281 74549 3315
rect 74583 3312 74595 3315
rect 77757 3315 77815 3321
rect 77757 3312 77769 3315
rect 74583 3284 77769 3312
rect 74583 3281 74595 3284
rect 74537 3275 74595 3281
rect 77757 3281 77769 3284
rect 77803 3281 77815 3315
rect 77757 3275 77815 3281
rect 77846 3272 77852 3324
rect 77904 3312 77910 3324
rect 78582 3312 78588 3324
rect 77904 3284 78588 3312
rect 77904 3272 77910 3284
rect 78582 3272 78588 3284
rect 78640 3272 78646 3324
rect 78953 3315 79011 3321
rect 78953 3281 78965 3315
rect 78999 3312 79011 3315
rect 81345 3315 81403 3321
rect 81345 3312 81357 3315
rect 78999 3284 81357 3312
rect 78999 3281 79011 3284
rect 78953 3275 79011 3281
rect 81345 3281 81357 3284
rect 81391 3281 81403 3315
rect 81345 3275 81403 3281
rect 81434 3272 81440 3324
rect 81492 3312 81498 3324
rect 82722 3312 82728 3324
rect 81492 3284 82728 3312
rect 81492 3272 81498 3284
rect 82722 3272 82728 3284
rect 82780 3272 82786 3324
rect 82817 3315 82875 3321
rect 82817 3281 82829 3315
rect 82863 3312 82875 3315
rect 191006 3312 191012 3324
rect 82863 3284 191012 3312
rect 82863 3281 82875 3284
rect 82817 3275 82875 3281
rect 191006 3272 191012 3284
rect 191064 3272 191070 3324
rect 45738 3204 45744 3256
rect 45796 3244 45802 3256
rect 69661 3247 69719 3253
rect 69661 3244 69673 3247
rect 45796 3216 69673 3244
rect 45796 3204 45802 3216
rect 69661 3213 69673 3216
rect 69707 3213 69719 3247
rect 69661 3207 69719 3213
rect 69753 3247 69811 3253
rect 69753 3213 69765 3247
rect 69799 3244 69811 3247
rect 71038 3244 71044 3256
rect 69799 3216 71044 3244
rect 69799 3213 69811 3216
rect 69753 3207 69811 3213
rect 71038 3204 71044 3216
rect 71096 3204 71102 3256
rect 84930 3204 84936 3256
rect 84988 3244 84994 3256
rect 85482 3244 85488 3256
rect 84988 3216 85488 3244
rect 84988 3204 84994 3216
rect 85482 3204 85488 3216
rect 85540 3204 85546 3256
rect 192570 3244 192576 3256
rect 87708 3216 192576 3244
rect 57606 3136 57612 3188
rect 57664 3176 57670 3188
rect 79413 3179 79471 3185
rect 79413 3176 79425 3179
rect 57664 3148 79425 3176
rect 57664 3136 57670 3148
rect 79413 3145 79425 3148
rect 79459 3145 79471 3179
rect 79413 3139 79471 3145
rect 79505 3179 79563 3185
rect 79505 3145 79517 3179
rect 79551 3176 79563 3179
rect 82541 3179 82599 3185
rect 82541 3176 82553 3179
rect 79551 3148 82553 3176
rect 79551 3145 79563 3148
rect 79505 3139 79563 3145
rect 82541 3145 82553 3148
rect 82587 3145 82599 3179
rect 82541 3139 82599 3145
rect 82630 3136 82636 3188
rect 82688 3176 82694 3188
rect 87708 3176 87736 3216
rect 192570 3204 192576 3216
rect 192628 3204 192634 3256
rect 196802 3204 196808 3256
rect 196860 3244 196866 3256
rect 204898 3244 204904 3256
rect 196860 3216 204904 3244
rect 196860 3204 196866 3216
rect 204898 3204 204904 3216
rect 204956 3204 204962 3256
rect 209866 3204 209872 3256
rect 209924 3244 209930 3256
rect 224880 3244 224908 3352
rect 224957 3349 224969 3352
rect 225003 3349 225015 3383
rect 224957 3343 225015 3349
rect 225049 3383 225107 3389
rect 225049 3349 225061 3383
rect 225095 3380 225107 3383
rect 226337 3383 226395 3389
rect 226337 3380 226349 3383
rect 225095 3352 226349 3380
rect 225095 3349 225107 3352
rect 225049 3343 225107 3349
rect 226337 3349 226349 3352
rect 226383 3349 226395 3383
rect 226444 3380 226472 3420
rect 226518 3408 226524 3460
rect 226576 3448 226582 3460
rect 227622 3448 227628 3460
rect 226576 3420 227628 3448
rect 226576 3408 226582 3420
rect 227622 3408 227628 3420
rect 227680 3408 227686 3460
rect 228729 3451 228787 3457
rect 228729 3417 228741 3451
rect 228775 3448 228787 3451
rect 232406 3448 232412 3460
rect 228775 3420 232412 3448
rect 228775 3417 228787 3420
rect 228729 3411 228787 3417
rect 232406 3408 232412 3420
rect 232464 3408 232470 3460
rect 232498 3408 232504 3460
rect 232556 3448 232562 3460
rect 249058 3448 249064 3460
rect 232556 3420 249064 3448
rect 232556 3408 232562 3420
rect 249058 3408 249064 3420
rect 249116 3408 249122 3460
rect 249150 3408 249156 3460
rect 249208 3448 249214 3460
rect 251910 3448 251916 3460
rect 249208 3420 251916 3448
rect 249208 3408 249214 3420
rect 251910 3408 251916 3420
rect 251968 3408 251974 3460
rect 263318 3408 263324 3460
rect 263376 3448 263382 3460
rect 271690 3448 271696 3460
rect 263376 3420 271696 3448
rect 263376 3408 263382 3420
rect 271690 3408 271696 3420
rect 271748 3408 271754 3460
rect 271800 3448 271828 3488
rect 272518 3476 272524 3528
rect 272576 3516 272582 3528
rect 275278 3516 275284 3528
rect 272576 3488 275284 3516
rect 272576 3476 272582 3488
rect 275278 3476 275284 3488
rect 275336 3476 275342 3528
rect 275741 3519 275799 3525
rect 275741 3485 275753 3519
rect 275787 3516 275799 3519
rect 278041 3519 278099 3525
rect 275787 3488 276796 3516
rect 275787 3485 275799 3488
rect 275741 3479 275799 3485
rect 276768 3448 276796 3488
rect 278041 3485 278053 3519
rect 278087 3516 278099 3519
rect 291930 3516 291936 3528
rect 278087 3488 291936 3516
rect 278087 3485 278099 3488
rect 278041 3479 278099 3485
rect 291930 3476 291936 3488
rect 291988 3476 291994 3528
rect 292482 3476 292488 3528
rect 292540 3516 292546 3528
rect 353754 3516 353760 3528
rect 292540 3488 353760 3516
rect 292540 3476 292546 3488
rect 353754 3476 353760 3488
rect 353812 3476 353818 3528
rect 368382 3476 368388 3528
rect 368440 3516 368446 3528
rect 575014 3516 575020 3528
rect 368440 3488 575020 3516
rect 368440 3476 368446 3488
rect 575014 3476 575020 3488
rect 575072 3476 575078 3528
rect 293126 3448 293132 3460
rect 271800 3420 276704 3448
rect 276768 3420 293132 3448
rect 231946 3380 231952 3392
rect 226444 3352 231952 3380
rect 226337 3343 226395 3349
rect 231946 3340 231952 3352
rect 232004 3340 232010 3392
rect 245562 3340 245568 3392
rect 245620 3380 245626 3392
rect 250530 3380 250536 3392
rect 245620 3352 250536 3380
rect 245620 3340 245626 3352
rect 250530 3340 250536 3352
rect 250588 3340 250594 3392
rect 266998 3340 267004 3392
rect 267056 3380 267062 3392
rect 274082 3380 274088 3392
rect 267056 3352 274088 3380
rect 267056 3340 267062 3352
rect 274082 3340 274088 3352
rect 274140 3340 274146 3392
rect 274174 3340 274180 3392
rect 274232 3380 274238 3392
rect 276676 3380 276704 3420
rect 293126 3408 293132 3420
rect 293184 3408 293190 3460
rect 293862 3408 293868 3460
rect 293920 3448 293926 3460
rect 297269 3451 297327 3457
rect 297269 3448 297281 3451
rect 293920 3420 297281 3448
rect 293920 3408 293926 3420
rect 297269 3417 297281 3420
rect 297315 3417 297327 3451
rect 297269 3411 297327 3417
rect 297358 3408 297364 3460
rect 297416 3448 297422 3460
rect 301406 3448 301412 3460
rect 297416 3420 301412 3448
rect 297416 3408 297422 3420
rect 301406 3408 301412 3420
rect 301464 3408 301470 3460
rect 301593 3451 301651 3457
rect 301593 3417 301605 3451
rect 301639 3448 301651 3451
rect 357342 3448 357348 3460
rect 301639 3420 357348 3448
rect 301639 3417 301651 3420
rect 301593 3411 301651 3417
rect 357342 3408 357348 3420
rect 357400 3408 357406 3460
rect 358078 3408 358084 3460
rect 358136 3448 358142 3460
rect 364981 3451 365039 3457
rect 364981 3448 364993 3451
rect 358136 3420 364993 3448
rect 358136 3408 358142 3420
rect 364981 3417 364993 3420
rect 365027 3417 365039 3451
rect 364981 3411 365039 3417
rect 369762 3408 369768 3460
rect 369820 3448 369826 3460
rect 582190 3448 582196 3460
rect 369820 3420 582196 3448
rect 369820 3408 369826 3420
rect 582190 3408 582196 3420
rect 582248 3408 582254 3460
rect 280062 3380 280068 3392
rect 274232 3352 274496 3380
rect 276676 3352 280068 3380
rect 274232 3340 274238 3352
rect 239398 3312 239404 3324
rect 209924 3216 224908 3244
rect 224972 3284 239404 3312
rect 209924 3204 209930 3216
rect 82688 3148 87736 3176
rect 82688 3136 82694 3148
rect 88518 3136 88524 3188
rect 88576 3176 88582 3188
rect 89622 3176 89628 3188
rect 88576 3148 89628 3176
rect 88576 3136 88582 3148
rect 89622 3136 89628 3148
rect 89680 3136 89686 3188
rect 192478 3176 192484 3188
rect 89732 3148 192484 3176
rect 50522 3068 50528 3120
rect 50580 3108 50586 3120
rect 77938 3108 77944 3120
rect 50580 3080 77944 3108
rect 50580 3068 50586 3080
rect 77938 3068 77944 3080
rect 77996 3068 78002 3120
rect 78033 3111 78091 3117
rect 78033 3077 78045 3111
rect 78079 3108 78091 3111
rect 78953 3111 79011 3117
rect 78953 3108 78965 3111
rect 78079 3080 78965 3108
rect 78079 3077 78091 3080
rect 78033 3071 78091 3077
rect 78953 3077 78965 3080
rect 78999 3077 79011 3111
rect 78953 3071 79011 3077
rect 79042 3068 79048 3120
rect 79100 3108 79106 3120
rect 86037 3111 86095 3117
rect 86037 3108 86049 3111
rect 79100 3080 86049 3108
rect 79100 3068 79106 3080
rect 86037 3077 86049 3080
rect 86083 3077 86095 3111
rect 86037 3071 86095 3077
rect 86126 3068 86132 3120
rect 86184 3108 86190 3120
rect 89732 3108 89760 3148
rect 192478 3136 192484 3148
rect 192536 3136 192542 3188
rect 207474 3136 207480 3188
rect 207532 3176 207538 3188
rect 208302 3176 208308 3188
rect 207532 3148 208308 3176
rect 207532 3136 207538 3148
rect 208302 3136 208308 3148
rect 208360 3136 208366 3188
rect 218146 3136 218152 3188
rect 218204 3176 218210 3188
rect 224972 3176 225000 3284
rect 239398 3272 239404 3284
rect 239456 3272 239462 3324
rect 250346 3272 250352 3324
rect 250404 3312 250410 3324
rect 255590 3312 255596 3324
rect 250404 3284 255596 3312
rect 250404 3272 250410 3284
rect 255590 3272 255596 3284
rect 255648 3272 255654 3324
rect 268838 3272 268844 3324
rect 268896 3312 268902 3324
rect 274361 3315 274419 3321
rect 274361 3312 274373 3315
rect 268896 3284 274373 3312
rect 268896 3272 268902 3284
rect 274361 3281 274373 3284
rect 274407 3281 274419 3315
rect 274468 3312 274496 3352
rect 280062 3340 280068 3352
rect 280120 3340 280126 3392
rect 309778 3380 309784 3392
rect 280172 3352 309784 3380
rect 277210 3312 277216 3324
rect 274468 3284 277216 3312
rect 274361 3275 274419 3281
rect 277210 3272 277216 3284
rect 277268 3272 277274 3324
rect 277302 3272 277308 3324
rect 277360 3312 277366 3324
rect 280172 3312 280200 3352
rect 309778 3340 309784 3352
rect 309836 3340 309842 3392
rect 312538 3340 312544 3392
rect 312596 3380 312602 3392
rect 313366 3380 313372 3392
rect 312596 3352 313372 3380
rect 312596 3340 312602 3352
rect 313366 3340 313372 3352
rect 313424 3340 313430 3392
rect 325234 3380 325240 3392
rect 313476 3352 325240 3380
rect 307386 3312 307392 3324
rect 277360 3284 280200 3312
rect 280264 3284 307392 3312
rect 277360 3272 277366 3284
rect 225049 3247 225107 3253
rect 225049 3213 225061 3247
rect 225095 3244 225107 3247
rect 228729 3247 228787 3253
rect 228729 3244 228741 3247
rect 225095 3216 228741 3244
rect 225095 3213 225107 3216
rect 225049 3207 225107 3213
rect 228729 3213 228741 3216
rect 228775 3213 228787 3247
rect 243538 3244 243544 3256
rect 228729 3207 228787 3213
rect 228836 3216 243544 3244
rect 218204 3148 225000 3176
rect 218204 3136 218210 3148
rect 86184 3080 89760 3108
rect 86184 3068 86190 3080
rect 93302 3068 93308 3120
rect 93360 3108 93366 3120
rect 193858 3108 193864 3120
rect 93360 3080 193864 3108
rect 93360 3068 93366 3080
rect 193858 3068 193864 3080
rect 193916 3068 193922 3120
rect 200390 3068 200396 3120
rect 200448 3108 200454 3120
rect 201402 3108 201408 3120
rect 200448 3080 201408 3108
rect 200448 3068 200454 3080
rect 201402 3068 201408 3080
rect 201460 3068 201466 3120
rect 202690 3068 202696 3120
rect 202748 3108 202754 3120
rect 209038 3108 209044 3120
rect 202748 3080 209044 3108
rect 202748 3068 202754 3080
rect 209038 3068 209044 3080
rect 209096 3068 209102 3120
rect 224126 3068 224132 3120
rect 224184 3108 224190 3120
rect 228836 3108 228864 3216
rect 243538 3204 243544 3216
rect 243596 3204 243602 3256
rect 253842 3204 253848 3256
rect 253900 3244 253906 3256
rect 256878 3244 256884 3256
rect 253900 3216 256884 3244
rect 253900 3204 253906 3216
rect 256878 3204 256884 3216
rect 256936 3204 256942 3256
rect 275922 3204 275928 3256
rect 275980 3244 275986 3256
rect 280264 3244 280292 3284
rect 307386 3272 307392 3284
rect 307444 3272 307450 3324
rect 309686 3272 309692 3324
rect 309744 3312 309750 3324
rect 313476 3312 313504 3352
rect 325234 3340 325240 3352
rect 325292 3340 325298 3392
rect 341518 3340 341524 3392
rect 341576 3380 341582 3392
rect 446582 3380 446588 3392
rect 341576 3352 446588 3380
rect 341576 3340 341582 3352
rect 446582 3340 446588 3352
rect 446640 3340 446646 3392
rect 494054 3340 494060 3392
rect 494112 3380 494118 3392
rect 495342 3380 495348 3392
rect 494112 3352 495348 3380
rect 494112 3340 494118 3352
rect 495342 3340 495348 3352
rect 495400 3340 495406 3392
rect 502334 3340 502340 3392
rect 502392 3380 502398 3392
rect 503622 3380 503628 3392
rect 502392 3352 503628 3380
rect 502392 3340 502398 3352
rect 503622 3340 503628 3352
rect 503680 3340 503686 3392
rect 309744 3284 313504 3312
rect 313553 3315 313611 3321
rect 309744 3272 309750 3284
rect 313553 3281 313565 3315
rect 313599 3312 313611 3315
rect 326430 3312 326436 3324
rect 313599 3284 326436 3312
rect 313599 3281 313611 3284
rect 313553 3275 313611 3281
rect 326430 3272 326436 3284
rect 326488 3272 326494 3324
rect 327718 3272 327724 3324
rect 327776 3312 327782 3324
rect 417970 3312 417976 3324
rect 327776 3284 417976 3312
rect 327776 3272 327782 3284
rect 417970 3272 417976 3284
rect 418028 3272 418034 3324
rect 275980 3216 280292 3244
rect 280341 3247 280399 3253
rect 275980 3204 275986 3216
rect 280341 3213 280353 3247
rect 280387 3244 280399 3247
rect 297177 3247 297235 3253
rect 297177 3244 297189 3247
rect 280387 3216 297189 3244
rect 280387 3213 280399 3216
rect 280341 3207 280399 3213
rect 297177 3213 297189 3216
rect 297223 3213 297235 3247
rect 297177 3207 297235 3213
rect 297453 3247 297511 3253
rect 297453 3213 297465 3247
rect 297499 3244 297511 3247
rect 301593 3247 301651 3253
rect 301593 3244 301605 3247
rect 297499 3216 301605 3244
rect 297499 3213 297511 3216
rect 297453 3207 297511 3213
rect 301593 3213 301605 3216
rect 301639 3213 301651 3247
rect 301593 3207 301651 3213
rect 302970 3204 302976 3256
rect 303028 3244 303034 3256
rect 306190 3244 306196 3256
rect 303028 3216 306196 3244
rect 303028 3204 303034 3216
rect 306190 3204 306196 3216
rect 306248 3204 306254 3256
rect 306285 3247 306343 3253
rect 306285 3213 306297 3247
rect 306331 3244 306343 3247
rect 322842 3244 322848 3256
rect 306331 3216 322848 3244
rect 306331 3213 306343 3216
rect 306285 3207 306343 3213
rect 322842 3204 322848 3216
rect 322900 3204 322906 3256
rect 340138 3204 340144 3256
rect 340196 3244 340202 3256
rect 425146 3244 425152 3256
rect 340196 3216 425152 3244
rect 340196 3204 340202 3216
rect 425146 3204 425152 3216
rect 425204 3204 425210 3256
rect 228910 3136 228916 3188
rect 228968 3176 228974 3188
rect 247678 3176 247684 3188
rect 228968 3148 247684 3176
rect 228968 3136 228974 3148
rect 247678 3136 247684 3148
rect 247736 3136 247742 3188
rect 271782 3136 271788 3188
rect 271840 3176 271846 3188
rect 275741 3179 275799 3185
rect 275741 3176 275753 3179
rect 271840 3148 275753 3176
rect 271840 3136 271846 3148
rect 275741 3145 275753 3148
rect 275787 3145 275799 3179
rect 300302 3176 300308 3188
rect 275741 3139 275799 3145
rect 278148 3148 300308 3176
rect 238018 3108 238024 3120
rect 224184 3080 228864 3108
rect 229848 3080 238024 3108
rect 224184 3068 224190 3080
rect 67913 3043 67971 3049
rect 67913 3009 67925 3043
rect 67959 3040 67971 3043
rect 69569 3043 69627 3049
rect 69569 3040 69581 3043
rect 67959 3012 69581 3040
rect 67959 3009 67971 3012
rect 67913 3003 67971 3009
rect 69569 3009 69581 3012
rect 69615 3009 69627 3043
rect 69569 3003 69627 3009
rect 69753 3043 69811 3049
rect 69753 3009 69765 3043
rect 69799 3040 69811 3043
rect 74537 3043 74595 3049
rect 74537 3040 74549 3043
rect 69799 3012 74549 3040
rect 69799 3009 69811 3012
rect 69753 3003 69811 3009
rect 74537 3009 74549 3012
rect 74583 3009 74595 3043
rect 74537 3003 74595 3009
rect 84105 3043 84163 3049
rect 84105 3009 84117 3043
rect 84151 3040 84163 3043
rect 95513 3043 95571 3049
rect 95513 3040 95525 3043
rect 84151 3012 95525 3040
rect 84151 3009 84163 3012
rect 84105 3003 84163 3009
rect 95513 3009 95525 3012
rect 95559 3009 95571 3043
rect 95513 3003 95571 3009
rect 95694 3000 95700 3052
rect 95752 3040 95758 3052
rect 96522 3040 96528 3052
rect 95752 3012 96528 3040
rect 95752 3000 95758 3012
rect 96522 3000 96528 3012
rect 96580 3000 96586 3052
rect 96890 3000 96896 3052
rect 96948 3040 96954 3052
rect 102594 3040 102600 3052
rect 96948 3012 102600 3040
rect 96948 3000 96954 3012
rect 102594 3000 102600 3012
rect 102652 3000 102658 3052
rect 102778 3000 102784 3052
rect 102836 3040 102842 3052
rect 103422 3040 103428 3052
rect 102836 3012 103428 3040
rect 102836 3000 102842 3012
rect 103422 3000 103428 3012
rect 103480 3000 103486 3052
rect 103974 3000 103980 3052
rect 104032 3040 104038 3052
rect 104802 3040 104808 3052
rect 104032 3012 104808 3040
rect 104032 3000 104038 3012
rect 104802 3000 104808 3012
rect 104860 3000 104866 3052
rect 106366 3000 106372 3052
rect 106424 3040 106430 3052
rect 107562 3040 107568 3052
rect 106424 3012 107568 3040
rect 106424 3000 106430 3012
rect 107562 3000 107568 3012
rect 107620 3000 107626 3052
rect 111150 3000 111156 3052
rect 111208 3040 111214 3052
rect 111702 3040 111708 3052
rect 111208 3012 111708 3040
rect 111208 3000 111214 3012
rect 111702 3000 111708 3012
rect 111760 3000 111766 3052
rect 195330 3040 195336 3052
rect 111812 3012 195336 3040
rect 46934 2932 46940 2984
rect 46992 2972 46998 2984
rect 64877 2975 64935 2981
rect 64877 2972 64889 2975
rect 46992 2944 64889 2972
rect 46992 2932 46998 2944
rect 64877 2941 64889 2944
rect 64923 2941 64935 2975
rect 64877 2935 64935 2941
rect 71866 2932 71872 2984
rect 71924 2972 71930 2984
rect 79321 2975 79379 2981
rect 79321 2972 79333 2975
rect 71924 2944 79333 2972
rect 71924 2932 71930 2944
rect 79321 2941 79333 2944
rect 79367 2941 79379 2975
rect 79321 2935 79379 2941
rect 79413 2975 79471 2981
rect 79413 2941 79425 2975
rect 79459 2972 79471 2975
rect 84838 2972 84844 2984
rect 79459 2944 84844 2972
rect 79459 2941 79471 2944
rect 79413 2935 79471 2941
rect 84838 2932 84844 2944
rect 84896 2932 84902 2984
rect 86037 2975 86095 2981
rect 86037 2941 86049 2975
rect 86083 2972 86095 2975
rect 88978 2972 88984 2984
rect 86083 2944 88984 2972
rect 86083 2941 86095 2944
rect 86037 2935 86095 2941
rect 88978 2932 88984 2944
rect 89036 2932 89042 2984
rect 89714 2932 89720 2984
rect 89772 2972 89778 2984
rect 95878 2972 95884 2984
rect 89772 2944 95884 2972
rect 89772 2932 89778 2944
rect 95878 2932 95884 2944
rect 95936 2932 95942 2984
rect 100478 2932 100484 2984
rect 100536 2972 100542 2984
rect 111812 2972 111840 3012
rect 195330 3000 195336 3012
rect 195388 3000 195394 3052
rect 222930 3000 222936 3052
rect 222988 3040 222994 3052
rect 229738 3040 229744 3052
rect 222988 3012 229744 3040
rect 222988 3000 222994 3012
rect 229738 3000 229744 3012
rect 229796 3000 229802 3052
rect 100536 2944 111840 2972
rect 100536 2932 100542 2944
rect 113542 2932 113548 2984
rect 113600 2972 113606 2984
rect 114462 2972 114468 2984
rect 113600 2944 114468 2972
rect 113600 2932 113606 2944
rect 114462 2932 114468 2944
rect 114520 2932 114526 2984
rect 120626 2932 120632 2984
rect 120684 2972 120690 2984
rect 121362 2972 121368 2984
rect 120684 2944 121368 2972
rect 120684 2932 120690 2944
rect 121362 2932 121368 2944
rect 121420 2932 121426 2984
rect 195238 2972 195244 2984
rect 121564 2944 195244 2972
rect 64782 2864 64788 2916
rect 64840 2904 64846 2916
rect 106918 2904 106924 2916
rect 64840 2876 106924 2904
rect 64840 2864 64846 2876
rect 106918 2864 106924 2876
rect 106976 2864 106982 2916
rect 114738 2864 114744 2916
rect 114796 2904 114802 2916
rect 121457 2907 121515 2913
rect 121457 2904 121469 2907
rect 114796 2876 121469 2904
rect 114796 2864 114802 2876
rect 121457 2873 121469 2876
rect 121503 2873 121515 2907
rect 121457 2867 121515 2873
rect 64877 2839 64935 2845
rect 64877 2805 64889 2839
rect 64923 2836 64935 2839
rect 69661 2839 69719 2845
rect 64923 2808 69612 2836
rect 64923 2805 64935 2808
rect 64877 2799 64935 2805
rect 69584 2768 69612 2808
rect 69661 2805 69673 2839
rect 69707 2836 69719 2839
rect 75178 2836 75184 2848
rect 69707 2808 75184 2836
rect 69707 2805 69719 2808
rect 69661 2799 69719 2805
rect 75178 2796 75184 2808
rect 75236 2796 75242 2848
rect 75454 2796 75460 2848
rect 75512 2836 75518 2848
rect 79321 2839 79379 2845
rect 75512 2808 79272 2836
rect 75512 2796 75518 2808
rect 69753 2771 69811 2777
rect 69753 2768 69765 2771
rect 69584 2740 69765 2768
rect 69753 2737 69765 2740
rect 69799 2737 69811 2771
rect 79244 2768 79272 2808
rect 79321 2805 79333 2839
rect 79367 2836 79379 2839
rect 86218 2836 86224 2848
rect 79367 2808 86224 2836
rect 79367 2805 79379 2808
rect 79321 2799 79379 2805
rect 86218 2796 86224 2808
rect 86276 2796 86282 2848
rect 95513 2839 95571 2845
rect 95513 2805 95525 2839
rect 95559 2836 95571 2839
rect 97258 2836 97264 2848
rect 95559 2808 97264 2836
rect 95559 2805 95571 2808
rect 95513 2799 95571 2805
rect 97258 2796 97264 2808
rect 97316 2796 97322 2848
rect 107562 2796 107568 2848
rect 107620 2836 107626 2848
rect 121564 2836 121592 2944
rect 195238 2932 195244 2944
rect 195296 2932 195302 2984
rect 121641 2907 121699 2913
rect 121641 2873 121653 2907
rect 121687 2904 121699 2907
rect 195422 2904 195428 2916
rect 121687 2876 195428 2904
rect 121687 2873 121699 2876
rect 121641 2867 121699 2873
rect 195422 2864 195428 2876
rect 195480 2864 195486 2916
rect 220538 2864 220544 2916
rect 220596 2904 220602 2916
rect 229848 2904 229876 3080
rect 238018 3068 238024 3080
rect 238076 3068 238082 3120
rect 273162 3068 273168 3120
rect 273220 3108 273226 3120
rect 278148 3108 278176 3148
rect 300302 3136 300308 3148
rect 300360 3136 300366 3188
rect 301498 3136 301504 3188
rect 301556 3176 301562 3188
rect 301556 3148 305132 3176
rect 301556 3136 301562 3148
rect 273220 3080 278176 3108
rect 278317 3111 278375 3117
rect 273220 3068 273226 3080
rect 278317 3077 278329 3111
rect 278363 3108 278375 3111
rect 299106 3108 299112 3120
rect 278363 3080 299112 3108
rect 278363 3077 278375 3080
rect 278317 3071 278375 3077
rect 299106 3068 299112 3080
rect 299164 3068 299170 3120
rect 300118 3068 300124 3120
rect 300176 3108 300182 3120
rect 304994 3108 305000 3120
rect 300176 3080 305000 3108
rect 300176 3068 300182 3080
rect 304994 3068 305000 3080
rect 305052 3068 305058 3120
rect 231302 3000 231308 3052
rect 231360 3040 231366 3052
rect 248598 3040 248604 3052
rect 231360 3012 248604 3040
rect 231360 3000 231366 3012
rect 248598 3000 248604 3012
rect 248656 3000 248662 3052
rect 252646 3000 252652 3052
rect 252704 3040 252710 3052
rect 254578 3040 254584 3052
rect 252704 3012 254584 3040
rect 252704 3000 252710 3012
rect 254578 3000 254584 3012
rect 254636 3000 254642 3052
rect 274542 3000 274548 3052
rect 274600 3040 274606 3052
rect 277857 3043 277915 3049
rect 277857 3040 277869 3043
rect 274600 3012 277869 3040
rect 274600 3000 274606 3012
rect 277857 3009 277869 3012
rect 277903 3009 277915 3043
rect 277857 3003 277915 3009
rect 278225 3043 278283 3049
rect 278225 3009 278237 3043
rect 278271 3040 278283 3043
rect 280341 3043 280399 3049
rect 280341 3040 280353 3043
rect 278271 3012 280353 3040
rect 278271 3009 278283 3012
rect 278225 3003 278283 3009
rect 280341 3009 280353 3012
rect 280387 3009 280399 3043
rect 280341 3003 280399 3009
rect 280430 3000 280436 3052
rect 280488 3040 280494 3052
rect 295518 3040 295524 3052
rect 280488 3012 295524 3040
rect 280488 3000 280494 3012
rect 295518 3000 295524 3012
rect 295576 3000 295582 3052
rect 298738 3000 298744 3052
rect 298796 3040 298802 3052
rect 302602 3040 302608 3052
rect 298796 3012 302608 3040
rect 298796 3000 298802 3012
rect 302602 3000 302608 3012
rect 302660 3000 302666 3052
rect 305104 3040 305132 3148
rect 326338 3136 326344 3188
rect 326396 3176 326402 3188
rect 410886 3176 410892 3188
rect 326396 3148 410892 3176
rect 326396 3136 326402 3148
rect 410886 3136 410892 3148
rect 410944 3136 410950 3188
rect 305638 3068 305644 3120
rect 305696 3108 305702 3120
rect 308309 3111 308367 3117
rect 308309 3108 308321 3111
rect 305696 3080 308321 3108
rect 305696 3068 305702 3080
rect 308309 3077 308321 3080
rect 308355 3077 308367 3111
rect 308309 3071 308367 3077
rect 308398 3068 308404 3120
rect 308456 3108 308462 3120
rect 313553 3111 313611 3117
rect 313553 3108 313565 3111
rect 308456 3080 313565 3108
rect 308456 3068 308462 3080
rect 313553 3077 313565 3080
rect 313599 3077 313611 3111
rect 313553 3071 313611 3077
rect 323578 3068 323584 3120
rect 323636 3108 323642 3120
rect 403710 3108 403716 3120
rect 323636 3080 403716 3108
rect 323636 3068 323642 3080
rect 403710 3068 403716 3080
rect 403768 3068 403774 3120
rect 308582 3040 308588 3052
rect 305104 3012 308588 3040
rect 308582 3000 308588 3012
rect 308640 3000 308646 3052
rect 319438 3000 319444 3052
rect 319496 3040 319502 3052
rect 360930 3040 360936 3052
rect 319496 3012 360936 3040
rect 319496 3000 319502 3012
rect 360930 3000 360936 3012
rect 360988 3000 360994 3052
rect 364981 3043 365039 3049
rect 364981 3009 364993 3043
rect 365027 3040 365039 3043
rect 432322 3040 432328 3052
rect 365027 3012 432328 3040
rect 365027 3009 365039 3012
rect 364981 3003 365039 3009
rect 432322 3000 432328 3012
rect 432380 3000 432386 3052
rect 244918 2972 244924 2984
rect 220596 2876 229876 2904
rect 229940 2944 244924 2972
rect 220596 2864 220602 2876
rect 107620 2808 121592 2836
rect 107620 2796 107626 2808
rect 121822 2796 121828 2848
rect 121880 2836 121886 2848
rect 122742 2836 122748 2848
rect 121880 2808 122748 2836
rect 121880 2796 121886 2808
rect 122742 2796 122748 2808
rect 122800 2796 122806 2848
rect 124214 2796 124220 2848
rect 124272 2836 124278 2848
rect 125502 2836 125508 2848
rect 124272 2808 125508 2836
rect 124272 2796 124278 2808
rect 125502 2796 125508 2808
rect 125560 2796 125566 2848
rect 196618 2836 196624 2848
rect 125612 2808 196624 2836
rect 79505 2771 79563 2777
rect 79505 2768 79517 2771
rect 79244 2740 79517 2768
rect 69753 2731 69811 2737
rect 79505 2737 79517 2740
rect 79551 2737 79563 2771
rect 79505 2731 79563 2737
rect 81345 2771 81403 2777
rect 81345 2737 81357 2771
rect 81391 2768 81403 2771
rect 84105 2771 84163 2777
rect 84105 2768 84117 2771
rect 81391 2740 84117 2768
rect 81391 2737 81403 2740
rect 81345 2731 81403 2737
rect 84105 2737 84117 2740
rect 84151 2737 84163 2771
rect 84105 2731 84163 2737
rect 125410 2728 125416 2780
rect 125468 2768 125474 2780
rect 125612 2768 125640 2808
rect 196618 2796 196624 2808
rect 196676 2796 196682 2848
rect 227714 2796 227720 2848
rect 227772 2836 227778 2848
rect 229940 2836 229968 2944
rect 244918 2932 244924 2944
rect 244976 2932 244982 2984
rect 270218 2932 270224 2984
rect 270276 2972 270282 2984
rect 289538 2972 289544 2984
rect 270276 2944 289544 2972
rect 270276 2932 270282 2944
rect 289538 2932 289544 2944
rect 289596 2932 289602 2984
rect 297177 2975 297235 2981
rect 297177 2941 297189 2975
rect 297223 2972 297235 2975
rect 303798 2972 303804 2984
rect 297223 2944 303804 2972
rect 297223 2941 297235 2944
rect 297177 2935 297235 2941
rect 303798 2932 303804 2944
rect 303856 2932 303862 2984
rect 305730 2932 305736 2984
rect 305788 2972 305794 2984
rect 306285 2975 306343 2981
rect 306285 2972 306297 2975
rect 305788 2944 306297 2972
rect 305788 2932 305794 2944
rect 306285 2941 306297 2944
rect 306331 2941 306343 2975
rect 306285 2935 306343 2941
rect 308309 2975 308367 2981
rect 308309 2941 308321 2975
rect 308355 2972 308367 2975
rect 319254 2972 319260 2984
rect 308355 2944 319260 2972
rect 308355 2941 308367 2944
rect 308309 2935 308367 2941
rect 319254 2932 319260 2944
rect 319312 2932 319318 2984
rect 322198 2932 322204 2984
rect 322256 2972 322262 2984
rect 396626 2972 396632 2984
rect 322256 2944 396632 2972
rect 322256 2932 322262 2944
rect 396626 2932 396632 2944
rect 396684 2932 396690 2984
rect 269022 2864 269028 2916
rect 269080 2904 269086 2916
rect 288342 2904 288348 2916
rect 269080 2876 288348 2904
rect 269080 2864 269086 2876
rect 288342 2864 288348 2876
rect 288400 2864 288406 2916
rect 290458 2864 290464 2916
rect 290516 2904 290522 2916
rect 297910 2904 297916 2916
rect 290516 2876 297916 2904
rect 290516 2864 290522 2876
rect 297910 2864 297916 2876
rect 297968 2864 297974 2916
rect 304258 2864 304264 2916
rect 304316 2904 304322 2916
rect 315758 2904 315764 2916
rect 304316 2876 315764 2904
rect 304316 2864 304322 2876
rect 315758 2864 315764 2876
rect 315816 2864 315822 2916
rect 334618 2864 334624 2916
rect 334676 2904 334682 2916
rect 382274 2904 382280 2916
rect 334676 2876 382280 2904
rect 334676 2864 334682 2876
rect 382274 2864 382280 2876
rect 382332 2864 382338 2916
rect 382366 2864 382372 2916
rect 382424 2904 382430 2916
rect 383562 2904 383568 2916
rect 382424 2876 383568 2904
rect 382424 2864 382430 2876
rect 383562 2864 383568 2876
rect 383620 2864 383626 2916
rect 390554 2864 390560 2916
rect 390612 2904 390618 2916
rect 391842 2904 391848 2916
rect 390612 2876 391848 2904
rect 390612 2864 390618 2876
rect 391842 2864 391848 2876
rect 391900 2864 391906 2916
rect 227772 2808 229968 2836
rect 227772 2796 227778 2808
rect 268930 2796 268936 2848
rect 268988 2836 268994 2848
rect 284754 2836 284760 2848
rect 268988 2808 284760 2836
rect 268988 2796 268994 2808
rect 284754 2796 284760 2808
rect 284812 2796 284818 2848
rect 294322 2836 294328 2848
rect 284864 2808 294328 2836
rect 125468 2740 125640 2768
rect 125468 2728 125474 2740
rect 283558 2728 283564 2780
rect 283616 2768 283622 2780
rect 284864 2768 284892 2808
rect 294322 2796 294328 2808
rect 294380 2796 294386 2848
rect 302878 2796 302884 2848
rect 302936 2836 302942 2848
rect 312170 2836 312176 2848
rect 302936 2808 312176 2836
rect 302936 2796 302942 2808
rect 312170 2796 312176 2808
rect 312228 2796 312234 2848
rect 345750 2796 345756 2848
rect 345808 2836 345814 2848
rect 389450 2836 389456 2848
rect 345808 2808 389456 2836
rect 345808 2796 345814 2808
rect 389450 2796 389456 2808
rect 389508 2796 389514 2848
rect 283616 2740 284892 2768
rect 283616 2728 283622 2740
rect 291838 892 291844 944
rect 291896 932 291902 944
rect 296714 932 296720 944
rect 291896 904 296720 932
rect 291896 892 291902 904
rect 296714 892 296720 904
rect 296772 892 296778 944
rect 367094 484 367100 536
rect 367152 524 367158 536
rect 368014 524 368020 536
rect 367152 496 368020 524
rect 367152 484 367158 496
rect 368014 484 368020 496
rect 368072 484 368078 536
rect 375374 484 375380 536
rect 375432 524 375438 536
rect 376386 524 376392 536
rect 375432 496 376392 524
rect 375432 484 375438 496
rect 376386 484 376392 496
rect 376444 484 376450 536
rect 376754 484 376760 536
rect 376812 524 376818 536
rect 377582 524 377588 536
rect 376812 496 377588 524
rect 376812 484 376818 496
rect 377582 484 377588 496
rect 377640 484 377646 536
rect 383654 484 383660 536
rect 383712 524 383718 536
rect 384666 524 384672 536
rect 383712 496 384672 524
rect 383712 484 383718 496
rect 384666 484 384672 496
rect 384724 484 384730 536
rect 385034 484 385040 536
rect 385092 524 385098 536
rect 385862 524 385868 536
rect 385092 496 385868 524
rect 385092 484 385098 496
rect 385862 484 385868 496
rect 385920 484 385926 536
rect 391934 484 391940 536
rect 391992 524 391998 536
rect 393038 524 393044 536
rect 391992 496 393044 524
rect 391992 484 391998 496
rect 393038 484 393044 496
rect 393096 484 393102 536
rect 463694 484 463700 536
rect 463752 524 463758 536
rect 464430 524 464436 536
rect 463752 496 464436 524
rect 463752 484 463758 496
rect 464430 484 464436 496
rect 464488 484 464494 536
rect 478874 484 478880 536
rect 478932 524 478938 536
rect 479886 524 479892 536
rect 478932 496 479892 524
rect 478932 484 478938 496
rect 479886 484 479892 496
rect 479944 484 479950 536
rect 485866 484 485872 536
rect 485924 524 485930 536
rect 486970 524 486976 536
rect 485924 496 486976 524
rect 485924 484 485930 496
rect 486970 484 486976 496
rect 487028 484 487034 536
rect 487154 484 487160 536
rect 487212 524 487218 536
rect 488166 524 488172 536
rect 487212 496 488172 524
rect 487212 484 487218 496
rect 488166 484 488172 496
rect 488224 484 488230 536
rect 489914 484 489920 536
rect 489972 524 489978 536
rect 490558 524 490564 536
rect 489972 496 490564 524
rect 489972 484 489978 496
rect 490558 484 490564 496
rect 490616 484 490622 536
rect 495434 484 495440 536
rect 495492 524 495498 536
rect 496538 524 496544 536
rect 495492 496 496544 524
rect 495492 484 495498 496
rect 496538 484 496544 496
rect 496596 484 496602 536
rect 496814 484 496820 536
rect 496872 524 496878 536
rect 497734 524 497740 536
rect 496872 496 497740 524
rect 496872 484 496878 496
rect 497734 484 497740 496
rect 497792 484 497798 536
rect 538214 484 538220 536
rect 538272 524 538278 536
rect 539318 524 539324 536
rect 538272 496 539324 524
rect 538272 484 538278 496
rect 539318 484 539324 496
rect 539376 484 539382 536
<< via1 >>
rect 137836 700952 137888 701004
rect 280160 700952 280212 701004
rect 262128 700884 262180 700936
rect 413652 700884 413704 700936
rect 105452 700816 105504 700868
rect 283012 700816 283064 700868
rect 89168 700748 89220 700800
rect 287244 700748 287296 700800
rect 255228 700680 255280 700732
rect 462320 700680 462372 700732
rect 72976 700612 73028 700664
rect 284300 700612 284352 700664
rect 256608 700544 256660 700596
rect 478512 700544 478564 700596
rect 40500 700476 40552 700528
rect 288440 700476 288492 700528
rect 24308 700408 24360 700460
rect 249708 700340 249760 700392
rect 527180 700340 527232 700392
rect 8116 700272 8168 700324
rect 290004 700272 290056 700324
rect 336004 700272 336056 700324
rect 429844 700272 429896 700324
rect 260748 700204 260800 700256
rect 397460 700204 397512 700256
rect 154120 700136 154172 700188
rect 281540 700136 281592 700188
rect 170312 700068 170364 700120
rect 277400 700068 277452 700120
rect 279424 700068 279476 700120
rect 364984 700068 365036 700120
rect 267648 700000 267700 700052
rect 269120 700000 269172 700052
rect 348792 700000 348844 700052
rect 202788 699932 202840 699984
rect 274640 699932 274692 699984
rect 264888 699864 264940 699916
rect 332508 699864 332560 699916
rect 218980 699796 219032 699848
rect 276020 699796 276072 699848
rect 235172 699728 235224 699780
rect 273260 699728 273312 699780
rect 267648 699660 267700 699712
rect 271788 699660 271840 699712
rect 283840 699660 283892 699712
rect 291384 698207 291436 698216
rect 291384 698173 291393 698207
rect 291393 698173 291427 698207
rect 291427 698173 291436 698207
rect 291384 698164 291436 698173
rect 245568 696940 245620 696992
rect 579896 696940 579948 696992
rect 269304 695444 269356 695496
rect 287244 695444 287296 695496
rect 290004 695444 290056 695496
rect 291384 695487 291436 695496
rect 291384 695453 291393 695487
rect 291393 695453 291427 695487
rect 291427 695453 291436 695487
rect 291384 695444 291436 695453
rect 267648 688712 267700 688764
rect 252284 688576 252336 688628
rect 252468 688576 252520 688628
rect 289912 688619 289964 688628
rect 289912 688585 289921 688619
rect 289921 688585 289955 688619
rect 289955 688585 289964 688619
rect 289912 688576 289964 688585
rect 291384 688619 291436 688628
rect 291384 688585 291393 688619
rect 291393 688585 291427 688619
rect 291427 688585 291436 688619
rect 291384 688576 291436 688585
rect 299664 688576 299716 688628
rect 300124 688576 300176 688628
rect 559104 688576 559156 688628
rect 559656 688576 559708 688628
rect 287152 688347 287204 688356
rect 287152 688313 287161 688347
rect 287161 688313 287195 688347
rect 287195 688313 287204 688347
rect 287152 688304 287204 688313
rect 267556 685967 267608 685976
rect 267556 685933 267565 685967
rect 267565 685933 267599 685967
rect 267599 685933 267608 685967
rect 267556 685924 267608 685933
rect 269212 685967 269264 685976
rect 269212 685933 269221 685967
rect 269221 685933 269255 685967
rect 269255 685933 269264 685967
rect 269212 685924 269264 685933
rect 246948 685856 247000 685908
rect 580080 685856 580132 685908
rect 252468 685788 252520 685840
rect 267556 684471 267608 684480
rect 267556 684437 267565 684471
rect 267565 684437 267599 684471
rect 267599 684437 267608 684471
rect 267556 684428 267608 684437
rect 269212 684471 269264 684480
rect 269212 684437 269221 684471
rect 269221 684437 269255 684471
rect 269255 684437 269264 684471
rect 269212 684428 269264 684437
rect 299572 684428 299624 684480
rect 559012 684428 559064 684480
rect 276020 683136 276072 683188
rect 276204 683136 276256 683188
rect 267648 682932 267700 682984
rect 3516 681708 3568 681760
rect 292580 681708 292632 681760
rect 291476 678988 291528 679040
rect 291384 678920 291436 678972
rect 252376 676243 252428 676252
rect 252376 676209 252385 676243
rect 252385 676209 252419 676243
rect 252419 676209 252428 676243
rect 252376 676200 252428 676209
rect 269304 676200 269356 676252
rect 287244 676132 287296 676184
rect 494060 676175 494112 676184
rect 494060 676141 494069 676175
rect 494069 676141 494103 676175
rect 494103 676141 494112 676175
rect 494060 676132 494112 676141
rect 267648 674772 267700 674824
rect 242808 673480 242860 673532
rect 580264 673480 580316 673532
rect 269304 669332 269356 669384
rect 252284 669264 252336 669316
rect 252468 669264 252520 669316
rect 276020 669264 276072 669316
rect 276204 669264 276256 669316
rect 269396 669196 269448 669248
rect 3424 667904 3476 667956
rect 296720 667904 296772 667956
rect 287152 666587 287204 666596
rect 287152 666553 287161 666587
rect 287161 666553 287195 666587
rect 287195 666553 287204 666587
rect 287152 666544 287204 666553
rect 299940 666544 299992 666596
rect 494152 666544 494204 666596
rect 559380 666544 559432 666596
rect 252468 666476 252520 666528
rect 276204 666476 276256 666528
rect 289820 666519 289872 666528
rect 289820 666485 289829 666519
rect 289829 666485 289863 666519
rect 289863 666485 289872 666519
rect 289820 666476 289872 666485
rect 267372 665295 267424 665304
rect 267372 665261 267381 665295
rect 267381 665261 267415 665295
rect 267415 665261 267424 665295
rect 267372 665252 267424 665261
rect 267372 665116 267424 665168
rect 269396 663731 269448 663740
rect 269396 663697 269405 663731
rect 269405 663697 269439 663731
rect 269439 663697 269448 663731
rect 269396 663688 269448 663697
rect 267556 659583 267608 659592
rect 267556 659549 267565 659583
rect 267565 659549 267599 659583
rect 267599 659549 267608 659583
rect 267556 659540 267608 659549
rect 252376 656931 252428 656940
rect 252376 656897 252385 656931
rect 252385 656897 252419 656931
rect 252419 656897 252428 656931
rect 252376 656888 252428 656897
rect 276112 656931 276164 656940
rect 276112 656897 276121 656931
rect 276121 656897 276155 656931
rect 276155 656897 276164 656931
rect 276112 656888 276164 656897
rect 289820 656931 289872 656940
rect 289820 656897 289829 656931
rect 289829 656897 289863 656931
rect 289863 656897 289872 656931
rect 289820 656888 289872 656897
rect 494060 654100 494112 654152
rect 494244 654100 494296 654152
rect 3056 652740 3108 652792
rect 295340 652740 295392 652792
rect 267556 650156 267608 650208
rect 240048 650020 240100 650072
rect 579896 650020 579948 650072
rect 252284 649952 252336 650004
rect 252468 649952 252520 650004
rect 269396 649927 269448 649936
rect 269396 649893 269405 649927
rect 269405 649893 269439 649927
rect 269439 649893 269448 649927
rect 269396 649884 269448 649893
rect 287244 649884 287296 649936
rect 287244 649748 287296 649800
rect 299664 647232 299716 647284
rect 299756 647232 299808 647284
rect 559104 647232 559156 647284
rect 559196 647232 559248 647284
rect 252468 647164 252520 647216
rect 289820 647207 289872 647216
rect 289820 647173 289829 647207
rect 289829 647173 289863 647207
rect 289863 647173 289872 647207
rect 289820 647164 289872 647173
rect 267464 645915 267516 645924
rect 267464 645881 267473 645915
rect 267473 645881 267507 645915
rect 267507 645881 267516 645915
rect 267464 645872 267516 645881
rect 276020 644444 276072 644496
rect 276204 644444 276256 644496
rect 269396 640364 269448 640416
rect 299664 640364 299716 640416
rect 299756 640364 299808 640416
rect 559104 640364 559156 640416
rect 559196 640364 559248 640416
rect 269304 640228 269356 640280
rect 241428 638936 241480 638988
rect 580080 638936 580132 638988
rect 252376 637619 252428 637628
rect 252376 637585 252385 637619
rect 252385 637585 252419 637619
rect 252419 637585 252428 637619
rect 252376 637576 252428 637585
rect 289820 637619 289872 637628
rect 289820 637585 289829 637619
rect 289829 637585 289863 637619
rect 289863 637585 289872 637619
rect 289820 637576 289872 637585
rect 291384 637508 291436 637560
rect 494060 634788 494112 634840
rect 494244 634788 494296 634840
rect 267556 630844 267608 630896
rect 287060 630640 287112 630692
rect 287244 630640 287296 630692
rect 299572 630640 299624 630692
rect 299756 630640 299808 630692
rect 559012 630640 559064 630692
rect 559196 630640 559248 630692
rect 291292 627963 291344 627972
rect 291292 627929 291301 627963
rect 291301 627929 291335 627963
rect 291335 627929 291344 627963
rect 291292 627920 291344 627929
rect 289912 627895 289964 627904
rect 289912 627861 289921 627895
rect 289921 627861 289955 627895
rect 289955 627861 289964 627895
rect 289912 627852 289964 627861
rect 267464 626671 267516 626680
rect 267464 626637 267473 626671
rect 267473 626637 267507 626671
rect 267507 626637 267516 626671
rect 267464 626628 267516 626637
rect 238668 626560 238720 626612
rect 580264 626560 580316 626612
rect 3424 623772 3476 623824
rect 298100 623772 298152 623824
rect 267464 623092 267516 623144
rect 267556 623092 267608 623144
rect 290004 618264 290056 618316
rect 291384 618196 291436 618248
rect 257988 617516 258040 617568
rect 336004 617516 336056 617568
rect 494060 615476 494112 615528
rect 494244 615476 494296 615528
rect 269304 611396 269356 611448
rect 276020 611328 276072 611380
rect 276204 611328 276256 611380
rect 287060 611328 287112 611380
rect 287244 611328 287296 611380
rect 289820 611328 289872 611380
rect 290004 611328 290056 611380
rect 299572 611328 299624 611380
rect 299756 611328 299808 611380
rect 559012 611328 559064 611380
rect 559196 611328 559248 611380
rect 269304 611260 269356 611312
rect 3424 609968 3476 610020
rect 302240 609968 302292 610020
rect 291292 608651 291344 608660
rect 291292 608617 291301 608651
rect 291301 608617 291335 608651
rect 291335 608617 291344 608651
rect 291292 608608 291344 608617
rect 287152 608583 287204 608592
rect 287152 608549 287161 608583
rect 287161 608549 287195 608583
rect 287195 608549 287204 608583
rect 287152 608540 287204 608549
rect 299664 608583 299716 608592
rect 299664 608549 299673 608583
rect 299673 608549 299707 608583
rect 299707 608549 299716 608583
rect 299664 608540 299716 608549
rect 559104 608583 559156 608592
rect 559104 608549 559113 608583
rect 559113 608549 559147 608583
rect 559147 608549 559156 608583
rect 559104 608540 559156 608549
rect 291292 607155 291344 607164
rect 291292 607121 291301 607155
rect 291301 607121 291335 607155
rect 291335 607121 291344 607155
rect 291292 607112 291344 607121
rect 234528 603100 234580 603152
rect 579896 603100 579948 603152
rect 276112 601740 276164 601792
rect 269120 601672 269172 601724
rect 269304 601672 269356 601724
rect 276204 601672 276256 601724
rect 299848 601672 299900 601724
rect 559288 601672 559340 601724
rect 287244 598952 287296 599004
rect 269120 598927 269172 598936
rect 269120 598893 269129 598927
rect 269129 598893 269163 598927
rect 269163 598893 269172 598927
rect 269120 598884 269172 598893
rect 276204 598927 276256 598936
rect 276204 598893 276213 598927
rect 276213 598893 276247 598927
rect 276247 598893 276256 598927
rect 276204 598884 276256 598893
rect 299848 598884 299900 598936
rect 559288 598927 559340 598936
rect 559288 598893 559297 598927
rect 559297 598893 559331 598927
rect 559331 598893 559340 598927
rect 559288 598884 559340 598893
rect 291384 597524 291436 597576
rect 494060 596164 494112 596216
rect 494244 596164 494296 596216
rect 3240 594804 3292 594856
rect 299572 594804 299624 594856
rect 267372 592084 267424 592136
rect 235908 592016 235960 592068
rect 580080 592016 580132 592068
rect 276204 591991 276256 592000
rect 276204 591957 276213 591991
rect 276213 591957 276247 591991
rect 276247 591957 276256 591991
rect 276204 591948 276256 591957
rect 267280 589407 267332 589416
rect 267280 589373 267289 589407
rect 267289 589373 267323 589407
rect 267323 589373 267332 589407
rect 267280 589364 267332 589373
rect 269212 589296 269264 589348
rect 299756 589339 299808 589348
rect 299756 589305 299765 589339
rect 299765 589305 299799 589339
rect 299799 589305 299808 589339
rect 299756 589296 299808 589305
rect 559380 589296 559432 589348
rect 276204 589271 276256 589280
rect 276204 589237 276213 589271
rect 276213 589237 276247 589271
rect 276247 589237 276256 589271
rect 276204 589228 276256 589237
rect 493876 589228 493928 589280
rect 494152 589228 494204 589280
rect 269212 587843 269264 587852
rect 269212 587809 269221 587843
rect 269221 587809 269255 587843
rect 269255 587809 269264 587843
rect 269212 587800 269264 587809
rect 267280 582360 267332 582412
rect 269304 582360 269356 582412
rect 299756 582360 299808 582412
rect 267372 582224 267424 582276
rect 276204 582267 276256 582276
rect 276204 582233 276213 582267
rect 276213 582233 276247 582267
rect 276247 582233 276256 582267
rect 276204 582224 276256 582233
rect 559380 582428 559432 582480
rect 559288 582292 559340 582344
rect 299848 582224 299900 582276
rect 233148 579640 233200 579692
rect 580264 579640 580316 579692
rect 291384 579615 291436 579624
rect 291384 579581 291393 579615
rect 291393 579581 291427 579615
rect 291427 579581 291436 579615
rect 291384 579572 291436 579581
rect 276020 572704 276072 572756
rect 276204 572704 276256 572756
rect 287060 572704 287112 572756
rect 287244 572704 287296 572756
rect 289820 572704 289872 572756
rect 290004 572704 290056 572756
rect 299480 572704 299532 572756
rect 299848 572704 299900 572756
rect 291476 569916 291528 569968
rect 494152 569891 494204 569900
rect 494152 569857 494161 569891
rect 494161 569857 494195 569891
rect 494195 569857 494204 569891
rect 494152 569848 494204 569857
rect 269120 568556 269172 568608
rect 269396 568556 269448 568608
rect 3424 567196 3476 567248
rect 303620 567196 303672 567248
rect 269396 563116 269448 563168
rect 291476 563116 291528 563168
rect 559012 563116 559064 563168
rect 494336 563048 494388 563100
rect 269304 562980 269356 563032
rect 291384 562980 291436 563032
rect 559012 562980 559064 563032
rect 267372 562912 267424 562964
rect 267556 562912 267608 562964
rect 559012 560235 559064 560244
rect 559012 560201 559021 560235
rect 559021 560201 559055 560235
rect 559055 560201 559064 560235
rect 559012 560192 559064 560201
rect 229008 556180 229060 556232
rect 579896 556180 579948 556232
rect 289820 553392 289872 553444
rect 290004 553392 290056 553444
rect 291292 553324 291344 553376
rect 299480 553324 299532 553376
rect 299940 553324 299992 553376
rect 291292 553188 291344 553240
rect 3148 552032 3200 552084
rect 306380 552032 306432 552084
rect 276020 550604 276072 550656
rect 276112 550604 276164 550656
rect 287060 550604 287112 550656
rect 287152 550604 287204 550656
rect 494152 550604 494204 550656
rect 494428 550604 494480 550656
rect 559196 550604 559248 550656
rect 269212 548836 269264 548888
rect 269488 548836 269540 548888
rect 292580 548020 292632 548072
rect 293316 548020 293368 548072
rect 231768 545096 231820 545148
rect 580080 545096 580132 545148
rect 299940 543804 299992 543856
rect 494428 543804 494480 543856
rect 299848 543668 299900 543720
rect 494336 543668 494388 543720
rect 559012 543600 559064 543652
rect 559196 543600 559248 543652
rect 287060 540880 287112 540932
rect 287244 540880 287296 540932
rect 276296 539588 276348 539640
rect 276388 539588 276440 539640
rect 3424 538228 3476 538280
rect 305000 538228 305052 538280
rect 251824 534080 251876 534132
rect 252376 534080 252428 534132
rect 287336 534080 287388 534132
rect 227628 532720 227680 532772
rect 580264 532720 580316 532772
rect 267188 531292 267240 531344
rect 267556 531292 267608 531344
rect 269304 531292 269356 531344
rect 269580 531292 269632 531344
rect 276296 531292 276348 531344
rect 276572 531292 276624 531344
rect 287152 531335 287204 531344
rect 287152 531301 287161 531335
rect 287161 531301 287195 531335
rect 287195 531301 287204 531335
rect 287152 531292 287204 531301
rect 291292 531292 291344 531344
rect 291844 531292 291896 531344
rect 293316 531292 293368 531344
rect 293500 531292 293552 531344
rect 299664 531292 299716 531344
rect 299940 531292 299992 531344
rect 494152 531292 494204 531344
rect 494428 531292 494480 531344
rect 230480 526464 230532 526516
rect 231768 526464 231820 526516
rect 231860 526464 231912 526516
rect 233148 526464 233200 526516
rect 233240 526464 233292 526516
rect 234528 526464 234580 526516
rect 234620 526464 234672 526516
rect 235908 526464 235960 526516
rect 237380 526464 237432 526516
rect 238668 526464 238720 526516
rect 276388 526328 276440 526380
rect 276572 526328 276624 526380
rect 263324 523880 263376 523932
rect 279424 523880 279476 523932
rect 268568 523812 268620 523864
rect 299940 523812 299992 523864
rect 253112 523744 253164 523796
rect 494428 523744 494480 523796
rect 248144 523676 248196 523728
rect 559196 523676 559248 523728
rect 219072 522928 219124 522980
rect 371056 522928 371108 522980
rect 213828 522860 213880 522912
rect 370780 522860 370832 522912
rect 190000 522792 190052 522844
rect 376024 522792 376076 522844
rect 2964 522724 3016 522776
rect 309140 522724 309192 522776
rect 4712 522656 4764 522708
rect 312452 522656 312504 522708
rect 3056 522588 3108 522640
rect 310612 522588 310664 522640
rect 3148 522520 3200 522572
rect 317420 522520 317472 522572
rect 3240 522452 3292 522504
rect 319260 522452 319312 522504
rect 5448 522384 5500 522436
rect 323032 522384 323084 522436
rect 325700 522384 325752 522436
rect 335268 522384 335320 522436
rect 6184 522316 6236 522368
rect 327724 522316 327776 522368
rect 4068 522248 4120 522300
rect 326068 522248 326120 522300
rect 19984 522180 20036 522232
rect 343180 522180 343232 522232
rect 345020 522180 345072 522232
rect 354588 522180 354640 522232
rect 10324 522112 10376 522164
rect 332876 522112 332928 522164
rect 13084 522044 13136 522096
rect 338120 522044 338172 522096
rect 5264 521976 5316 522028
rect 331220 521976 331272 522028
rect 21364 521908 21416 521960
rect 348332 521908 348384 521960
rect 3884 521840 3936 521892
rect 334532 521840 334584 521892
rect 3792 521772 3844 521824
rect 336372 521772 336424 521824
rect 5080 521704 5132 521756
rect 346492 521704 346544 521756
rect 186136 521636 186188 521688
rect 580724 521636 580776 521688
rect 311808 521568 311860 521620
rect 311992 521568 312044 521620
rect 224224 520820 224276 520872
rect 369768 520820 369820 520872
rect 220728 520752 220780 520804
rect 370964 520752 371016 520804
rect 217232 520684 217284 520736
rect 370872 520684 370924 520736
rect 212080 520616 212132 520668
rect 370596 520616 370648 520668
rect 208768 520548 208820 520600
rect 369676 520548 369728 520600
rect 206928 520480 206980 520532
rect 369584 520480 369636 520532
rect 203616 520412 203668 520464
rect 369492 520412 369544 520464
rect 188160 520344 188212 520396
rect 580908 520344 580960 520396
rect 183192 520276 183244 520328
rect 580540 520276 580592 520328
rect 179420 519571 179472 519580
rect 179420 519537 179429 519571
rect 179429 519537 179463 519571
rect 179463 519537 179472 519571
rect 179420 519528 179472 519537
rect 215576 519528 215628 519580
rect 370688 519528 370740 519580
rect 6368 519460 6420 519512
rect 314108 519460 314160 519512
rect 5356 519392 5408 519444
rect 320916 519392 320968 519444
rect 3332 519324 3384 519376
rect 324412 519324 324464 519376
rect 339684 519324 339736 519376
rect 3976 519256 4028 519308
rect 329656 519256 329708 519308
rect 345020 519256 345072 519308
rect 349988 519299 350040 519308
rect 349988 519265 349997 519299
rect 349997 519265 350031 519299
rect 350031 519265 350040 519299
rect 349988 519256 350040 519265
rect 351828 519299 351880 519308
rect 351828 519265 351837 519299
rect 351837 519265 351871 519299
rect 351871 519265 351880 519299
rect 351828 519256 351880 519265
rect 355140 519299 355192 519308
rect 355140 519265 355149 519299
rect 355149 519265 355183 519299
rect 355183 519265 355192 519299
rect 355140 519256 355192 519265
rect 3700 519188 3752 519240
rect 5172 519120 5224 519172
rect 4988 519052 5040 519104
rect 360292 519256 360344 519308
rect 3424 518984 3476 519036
rect 4804 518916 4856 518968
rect 370320 518644 370372 518696
rect 375288 518644 375340 518696
rect 3516 518236 3568 518288
rect 580356 518168 580408 518220
rect 50988 517828 51040 517880
rect 57888 517828 57940 517880
rect 70308 517828 70360 517880
rect 77208 517828 77260 517880
rect 89628 517828 89680 517880
rect 96528 517828 96580 517880
rect 108948 517828 109000 517880
rect 115848 517828 115900 517880
rect 128268 517828 128320 517880
rect 135168 517828 135220 517880
rect 147588 517828 147640 517880
rect 154488 517828 154540 517880
rect 27620 517556 27672 517608
rect 37188 517556 37240 517608
rect 369768 510552 369820 510604
rect 579988 510552 580040 510604
rect 579712 510212 579764 510264
rect 579988 510212 580040 510264
rect 371148 499468 371200 499520
rect 579896 499468 579948 499520
rect 2780 495524 2832 495576
rect 4712 495524 4764 495576
rect 398748 486004 398800 486056
rect 405648 486004 405700 486056
rect 371056 463632 371108 463684
rect 579896 463632 579948 463684
rect 370964 452548 371016 452600
rect 579896 452548 579948 452600
rect 3056 452412 3108 452464
rect 6368 452412 6420 452464
rect 370872 440172 370924 440224
rect 579896 440172 579948 440224
rect 3148 424056 3200 424108
rect 6276 424056 6328 424108
rect 370780 416712 370832 416764
rect 579896 416712 579948 416764
rect 370688 405628 370740 405680
rect 579896 405628 579948 405680
rect 370596 393252 370648 393304
rect 579896 393252 579948 393304
rect 2780 380604 2832 380656
rect 5448 380604 5500 380656
rect 369676 369792 369728 369844
rect 579896 369792 579948 369844
rect 2780 366936 2832 366988
rect 5356 366936 5408 366988
rect 369584 346332 369636 346384
rect 580080 346332 580132 346384
rect 3148 324164 3200 324216
rect 6184 324164 6236 324216
rect 369676 322872 369728 322924
rect 580080 322872 580132 322924
rect 3332 280100 3384 280152
rect 10324 280100 10376 280152
rect 2780 266024 2832 266076
rect 5264 266024 5316 266076
rect 3332 237328 3384 237380
rect 13084 237328 13136 237380
rect 315764 219376 315816 219428
rect 315948 219376 316000 219428
rect 334624 218152 334676 218204
rect 223764 218084 223816 218136
rect 223948 218084 224000 218136
rect 88984 217948 89036 218000
rect 197084 217948 197136 218000
rect 218704 217948 218756 218000
rect 224040 217948 224092 218000
rect 224592 217948 224644 218000
rect 330484 218016 330536 218068
rect 340144 218084 340196 218136
rect 244464 217948 244516 218000
rect 266912 217948 266964 218000
rect 279424 217948 279476 218000
rect 282000 217948 282052 218000
rect 308404 217948 308456 218000
rect 315856 217948 315908 218000
rect 334624 218016 334676 218068
rect 86224 217880 86276 217932
rect 194692 217880 194744 217932
rect 196624 217880 196676 217932
rect 213000 217880 213052 217932
rect 215208 217880 215260 217932
rect 243636 217880 243688 217932
rect 271788 217880 271840 217932
rect 283196 217880 283248 217932
rect 284116 217880 284168 217932
rect 284484 217880 284536 217932
rect 285496 217880 285548 217932
rect 286508 217880 286560 217932
rect 286968 217880 287020 217932
rect 287704 217880 287756 217932
rect 288348 217880 288400 217932
rect 289360 217880 289412 217932
rect 289728 217880 289780 217932
rect 290556 217880 290608 217932
rect 291016 217880 291068 217932
rect 291384 217880 291436 217932
rect 292488 217880 292540 217932
rect 293868 217880 293920 217932
rect 319444 217880 319496 217932
rect 320824 217880 320876 217932
rect 321652 217880 321704 217932
rect 322664 217880 322716 217932
rect 329380 217880 329432 217932
rect 77944 217812 77996 217864
rect 187332 217812 187384 217864
rect 212356 217812 212408 217864
rect 240784 217812 240836 217864
rect 298744 217812 298796 217864
rect 301228 217812 301280 217864
rect 335452 217812 335504 217864
rect 336648 217812 336700 217864
rect 336740 217812 336792 217864
rect 337752 217812 337804 217864
rect 340788 217812 340840 217864
rect 345572 217812 345624 217864
rect 345664 217812 345716 217864
rect 346308 217812 346360 217864
rect 346492 217812 346544 217864
rect 347504 217812 347556 217864
rect 348148 217812 348200 217864
rect 349068 217812 349120 217864
rect 349344 217948 349396 218000
rect 350448 217948 350500 218000
rect 358728 217948 358780 218000
rect 469864 217948 469916 218000
rect 358084 217880 358136 217932
rect 366088 217880 366140 217932
rect 478144 217880 478196 217932
rect 352564 217812 352616 217864
rect 355048 217812 355100 217864
rect 355600 217812 355652 217864
rect 362040 217812 362092 217864
rect 362592 217812 362644 217864
rect 363696 217812 363748 217864
rect 475384 217812 475436 217864
rect 75184 217744 75236 217796
rect 185676 217744 185728 217796
rect 191196 217744 191248 217796
rect 195888 217744 195940 217796
rect 209044 217744 209096 217796
rect 239588 217744 239640 217796
rect 275928 217744 275980 217796
rect 278320 217744 278372 217796
rect 304264 217744 304316 217796
rect 318340 217744 318392 217796
rect 350632 217744 350684 217796
rect 351828 217744 351880 217796
rect 354680 217744 354732 217796
rect 355876 217744 355928 217796
rect 356704 217744 356756 217796
rect 357348 217744 357400 217796
rect 357900 217744 357952 217796
rect 358728 217744 358780 217796
rect 361580 217744 361632 217796
rect 362776 217744 362828 217796
rect 364892 217744 364944 217796
rect 365628 217744 365680 217796
rect 365720 217744 365772 217796
rect 366824 217744 366876 217796
rect 367284 217744 367336 217796
rect 368388 217744 368440 217796
rect 368572 217744 368624 217796
rect 480904 217744 480956 217796
rect 71044 217676 71096 217728
rect 175464 217676 175516 217728
rect 210148 217676 210200 217728
rect 242808 217676 242860 217728
rect 256608 217676 256660 217728
rect 257896 217676 257948 217728
rect 262864 217676 262916 217728
rect 263508 217676 263560 217728
rect 264888 217676 264940 217728
rect 265624 217676 265676 217728
rect 267740 217676 267792 217728
rect 268936 217676 268988 217728
rect 270592 217676 270644 217728
rect 271788 217676 271840 217728
rect 277952 217676 278004 217728
rect 278688 217676 278740 217728
rect 279148 217676 279200 217728
rect 280068 217676 280120 217728
rect 280344 217676 280396 217728
rect 281448 217676 281500 217728
rect 292672 217676 292724 217728
rect 293868 217676 293920 217728
rect 295892 217676 295944 217728
rect 296536 217676 296588 217728
rect 296720 217676 296772 217728
rect 298008 217676 298060 217728
rect 300400 217676 300452 217728
rect 300768 217676 300820 217728
rect 301596 217676 301648 217728
rect 302148 217676 302200 217728
rect 303620 217676 303672 217728
rect 331312 217676 331364 217728
rect 331404 217676 331456 217728
rect 332416 217676 332468 217728
rect 333428 217676 333480 217728
rect 333796 217676 333848 217728
rect 334716 217676 334768 217728
rect 335268 217676 335320 217728
rect 335912 217676 335964 217728
rect 336556 217676 336608 217728
rect 337568 217676 337620 217728
rect 337936 217676 337988 217728
rect 338304 217676 338356 217728
rect 339408 217676 339460 217728
rect 341064 217676 341116 217728
rect 341156 217676 341208 217728
rect 342076 217676 342128 217728
rect 342444 217676 342496 217728
rect 343456 217676 343508 217728
rect 345296 217676 345348 217728
rect 346124 217676 346176 217728
rect 347412 217676 347464 217728
rect 347688 217676 347740 217728
rect 348516 217676 348568 217728
rect 348976 217676 349028 217728
rect 349804 217676 349856 217728
rect 350356 217676 350408 217728
rect 351000 217676 351052 217728
rect 351644 217676 351696 217728
rect 352196 217676 352248 217728
rect 353116 217676 353168 217728
rect 353484 217676 353536 217728
rect 354496 217676 354548 217728
rect 355508 217676 355560 217728
rect 355968 217676 356020 217728
rect 356336 217676 356388 217728
rect 357164 217676 357216 217728
rect 357532 217676 357584 217728
rect 358544 217676 358596 217728
rect 359188 217676 359240 217728
rect 360016 217676 360068 217728
rect 360384 217676 360436 217728
rect 361488 217676 361540 217728
rect 362408 217676 362460 217728
rect 362868 217676 362920 217728
rect 363236 217676 363288 217728
rect 364156 217676 364208 217728
rect 364432 217676 364484 217728
rect 365444 217676 365496 217728
rect 366548 217676 366600 217728
rect 367008 217676 367060 217728
rect 367744 217676 367796 217728
rect 368296 217676 368348 217728
rect 368940 217676 368992 217728
rect 369676 217676 369728 217728
rect 474004 217676 474056 217728
rect 42064 217608 42116 217660
rect 183652 217608 183704 217660
rect 188344 217608 188396 217660
rect 193404 217608 193456 217660
rect 195428 217608 195480 217660
rect 209320 217608 209372 217660
rect 212264 217608 212316 217660
rect 242440 217608 242492 217660
rect 247776 217608 247828 217660
rect 250628 217608 250680 217660
rect 255228 217608 255280 217660
rect 257528 217608 257580 217660
rect 260748 217608 260800 217660
rect 261576 217608 261628 217660
rect 264428 217608 264480 217660
rect 272524 217608 272576 217660
rect 279608 217608 279660 217660
rect 295524 217608 295576 217660
rect 296628 217608 296680 217660
rect 299572 217608 299624 217660
rect 300584 217608 300636 217660
rect 35164 217540 35216 217592
rect 181168 217540 181220 217592
rect 181352 217540 181404 217592
rect 181904 217540 181956 217592
rect 195244 217540 195296 217592
rect 206928 217540 206980 217592
rect 208308 217540 208360 217592
rect 241152 217540 241204 217592
rect 245568 217540 245620 217592
rect 253848 217540 253900 217592
rect 277124 217540 277176 217592
rect 302884 217608 302936 217660
rect 319536 217608 319588 217660
rect 434720 217608 434772 217660
rect 322388 217540 322440 217592
rect 322848 217540 322900 217592
rect 324872 217540 324924 217592
rect 325608 217540 325660 217592
rect 326068 217540 326120 217592
rect 326988 217540 327040 217592
rect 327356 217540 327408 217592
rect 328368 217540 328420 217592
rect 328552 217540 328604 217592
rect 329656 217540 329708 217592
rect 330208 217540 330260 217592
rect 331036 217540 331088 217592
rect 443000 217540 443052 217592
rect 32404 217472 32456 217524
rect 31024 217404 31076 217456
rect 24124 217336 24176 217388
rect 183192 217472 183244 217524
rect 186964 217472 187016 217524
rect 191012 217472 191064 217524
rect 195336 217472 195388 217524
rect 204444 217472 204496 217524
rect 204904 217472 204956 217524
rect 237564 217472 237616 217524
rect 238024 217472 238076 217524
rect 245660 217472 245712 217524
rect 248328 217472 248380 217524
rect 255044 217472 255096 217524
rect 281632 217472 281684 217524
rect 309784 217472 309836 217524
rect 317144 217472 317196 217524
rect 323676 217472 323728 217524
rect 324228 217472 324280 217524
rect 324504 217472 324556 217524
rect 449900 217472 449952 217524
rect 178776 217404 178828 217456
rect 203524 217404 203576 217456
rect 238300 217404 238352 217456
rect 238668 217404 238720 217456
rect 251824 217404 251876 217456
rect 260012 217404 260064 217456
rect 261484 217404 261536 217456
rect 269396 217404 269448 217456
rect 270224 217404 270276 217456
rect 273812 217404 273864 217456
rect 17224 217268 17276 217320
rect 175096 217336 175148 217388
rect 204168 217336 204220 217388
rect 239956 217336 240008 217388
rect 240784 217336 240836 217388
rect 249892 217336 249944 217388
rect 264060 217336 264112 217388
rect 267004 217336 267056 217388
rect 276296 217336 276348 217388
rect 277308 217336 277360 217388
rect 277492 217336 277544 217388
rect 301504 217404 301556 217456
rect 306104 217404 306156 217456
rect 322204 217404 322256 217456
rect 323216 217404 323268 217456
rect 302976 217336 303028 217388
rect 310980 217336 311032 217388
rect 178316 217268 178368 217320
rect 192208 217268 192260 217320
rect 192484 217268 192536 217320
rect 199568 217268 199620 217320
rect 201408 217268 201460 217320
rect 238760 217268 238812 217320
rect 241428 217268 241480 217320
rect 252652 217268 252704 217320
rect 265256 217268 265308 217320
rect 276664 217268 276716 217320
rect 280804 217268 280856 217320
rect 84844 217200 84896 217252
rect 189724 217200 189776 217252
rect 192576 217200 192628 217252
rect 198372 217200 198424 217252
rect 219348 217200 219400 217252
rect 245292 217200 245344 217252
rect 278780 217200 278832 217252
rect 283656 217200 283708 217252
rect 285680 217200 285732 217252
rect 286876 217200 286928 217252
rect 288532 217268 288584 217320
rect 289636 217268 289688 217320
rect 290188 217268 290240 217320
rect 291108 217268 291160 217320
rect 312544 217268 312596 217320
rect 313464 217336 313516 217388
rect 327724 217336 327776 217388
rect 328184 217336 328236 217388
rect 332600 217404 332652 217456
rect 333704 217404 333756 217456
rect 337108 217404 337160 217456
rect 338028 217404 338080 217456
rect 339960 217404 340012 217456
rect 340604 217404 340656 217456
rect 456800 217404 456852 217456
rect 338764 217336 338816 217388
rect 339316 217336 339368 217388
rect 326344 217268 326396 217320
rect 326896 217268 326948 217320
rect 463700 217336 463752 217388
rect 477500 217268 477552 217320
rect 305736 217200 305788 217252
rect 313832 217200 313884 217252
rect 314568 217200 314620 217252
rect 95884 217132 95936 217184
rect 200764 217132 200816 217184
rect 226248 217132 226300 217184
rect 247316 217132 247368 217184
rect 275100 217132 275152 217184
rect 104808 217064 104860 217116
rect 205640 217064 205692 217116
rect 227628 217064 227680 217116
rect 247684 217064 247736 217116
rect 261208 217064 261260 217116
rect 102784 216996 102836 217048
rect 203248 216996 203300 217048
rect 230388 216996 230440 217048
rect 248972 216996 249024 217048
rect 249340 216996 249392 217048
rect 253020 216996 253072 217048
rect 262404 216996 262456 217048
rect 263416 216996 263468 217048
rect 274640 217064 274692 217116
rect 265256 216996 265308 217048
rect 266544 216996 266596 217048
rect 267648 216996 267700 217048
rect 272248 216996 272300 217048
rect 111708 216928 111760 216980
rect 208124 216928 208176 216980
rect 229744 216928 229796 216980
rect 246488 216928 246540 216980
rect 252468 216928 252520 216980
rect 256332 216928 256384 216980
rect 270960 216928 271012 216980
rect 283564 216928 283616 216980
rect 287336 216996 287388 217048
rect 288256 216996 288308 217048
rect 290464 216928 290516 216980
rect 293040 217064 293092 217116
rect 293776 217064 293828 217116
rect 297088 217132 297140 217184
rect 297824 217132 297876 217184
rect 300124 217132 300176 217184
rect 310060 217132 310112 217184
rect 427820 217200 427872 217252
rect 314844 217132 314896 217184
rect 420920 217132 420972 217184
rect 298376 217064 298428 217116
rect 299296 217064 299348 217116
rect 316684 217064 316736 217116
rect 294236 216996 294288 217048
rect 295248 216996 295300 217048
rect 297364 216928 297416 216980
rect 302424 216996 302476 217048
rect 307300 216996 307352 217048
rect 305644 216928 305696 216980
rect 308588 216928 308640 216980
rect 312176 216996 312228 217048
rect 414020 217064 414072 217116
rect 318156 216996 318208 217048
rect 318524 216996 318576 217048
rect 407120 216996 407172 217048
rect 400220 216928 400272 216980
rect 118608 216860 118660 216912
rect 210608 216860 210660 216912
rect 237288 216860 237340 216912
rect 251364 216860 251416 216912
rect 251916 216860 251968 216912
rect 255504 216860 255556 216912
rect 263692 216860 263744 216912
rect 269764 216860 269816 216912
rect 273444 216860 273496 216912
rect 282828 216860 282880 216912
rect 304908 216860 304960 216912
rect 391940 216860 391992 216912
rect 122748 216792 122800 216844
rect 211528 216792 211580 216844
rect 232504 216792 232556 216844
rect 241980 216792 242032 216844
rect 243544 216792 243596 216844
rect 246948 216792 247000 216844
rect 250904 216792 250956 216844
rect 254216 216792 254268 216844
rect 254584 216792 254636 216844
rect 256700 216792 256752 216844
rect 271420 216792 271472 216844
rect 273904 216792 273956 216844
rect 385040 216792 385092 216844
rect 97264 216724 97316 216776
rect 186136 216724 186188 216776
rect 244924 216724 244976 216776
rect 248144 216724 248196 216776
rect 250812 216724 250864 216776
rect 252192 216724 252244 216776
rect 291844 216724 291896 216776
rect 292396 216724 292448 216776
rect 302792 216724 302844 216776
rect 303528 216724 303580 216776
rect 304080 216724 304132 216776
rect 304908 216724 304960 216776
rect 305276 216724 305328 216776
rect 306196 216724 306248 216776
rect 306472 216724 306524 216776
rect 307576 216724 307628 216776
rect 307760 216724 307812 216776
rect 308864 216724 308916 216776
rect 311440 216724 311492 216776
rect 311808 216724 311860 216776
rect 106924 216656 106976 216708
rect 185584 216656 185636 216708
rect 188528 216656 188580 216708
rect 211804 216656 211856 216708
rect 212264 216656 212316 216708
rect 239404 216656 239456 216708
rect 244832 216656 244884 216708
rect 245016 216656 245068 216708
rect 246120 216656 246172 216708
rect 247684 216656 247736 216708
rect 248512 216656 248564 216708
rect 249156 216656 249208 216708
rect 249800 216656 249852 216708
rect 251824 216656 251876 216708
rect 253480 216656 253532 216708
rect 306932 216656 306984 216708
rect 307668 216656 307720 216708
rect 308128 216656 308180 216708
rect 308956 216656 309008 216708
rect 309324 216656 309376 216708
rect 310336 216656 310388 216708
rect 310612 216656 310664 216708
rect 311624 216656 311676 216708
rect 312636 216656 312688 216708
rect 313188 216656 313240 216708
rect 315120 216656 315172 216708
rect 315948 216656 316000 216708
rect 316316 216656 316368 216708
rect 317328 216656 317380 216708
rect 317512 216656 317564 216708
rect 318616 216656 318668 216708
rect 319168 216656 319220 216708
rect 319996 216656 320048 216708
rect 320364 216656 320416 216708
rect 321376 216656 321428 216708
rect 322020 216724 322072 216776
rect 323584 216656 323636 216708
rect 325700 216656 325752 216708
rect 330576 216724 330628 216776
rect 337384 216724 337436 216776
rect 339592 216724 339644 216776
rect 340788 216724 340840 216776
rect 341064 216724 341116 216776
rect 341524 216724 341576 216776
rect 343640 216724 343692 216776
rect 344744 216724 344796 216776
rect 361212 216724 361264 216776
rect 345664 216656 345716 216708
rect 194692 216316 194744 216368
rect 195520 216316 195572 216368
rect 219808 215704 219860 215756
rect 220360 215704 220412 215756
rect 216864 215568 216916 215620
rect 217508 215568 217560 215620
rect 173992 215296 174044 215348
rect 174636 215296 174688 215348
rect 209872 215296 209924 215348
rect 210792 215296 210844 215348
rect 217140 215296 217192 215348
rect 291936 215203 291988 215212
rect 291936 215169 291945 215203
rect 291945 215169 291979 215203
rect 291979 215169 291988 215203
rect 291936 215160 291988 215169
rect 205732 214548 205784 214600
rect 206192 214548 206244 214600
rect 208492 214548 208544 214600
rect 208676 214548 208728 214600
rect 212816 214548 212868 214600
rect 213552 214548 213604 214600
rect 214012 214548 214064 214600
rect 214748 214548 214800 214600
rect 333336 214548 333388 214600
rect 333888 214548 333940 214600
rect 179420 213800 179472 213852
rect 179972 213800 180024 213852
rect 193864 212848 193916 212900
rect 202052 212848 202104 212900
rect 171416 212508 171468 212560
rect 171784 212508 171836 212560
rect 173256 212508 173308 212560
rect 173808 212508 173860 212560
rect 177304 212508 177356 212560
rect 177948 212508 178000 212560
rect 178868 212508 178920 212560
rect 179144 212508 179196 212560
rect 180156 212551 180208 212560
rect 180156 212517 180165 212551
rect 180165 212517 180199 212551
rect 180199 212517 180208 212551
rect 180156 212508 180208 212517
rect 184020 212508 184072 212560
rect 184480 212508 184532 212560
rect 189356 212508 189408 212560
rect 190184 212508 190236 212560
rect 192392 212508 192444 212560
rect 192668 212508 192720 212560
rect 200856 212508 200908 212560
rect 201224 212508 201276 212560
rect 201868 212508 201920 212560
rect 202420 212508 202472 212560
rect 203432 212508 203484 212560
rect 203616 212508 203668 212560
rect 212356 212551 212408 212560
rect 212356 212517 212365 212551
rect 212365 212517 212399 212551
rect 212399 212517 212408 212551
rect 212356 212508 212408 212517
rect 216956 212551 217008 212560
rect 216956 212517 216965 212551
rect 216965 212517 216999 212551
rect 216999 212517 217008 212551
rect 216956 212508 217008 212517
rect 236276 212508 236328 212560
rect 236736 212508 236788 212560
rect 283748 212508 283800 212560
rect 284024 212508 284076 212560
rect 284852 212508 284904 212560
rect 285312 212508 285364 212560
rect 286140 212508 286192 212560
rect 286600 212508 286652 212560
rect 288992 212508 289044 212560
rect 289360 212508 289412 212560
rect 294696 212508 294748 212560
rect 295064 212508 295116 212560
rect 299940 212508 299992 212560
rect 300492 212508 300544 212560
rect 360752 212508 360804 212560
rect 361304 212508 361356 212560
rect 211896 212483 211948 212492
rect 211896 212449 211905 212483
rect 211905 212449 211939 212483
rect 211939 212449 211948 212483
rect 211896 212440 211948 212449
rect 261944 211896 261996 211948
rect 266544 211896 266596 211948
rect 260380 211216 260432 211268
rect 262588 211216 262640 211268
rect 259552 211148 259604 211200
rect 261116 211148 261168 211200
rect 217048 211123 217100 211132
rect 217048 211089 217057 211123
rect 217057 211089 217091 211123
rect 217091 211089 217100 211123
rect 217048 211080 217100 211089
rect 262588 211123 262640 211132
rect 262588 211089 262597 211123
rect 262597 211089 262631 211123
rect 262631 211089 262640 211123
rect 262588 211080 262640 211089
rect 266544 211080 266596 211132
rect 266728 211080 266780 211132
rect 283840 211080 283892 211132
rect 284024 211080 284076 211132
rect 328092 211123 328144 211132
rect 328092 211089 328101 211123
rect 328101 211089 328135 211123
rect 328135 211089 328144 211123
rect 328092 211080 328144 211089
rect 341800 211080 341852 211132
rect 341984 211080 342036 211132
rect 343272 211123 343324 211132
rect 343272 211089 343281 211123
rect 343281 211089 343315 211123
rect 343315 211089 343324 211123
rect 343272 211080 343324 211089
rect 344560 211123 344612 211132
rect 344560 211089 344569 211123
rect 344569 211089 344603 211123
rect 344603 211089 344612 211123
rect 344560 211080 344612 211089
rect 354128 211080 354180 211132
rect 354220 211080 354272 211132
rect 355416 211080 355468 211132
rect 355600 211080 355652 211132
rect 194692 210876 194744 210928
rect 195152 210876 195204 210928
rect 169944 210468 169996 210520
rect 170680 210468 170732 210520
rect 220912 210468 220964 210520
rect 221740 210468 221792 210520
rect 169852 210400 169904 210452
rect 170312 210400 170364 210452
rect 175372 210400 175424 210452
rect 176016 210400 176068 210452
rect 179512 210400 179564 210452
rect 180064 210400 180116 210452
rect 180892 210400 180944 210452
rect 181260 210400 181312 210452
rect 186412 210400 186464 210452
rect 186596 210400 186648 210452
rect 187976 210400 188028 210452
rect 188620 210400 188672 210452
rect 192024 210400 192076 210452
rect 192760 210400 192812 210452
rect 193312 210400 193364 210452
rect 193956 210400 194008 210452
rect 201684 210400 201736 210452
rect 202512 210400 202564 210452
rect 202972 210400 203024 210452
rect 203708 210400 203760 210452
rect 204352 210400 204404 210452
rect 204996 210400 205048 210452
rect 215392 210400 215444 210452
rect 216036 210400 216088 210452
rect 218060 210400 218112 210452
rect 218796 210400 218848 210452
rect 221004 210400 221056 210452
rect 221372 210400 221424 210452
rect 222292 210400 222344 210452
rect 222476 210400 222528 210452
rect 224960 210400 225012 210452
rect 225788 210400 225840 210452
rect 226340 210400 226392 210452
rect 227076 210400 227128 210452
rect 227904 210400 227956 210452
rect 228640 210400 228692 210452
rect 229100 210400 229152 210452
rect 229468 210400 229520 210452
rect 230480 210400 230532 210452
rect 231124 210400 231176 210452
rect 231860 210400 231912 210452
rect 232780 210400 232832 210452
rect 233332 210400 233384 210452
rect 233976 210400 234028 210452
rect 236000 210400 236052 210452
rect 236828 210400 236880 210452
rect 242992 210400 243044 210452
rect 243820 210400 243872 210452
rect 270132 210400 270184 210452
rect 270316 210400 270368 210452
rect 346952 210400 347004 210452
rect 347688 210400 347740 210452
rect 234620 210332 234672 210384
rect 234896 210332 234948 210384
rect 207112 209788 207164 209840
rect 207388 209788 207440 209840
rect 225144 209720 225196 209772
rect 225420 209720 225472 209772
rect 275836 209720 275888 209772
rect 276112 209720 276164 209772
rect 329380 209763 329432 209772
rect 329380 209729 329389 209763
rect 329389 209729 329423 209763
rect 329423 209729 329432 209763
rect 329380 209720 329432 209729
rect 223580 208496 223632 208548
rect 224132 208496 224184 208548
rect 183836 208360 183888 208412
rect 184572 208360 184624 208412
rect 198832 208292 198884 208344
rect 199660 208292 199712 208344
rect 258264 207723 258316 207732
rect 258264 207689 258273 207723
rect 258273 207689 258307 207723
rect 258307 207689 258316 207723
rect 258264 207680 258316 207689
rect 229192 207000 229244 207052
rect 229836 207000 229888 207052
rect 222200 206456 222252 206508
rect 222936 206456 222988 206508
rect 230664 205844 230716 205896
rect 230848 205844 230900 205896
rect 197452 205708 197504 205760
rect 197636 205708 197688 205760
rect 234804 205708 234856 205760
rect 182272 205640 182324 205692
rect 182548 205640 182600 205692
rect 196072 205640 196124 205692
rect 196348 205640 196400 205692
rect 219808 205683 219860 205692
rect 219808 205649 219817 205683
rect 219817 205649 219851 205683
rect 219851 205649 219860 205683
rect 219808 205640 219860 205649
rect 286600 205640 286652 205692
rect 315856 205683 315908 205692
rect 315856 205649 315865 205683
rect 315865 205649 315899 205683
rect 315899 205649 315908 205683
rect 315856 205640 315908 205649
rect 171416 205572 171468 205624
rect 171600 205572 171652 205624
rect 234804 205572 234856 205624
rect 236276 205572 236328 205624
rect 236460 205572 236512 205624
rect 262588 205615 262640 205624
rect 262588 205581 262597 205615
rect 262597 205581 262631 205615
rect 262631 205581 262640 205615
rect 262588 205572 262640 205581
rect 282644 205504 282696 205556
rect 282828 205504 282880 205556
rect 328184 205572 328236 205624
rect 343272 205615 343324 205624
rect 343272 205581 343281 205615
rect 343281 205581 343315 205615
rect 343315 205581 343324 205615
rect 343272 205572 343324 205581
rect 344560 205615 344612 205624
rect 344560 205581 344569 205615
rect 344569 205581 344603 205615
rect 344603 205581 344612 205615
rect 344560 205572 344612 205581
rect 286692 205504 286744 205556
rect 173348 202852 173400 202904
rect 173440 202852 173492 202904
rect 211988 202852 212040 202904
rect 212172 202852 212224 202904
rect 212448 202852 212500 202904
rect 219808 202895 219860 202904
rect 219808 202861 219817 202895
rect 219817 202861 219851 202895
rect 219851 202861 219860 202895
rect 219808 202852 219860 202861
rect 232136 202852 232188 202904
rect 232320 202852 232372 202904
rect 258356 202852 258408 202904
rect 289176 202852 289228 202904
rect 289452 202852 289504 202904
rect 315856 202895 315908 202904
rect 315856 202861 315865 202895
rect 315865 202861 315899 202895
rect 315899 202861 315908 202895
rect 315856 202852 315908 202861
rect 352840 202852 352892 202904
rect 353024 202852 353076 202904
rect 217140 201492 217192 201544
rect 184112 201424 184164 201476
rect 184296 201424 184348 201476
rect 192392 201424 192444 201476
rect 282828 201467 282880 201476
rect 282828 201433 282837 201467
rect 282837 201433 282871 201467
rect 282871 201433 282880 201467
rect 282828 201424 282880 201433
rect 329472 201424 329524 201476
rect 362592 201424 362644 201476
rect 229468 200064 229520 200116
rect 229560 200064 229612 200116
rect 230848 200064 230900 200116
rect 231400 200064 231452 200116
rect 277216 200107 277268 200116
rect 277216 200073 277225 200107
rect 277225 200073 277259 200107
rect 277259 200073 277268 200107
rect 277216 200064 277268 200073
rect 232136 198092 232188 198144
rect 232044 198024 232096 198076
rect 234988 198024 235040 198076
rect 235632 198024 235684 198076
rect 234804 197956 234856 198008
rect 235172 197956 235224 198008
rect 262404 196596 262456 196648
rect 262680 196596 262732 196648
rect 315856 196052 315908 196104
rect 171508 196027 171560 196036
rect 171508 195993 171517 196027
rect 171517 195993 171551 196027
rect 171551 195993 171560 196027
rect 171508 195984 171560 195993
rect 219808 195984 219860 196036
rect 219716 195916 219768 195968
rect 275836 195236 275888 195288
rect 276112 195236 276164 195288
rect 180064 195168 180116 195220
rect 180156 195168 180208 195220
rect 3148 194488 3200 194540
rect 19984 194488 20036 194540
rect 171508 193239 171560 193248
rect 171508 193205 171517 193239
rect 171517 193205 171551 193239
rect 171551 193205 171560 193239
rect 171508 193196 171560 193205
rect 173164 193196 173216 193248
rect 173532 193196 173584 193248
rect 203248 193196 203300 193248
rect 203340 193196 203392 193248
rect 216680 193196 216732 193248
rect 216956 193196 217008 193248
rect 286508 193196 286560 193248
rect 286692 193196 286744 193248
rect 289268 193196 289320 193248
rect 289452 193196 289504 193248
rect 192116 193171 192168 193180
rect 192116 193137 192125 193171
rect 192125 193137 192159 193171
rect 192159 193137 192168 193171
rect 192116 193128 192168 193137
rect 217140 193128 217192 193180
rect 217232 193128 217284 193180
rect 282828 193171 282880 193180
rect 282828 193137 282837 193171
rect 282837 193137 282871 193171
rect 282871 193137 282880 193171
rect 282828 193128 282880 193137
rect 328276 193060 328328 193112
rect 315764 191879 315816 191888
rect 315764 191845 315773 191879
rect 315773 191845 315807 191879
rect 315807 191845 315816 191879
rect 315764 191836 315816 191845
rect 362500 191879 362552 191888
rect 362500 191845 362509 191879
rect 362509 191845 362543 191879
rect 362543 191845 362552 191879
rect 362500 191836 362552 191845
rect 262496 191811 262548 191820
rect 262496 191777 262505 191811
rect 262505 191777 262539 191811
rect 262539 191777 262548 191811
rect 262496 191768 262548 191777
rect 283840 191768 283892 191820
rect 284024 191768 284076 191820
rect 329564 191811 329616 191820
rect 329564 191777 329573 191811
rect 329573 191777 329607 191811
rect 329607 191777 329616 191811
rect 329564 191768 329616 191777
rect 342996 191768 343048 191820
rect 343180 191768 343232 191820
rect 354220 191811 354272 191820
rect 354220 191777 354229 191811
rect 354229 191777 354263 191811
rect 354263 191777 354272 191811
rect 354220 191768 354272 191777
rect 355416 191768 355468 191820
rect 355508 191768 355560 191820
rect 315764 191700 315816 191752
rect 230572 191088 230624 191140
rect 230756 191088 230808 191140
rect 225236 190408 225288 190460
rect 225420 190408 225472 190460
rect 270132 189864 270184 189916
rect 270316 189864 270368 189916
rect 180064 188980 180116 189032
rect 178868 187756 178920 187808
rect 178224 187688 178276 187740
rect 178224 186396 178276 186448
rect 181168 186328 181220 186380
rect 182180 186371 182232 186380
rect 182180 186337 182189 186371
rect 182189 186337 182223 186371
rect 182223 186337 182232 186371
rect 182180 186328 182232 186337
rect 189448 186328 189500 186380
rect 223948 186328 224000 186380
rect 178132 186260 178184 186312
rect 181076 186260 181128 186312
rect 189540 186192 189592 186244
rect 231032 186396 231084 186448
rect 230940 186260 230992 186312
rect 262496 186303 262548 186312
rect 262496 186269 262505 186303
rect 262505 186269 262539 186303
rect 262539 186269 262548 186303
rect 262496 186260 262548 186269
rect 328184 186303 328236 186312
rect 328184 186269 328193 186303
rect 328193 186269 328227 186303
rect 328227 186269 328236 186303
rect 328184 186260 328236 186269
rect 224040 186192 224092 186244
rect 184020 183608 184072 183660
rect 184112 183608 184164 183660
rect 275836 183608 275888 183660
rect 192116 183540 192168 183592
rect 192208 183540 192260 183592
rect 232136 183540 232188 183592
rect 232228 183540 232280 183592
rect 234988 183540 235040 183592
rect 235080 183540 235132 183592
rect 286692 183608 286744 183660
rect 344376 183608 344428 183660
rect 344560 183608 344612 183660
rect 277216 183583 277268 183592
rect 277216 183549 277225 183583
rect 277225 183549 277259 183583
rect 277259 183549 277268 183583
rect 277216 183540 277268 183549
rect 282736 183540 282788 183592
rect 282920 183540 282972 183592
rect 286600 183540 286652 183592
rect 289268 183540 289320 183592
rect 289452 183540 289504 183592
rect 291660 183540 291712 183592
rect 291936 183540 291988 183592
rect 275836 183472 275888 183524
rect 354220 183515 354272 183524
rect 354220 183481 354229 183515
rect 354229 183481 354263 183515
rect 354263 183481 354272 183515
rect 354220 183472 354272 183481
rect 182180 182223 182232 182232
rect 182180 182189 182189 182223
rect 182189 182189 182223 182223
rect 182223 182189 182232 182223
rect 315672 182223 315724 182232
rect 182180 182180 182232 182189
rect 315672 182189 315681 182223
rect 315681 182189 315715 182223
rect 315715 182189 315724 182223
rect 315672 182180 315724 182189
rect 184112 182112 184164 182164
rect 184204 182112 184256 182164
rect 192208 182155 192260 182164
rect 192208 182121 192217 182155
rect 192217 182121 192251 182155
rect 192251 182121 192260 182155
rect 192208 182112 192260 182121
rect 224040 182155 224092 182164
rect 224040 182121 224049 182155
rect 224049 182121 224083 182155
rect 224083 182121 224092 182155
rect 224040 182112 224092 182121
rect 228272 182112 228324 182164
rect 228364 182112 228416 182164
rect 229284 182112 229336 182164
rect 229468 182112 229520 182164
rect 230940 182112 230992 182164
rect 231032 182112 231084 182164
rect 236276 182112 236328 182164
rect 236460 182112 236512 182164
rect 261116 182112 261168 182164
rect 261300 182112 261352 182164
rect 277216 182112 277268 182164
rect 282828 182112 282880 182164
rect 282920 182112 282972 182164
rect 285220 182155 285272 182164
rect 285220 182121 285229 182155
rect 285229 182121 285263 182155
rect 285263 182121 285272 182155
rect 285220 182112 285272 182121
rect 354312 182155 354364 182164
rect 354312 182121 354321 182155
rect 354321 182121 354355 182155
rect 354355 182121 354364 182155
rect 354312 182112 354364 182121
rect 355600 182155 355652 182164
rect 355600 182121 355609 182155
rect 355609 182121 355643 182155
rect 355643 182121 355652 182155
rect 355600 182112 355652 182121
rect 360936 182112 360988 182164
rect 361212 182112 361264 182164
rect 362592 182112 362644 182164
rect 262588 182087 262640 182096
rect 262588 182053 262597 182087
rect 262597 182053 262631 182087
rect 262631 182053 262640 182087
rect 262588 182044 262640 182053
rect 182180 182019 182232 182028
rect 182180 181985 182189 182019
rect 182189 181985 182223 182019
rect 182223 181985 182232 182019
rect 182180 181976 182232 181985
rect 329380 181568 329432 181620
rect 230572 181432 230624 181484
rect 230756 181432 230808 181484
rect 270132 181432 270184 181484
rect 270316 181432 270368 181484
rect 217324 180795 217376 180804
rect 217324 180761 217333 180795
rect 217333 180761 217367 180795
rect 217367 180761 217376 180795
rect 217324 180752 217376 180761
rect 275836 180795 275888 180804
rect 275836 180761 275845 180795
rect 275845 180761 275879 180795
rect 275879 180761 275888 180795
rect 275836 180752 275888 180761
rect 179972 179435 180024 179444
rect 179972 179401 179981 179435
rect 179981 179401 180015 179435
rect 180015 179401 180024 179435
rect 179972 179392 180024 179401
rect 177120 179324 177172 179376
rect 181076 179367 181128 179376
rect 181076 179333 181085 179367
rect 181085 179333 181119 179367
rect 181119 179333 181128 179367
rect 181076 179324 181128 179333
rect 291936 176740 291988 176792
rect 211712 176672 211764 176724
rect 211988 176672 212040 176724
rect 344560 176604 344612 176656
rect 355600 176647 355652 176656
rect 355600 176613 355609 176647
rect 355609 176613 355643 176647
rect 355643 176613 355652 176647
rect 355600 176604 355652 176613
rect 182272 176536 182324 176588
rect 291936 176536 291988 176588
rect 344468 176536 344520 176588
rect 354404 176536 354456 176588
rect 192208 176103 192260 176112
rect 192208 176069 192217 176103
rect 192217 176069 192251 176103
rect 192251 176069 192260 176103
rect 192208 176060 192260 176069
rect 232136 173952 232188 174004
rect 232228 173952 232280 174004
rect 173072 173884 173124 173936
rect 173164 173884 173216 173936
rect 216680 173884 216732 173936
rect 216956 173884 217008 173936
rect 219808 173884 219860 173936
rect 219992 173884 220044 173936
rect 286508 173884 286560 173936
rect 289268 173884 289320 173936
rect 289452 173884 289504 173936
rect 329380 173884 329432 173936
rect 329564 173884 329616 173936
rect 286600 173748 286652 173800
rect 177120 173136 177172 173188
rect 189448 172524 189500 172576
rect 189540 172524 189592 172576
rect 194968 172524 195020 172576
rect 195060 172524 195112 172576
rect 224040 172567 224092 172576
rect 224040 172533 224049 172567
rect 224049 172533 224083 172567
rect 224083 172533 224092 172567
rect 224040 172524 224092 172533
rect 262588 172567 262640 172576
rect 262588 172533 262597 172567
rect 262597 172533 262631 172567
rect 262631 172533 262640 172567
rect 262588 172524 262640 172533
rect 277124 172567 277176 172576
rect 277124 172533 277133 172567
rect 277133 172533 277167 172567
rect 277167 172533 277176 172567
rect 277124 172524 277176 172533
rect 225420 172499 225472 172508
rect 225420 172465 225429 172499
rect 225429 172465 225463 172499
rect 225463 172465 225472 172499
rect 225420 172456 225472 172465
rect 229376 172499 229428 172508
rect 229376 172465 229385 172499
rect 229385 172465 229419 172499
rect 229419 172465 229428 172499
rect 229376 172456 229428 172465
rect 283840 172456 283892 172508
rect 284024 172456 284076 172508
rect 345480 172456 345532 172508
rect 345664 172456 345716 172508
rect 361120 172456 361172 172508
rect 361396 172456 361448 172508
rect 362316 171164 362368 171216
rect 203156 171096 203208 171148
rect 203248 171096 203300 171148
rect 217416 171096 217468 171148
rect 275928 171096 275980 171148
rect 182272 171028 182324 171080
rect 211712 171028 211764 171080
rect 236368 171071 236420 171080
rect 236368 171037 236377 171071
rect 236377 171037 236411 171071
rect 236411 171037 236420 171071
rect 236368 171028 236420 171037
rect 362408 171071 362460 171080
rect 362408 171037 362417 171071
rect 362417 171037 362451 171071
rect 362451 171037 362460 171071
rect 362408 171028 362460 171037
rect 376024 171028 376076 171080
rect 580172 171028 580224 171080
rect 270132 170552 270184 170604
rect 270316 170552 270368 170604
rect 181352 169736 181404 169788
rect 343272 169668 343324 169720
rect 343364 169668 343416 169720
rect 318524 169124 318576 169176
rect 328000 169056 328052 169108
rect 328184 169056 328236 169108
rect 329288 169056 329340 169108
rect 329472 169056 329524 169108
rect 177120 168351 177172 168360
rect 177120 168317 177129 168351
rect 177129 168317 177163 168351
rect 177163 168317 177172 168351
rect 177120 168308 177172 168317
rect 344652 167492 344704 167544
rect 232136 167084 232188 167136
rect 258172 167016 258224 167068
rect 258356 167016 258408 167068
rect 232136 166948 232188 167000
rect 273076 167084 273128 167136
rect 317052 167016 317104 167068
rect 355692 167016 355744 167068
rect 317144 166948 317196 167000
rect 272984 166880 273036 166932
rect 285312 166880 285364 166932
rect 2780 165452 2832 165504
rect 5172 165452 5224 165504
rect 217232 164228 217284 164280
rect 217416 164228 217468 164280
rect 235264 164228 235316 164280
rect 235356 164228 235408 164280
rect 315672 164228 315724 164280
rect 315764 164228 315816 164280
rect 318432 164271 318484 164280
rect 318432 164237 318441 164271
rect 318441 164237 318475 164271
rect 318475 164237 318484 164271
rect 318432 164228 318484 164237
rect 354312 164228 354364 164280
rect 354404 164228 354456 164280
rect 355600 164271 355652 164280
rect 355600 164237 355609 164271
rect 355609 164237 355643 164271
rect 355643 164237 355652 164271
rect 355600 164228 355652 164237
rect 171416 164160 171468 164212
rect 171600 164160 171652 164212
rect 173072 164160 173124 164212
rect 173256 164160 173308 164212
rect 184020 164160 184072 164212
rect 184112 164160 184164 164212
rect 189356 164160 189408 164212
rect 189448 164160 189500 164212
rect 212448 164203 212500 164212
rect 212448 164169 212457 164203
rect 212457 164169 212491 164203
rect 212491 164169 212500 164203
rect 212448 164160 212500 164169
rect 229376 164203 229428 164212
rect 229376 164169 229385 164203
rect 229385 164169 229419 164203
rect 229419 164169 229428 164203
rect 229376 164160 229428 164169
rect 235080 164160 235132 164212
rect 258264 164203 258316 164212
rect 258264 164169 258273 164203
rect 258273 164169 258307 164203
rect 258307 164169 258316 164203
rect 258264 164160 258316 164169
rect 262312 164160 262364 164212
rect 262496 164160 262548 164212
rect 286600 164160 286652 164212
rect 286692 164160 286744 164212
rect 289360 164160 289412 164212
rect 289452 164160 289504 164212
rect 235172 164092 235224 164144
rect 344560 162911 344612 162920
rect 344560 162877 344569 162911
rect 344569 162877 344603 162911
rect 344603 162877 344612 162911
rect 344560 162868 344612 162877
rect 229468 162800 229520 162852
rect 261116 162843 261168 162852
rect 261116 162809 261125 162843
rect 261125 162809 261159 162843
rect 261159 162809 261168 162843
rect 261116 162800 261168 162809
rect 275836 162800 275888 162852
rect 275928 162800 275980 162852
rect 282644 162800 282696 162852
rect 282828 162800 282880 162852
rect 286692 162843 286744 162852
rect 286692 162809 286701 162843
rect 286701 162809 286735 162843
rect 286735 162809 286744 162843
rect 286692 162800 286744 162809
rect 289268 162800 289320 162852
rect 289452 162800 289504 162852
rect 317144 162843 317196 162852
rect 317144 162809 317153 162843
rect 317153 162809 317187 162843
rect 317187 162809 317196 162843
rect 317144 162800 317196 162809
rect 318432 162843 318484 162852
rect 318432 162809 318441 162843
rect 318441 162809 318475 162843
rect 318475 162809 318484 162843
rect 318432 162800 318484 162809
rect 341984 162843 342036 162852
rect 341984 162809 341993 162843
rect 341993 162809 342027 162843
rect 342027 162809 342036 162843
rect 341984 162800 342036 162809
rect 354312 162843 354364 162852
rect 354312 162809 354321 162843
rect 354321 162809 354355 162843
rect 354355 162809 354364 162843
rect 354312 162800 354364 162809
rect 355600 162800 355652 162852
rect 225420 162707 225472 162716
rect 225420 162673 225429 162707
rect 225429 162673 225463 162707
rect 225463 162673 225472 162707
rect 225420 162664 225472 162673
rect 270132 162120 270184 162172
rect 270316 162120 270368 162172
rect 182180 161483 182232 161492
rect 182180 161449 182189 161483
rect 182189 161449 182223 161483
rect 182223 161449 182232 161483
rect 182180 161440 182232 161449
rect 362408 161483 362460 161492
rect 362408 161449 362417 161483
rect 362417 161449 362451 161483
rect 362451 161449 362460 161483
rect 362408 161440 362460 161449
rect 181076 161415 181128 161424
rect 181076 161381 181085 161415
rect 181085 161381 181119 161415
rect 181119 161381 181128 161415
rect 181076 161372 181128 161381
rect 203156 161415 203208 161424
rect 203156 161381 203165 161415
rect 203165 161381 203199 161415
rect 203199 161381 203208 161415
rect 203156 161372 203208 161381
rect 217232 161372 217284 161424
rect 345664 161415 345716 161424
rect 345664 161381 345673 161415
rect 345673 161381 345707 161415
rect 345707 161381 345716 161415
rect 345664 161372 345716 161381
rect 182180 161347 182232 161356
rect 182180 161313 182189 161347
rect 182189 161313 182223 161347
rect 182223 161313 182232 161347
rect 182180 161304 182232 161313
rect 236276 160080 236328 160132
rect 225420 160012 225472 160064
rect 225604 160012 225656 160064
rect 361212 160055 361264 160064
rect 361212 160021 361221 160055
rect 361221 160021 361255 160055
rect 361255 160021 361264 160055
rect 361212 160012 361264 160021
rect 177120 158763 177172 158772
rect 177120 158729 177129 158763
rect 177129 158729 177163 158763
rect 177163 158729 177172 158763
rect 177120 158720 177172 158729
rect 178040 158652 178092 158704
rect 178132 158652 178184 158704
rect 225604 158695 225656 158704
rect 225604 158661 225613 158695
rect 225613 158661 225647 158695
rect 225647 158661 225656 158695
rect 225604 158652 225656 158661
rect 228364 158652 228416 158704
rect 228548 158652 228600 158704
rect 343272 158695 343324 158704
rect 343272 158661 343281 158695
rect 343281 158661 343315 158695
rect 343315 158661 343324 158695
rect 343272 158652 343324 158661
rect 272984 157972 273036 158024
rect 273260 157972 273312 158024
rect 328184 157360 328236 157412
rect 329472 157360 329524 157412
rect 228548 157292 228600 157344
rect 258264 157335 258316 157344
rect 258264 157301 258273 157335
rect 258273 157301 258307 157335
rect 258307 157301 258316 157335
rect 258264 157292 258316 157301
rect 291936 157292 291988 157344
rect 317144 157335 317196 157344
rect 317144 157301 317153 157335
rect 317153 157301 317187 157335
rect 317187 157301 317196 157335
rect 317144 157292 317196 157301
rect 318432 157335 318484 157344
rect 318432 157301 318441 157335
rect 318441 157301 318475 157335
rect 318475 157301 318484 157335
rect 318432 157292 318484 157301
rect 232136 157224 232188 157276
rect 328276 157224 328328 157276
rect 354312 157335 354364 157344
rect 354312 157301 354321 157335
rect 354321 157301 354355 157335
rect 354355 157301 354364 157335
rect 354312 157292 354364 157301
rect 329564 157224 329616 157276
rect 291936 157156 291988 157208
rect 232044 157088 232096 157140
rect 192208 156791 192260 156800
rect 192208 156757 192217 156791
rect 192217 156757 192251 156791
rect 192251 156757 192260 156791
rect 192208 156748 192260 156757
rect 182180 156723 182232 156732
rect 182180 156689 182189 156723
rect 182189 156689 182223 156723
rect 182223 156689 182232 156723
rect 182180 156680 182232 156689
rect 362408 156655 362460 156664
rect 362408 156621 362417 156655
rect 362417 156621 362451 156655
rect 362451 156621 362460 156655
rect 362408 156612 362460 156621
rect 273168 154640 273220 154692
rect 211896 154615 211948 154624
rect 211896 154581 211905 154615
rect 211905 154581 211939 154615
rect 211939 154581 211948 154615
rect 211896 154572 211948 154581
rect 212448 154615 212500 154624
rect 212448 154581 212457 154615
rect 212457 154581 212491 154615
rect 212491 154581 212500 154615
rect 212448 154572 212500 154581
rect 234988 154504 235040 154556
rect 235172 154504 235224 154556
rect 273168 154504 273220 154556
rect 291936 154547 291988 154556
rect 291936 154513 291945 154547
rect 291945 154513 291979 154547
rect 291979 154513 291988 154547
rect 291936 154504 291988 154513
rect 315764 153280 315816 153332
rect 315856 153280 315908 153332
rect 192116 153212 192168 153264
rect 229284 153255 229336 153264
rect 229284 153221 229293 153255
rect 229293 153221 229327 153255
rect 229327 153221 229336 153255
rect 229284 153212 229336 153221
rect 261116 153255 261168 153264
rect 261116 153221 261125 153255
rect 261125 153221 261159 153255
rect 261159 153221 261168 153255
rect 261116 153212 261168 153221
rect 283840 153212 283892 153264
rect 283932 153212 283984 153264
rect 286692 153255 286744 153264
rect 286692 153221 286701 153255
rect 286701 153221 286735 153255
rect 286735 153221 286744 153255
rect 286692 153212 286744 153221
rect 341984 153255 342036 153264
rect 341984 153221 341993 153255
rect 341993 153221 342027 153255
rect 342027 153221 342036 153255
rect 341984 153212 342036 153221
rect 355508 153255 355560 153264
rect 355508 153221 355517 153255
rect 355517 153221 355551 153255
rect 355551 153221 355560 153255
rect 355508 153212 355560 153221
rect 191104 153144 191156 153196
rect 191196 153144 191248 153196
rect 230940 153187 230992 153196
rect 230940 153153 230949 153187
rect 230949 153153 230983 153187
rect 230983 153153 230992 153187
rect 230940 153144 230992 153153
rect 231768 153144 231820 153196
rect 232044 153144 232096 153196
rect 277032 153144 277084 153196
rect 277124 153144 277176 153196
rect 270132 152464 270184 152516
rect 270316 152464 270368 152516
rect 230572 152056 230624 152108
rect 230756 152056 230808 152108
rect 179880 151784 179932 151836
rect 179972 151784 180024 151836
rect 181076 151827 181128 151836
rect 181076 151793 181085 151827
rect 181085 151793 181119 151827
rect 181119 151793 181128 151827
rect 181076 151784 181128 151793
rect 217140 151827 217192 151836
rect 217140 151793 217149 151827
rect 217149 151793 217183 151827
rect 217183 151793 217192 151827
rect 217140 151784 217192 151793
rect 344468 151784 344520 151836
rect 344560 151784 344612 151836
rect 345664 151827 345716 151836
rect 345664 151793 345673 151827
rect 345673 151793 345707 151827
rect 345707 151793 345716 151827
rect 345664 151784 345716 151793
rect 3332 151716 3384 151768
rect 21364 151716 21416 151768
rect 361304 150424 361356 150476
rect 225604 150331 225656 150340
rect 225604 150297 225613 150331
rect 225613 150297 225647 150331
rect 225647 150297 225656 150331
rect 225604 150288 225656 150297
rect 177120 149039 177172 149048
rect 177120 149005 177129 149039
rect 177129 149005 177163 149039
rect 177163 149005 177172 149039
rect 177120 148996 177172 149005
rect 178132 149039 178184 149048
rect 178132 149005 178141 149039
rect 178141 149005 178175 149039
rect 178175 149005 178184 149039
rect 178132 148996 178184 149005
rect 299204 147815 299256 147824
rect 299204 147781 299213 147815
rect 299213 147781 299247 147815
rect 299247 147781 299256 147815
rect 299204 147772 299256 147781
rect 300492 147815 300544 147824
rect 300492 147781 300501 147815
rect 300501 147781 300535 147815
rect 300535 147781 300544 147815
rect 300492 147772 300544 147781
rect 354404 147772 354456 147824
rect 184020 147704 184072 147756
rect 189356 147704 189408 147756
rect 200396 147704 200448 147756
rect 201868 147704 201920 147756
rect 273076 147704 273128 147756
rect 273260 147704 273312 147756
rect 315764 147704 315816 147756
rect 211896 147636 211948 147688
rect 217140 147636 217192 147688
rect 258172 147636 258224 147688
rect 258356 147636 258408 147688
rect 184020 147568 184072 147620
rect 189356 147568 189408 147620
rect 200396 147568 200448 147620
rect 201868 147568 201920 147620
rect 211988 147568 212040 147620
rect 317236 147679 317288 147688
rect 317236 147645 317245 147679
rect 317245 147645 317279 147679
rect 317279 147645 317288 147679
rect 317236 147636 317288 147645
rect 328276 147679 328328 147688
rect 328276 147645 328285 147679
rect 328285 147645 328319 147679
rect 328319 147645 328328 147679
rect 328276 147636 328328 147645
rect 354404 147636 354456 147688
rect 217232 147568 217284 147620
rect 315764 147568 315816 147620
rect 291936 145027 291988 145036
rect 291936 144993 291945 145027
rect 291945 144993 291979 145027
rect 291979 144993 291988 145027
rect 291936 144984 291988 144993
rect 224040 144916 224092 144968
rect 224132 144916 224184 144968
rect 299204 144959 299256 144968
rect 299204 144925 299213 144959
rect 299213 144925 299247 144959
rect 299247 144925 299256 144959
rect 299204 144916 299256 144925
rect 300492 144959 300544 144968
rect 300492 144925 300501 144959
rect 300501 144925 300535 144959
rect 300535 144925 300544 144959
rect 300492 144916 300544 144925
rect 328276 144959 328328 144968
rect 328276 144925 328285 144959
rect 328285 144925 328319 144959
rect 328319 144925 328328 144959
rect 328276 144916 328328 144925
rect 171416 144848 171468 144900
rect 171600 144848 171652 144900
rect 173072 144848 173124 144900
rect 173256 144848 173308 144900
rect 203156 144891 203208 144900
rect 203156 144857 203165 144891
rect 203165 144857 203199 144891
rect 203199 144857 203208 144891
rect 203156 144848 203208 144857
rect 211988 144848 212040 144900
rect 230940 144891 230992 144900
rect 230940 144857 230949 144891
rect 230949 144857 230983 144891
rect 230983 144857 230992 144891
rect 230940 144848 230992 144857
rect 258264 144891 258316 144900
rect 258264 144857 258273 144891
rect 258273 144857 258307 144891
rect 258307 144857 258316 144891
rect 258264 144848 258316 144857
rect 329564 144891 329616 144900
rect 329564 144857 329573 144891
rect 329573 144857 329607 144891
rect 329607 144857 329616 144891
rect 329564 144848 329616 144857
rect 362408 144891 362460 144900
rect 362408 144857 362417 144891
rect 362417 144857 362451 144891
rect 362451 144857 362460 144891
rect 362408 144848 362460 144857
rect 317236 143599 317288 143608
rect 317236 143565 317245 143599
rect 317245 143565 317279 143599
rect 317279 143565 317288 143599
rect 317236 143556 317288 143565
rect 261116 143531 261168 143540
rect 261116 143497 261125 143531
rect 261125 143497 261159 143531
rect 261159 143497 261168 143531
rect 261116 143488 261168 143497
rect 275928 143488 275980 143540
rect 285312 143531 285364 143540
rect 285312 143497 285321 143531
rect 285321 143497 285355 143531
rect 285355 143497 285364 143531
rect 285312 143488 285364 143497
rect 286600 143531 286652 143540
rect 286600 143497 286609 143531
rect 286609 143497 286643 143531
rect 286643 143497 286652 143531
rect 286600 143488 286652 143497
rect 289360 143531 289412 143540
rect 289360 143497 289369 143531
rect 289369 143497 289403 143531
rect 289403 143497 289412 143531
rect 289360 143488 289412 143497
rect 291844 143488 291896 143540
rect 291936 143488 291988 143540
rect 318524 143488 318576 143540
rect 230572 142808 230624 142860
rect 230756 142808 230808 142860
rect 234988 142808 235040 142860
rect 235264 142808 235316 142860
rect 270132 142808 270184 142860
rect 270316 142808 270368 142860
rect 236184 142196 236236 142248
rect 236276 142196 236328 142248
rect 341984 142171 342036 142180
rect 341984 142137 341993 142171
rect 341993 142137 342027 142171
rect 342027 142137 342036 142171
rect 341984 142128 342036 142137
rect 181076 142103 181128 142112
rect 181076 142069 181085 142103
rect 181085 142069 181119 142103
rect 181119 142069 181128 142103
rect 181076 142060 181128 142069
rect 182180 142103 182232 142112
rect 182180 142069 182189 142103
rect 182189 142069 182223 142103
rect 182223 142069 182232 142103
rect 182180 142060 182232 142069
rect 229284 142060 229336 142112
rect 229376 142060 229428 142112
rect 235080 142060 235132 142112
rect 236184 142060 236236 142112
rect 315856 142103 315908 142112
rect 315856 142069 315865 142103
rect 315865 142069 315899 142103
rect 315899 142069 315908 142103
rect 315856 142060 315908 142069
rect 361396 142103 361448 142112
rect 361396 142069 361405 142103
rect 361405 142069 361439 142103
rect 361439 142069 361448 142103
rect 361396 142060 361448 142069
rect 235172 141992 235224 142044
rect 225236 140768 225288 140820
rect 225604 140768 225656 140820
rect 341984 140811 342036 140820
rect 341984 140777 341993 140811
rect 341993 140777 342027 140811
rect 342027 140777 342036 140811
rect 341984 140768 342036 140777
rect 343364 140768 343416 140820
rect 344284 140768 344336 140820
rect 344376 140768 344428 140820
rect 179972 140743 180024 140752
rect 179972 140709 179981 140743
rect 179981 140709 180015 140743
rect 180015 140709 180024 140743
rect 179972 140700 180024 140709
rect 194968 140700 195020 140752
rect 212356 140700 212408 140752
rect 177120 139519 177172 139528
rect 177120 139485 177129 139519
rect 177129 139485 177163 139519
rect 177163 139485 177172 139519
rect 177120 139476 177172 139485
rect 178132 139519 178184 139528
rect 178132 139485 178141 139519
rect 178141 139485 178175 139519
rect 178175 139485 178184 139519
rect 178132 139476 178184 139485
rect 228180 139451 228232 139460
rect 228180 139417 228189 139451
rect 228189 139417 228223 139451
rect 228223 139417 228232 139451
rect 228180 139408 228232 139417
rect 177120 139383 177172 139392
rect 177120 139349 177129 139383
rect 177129 139349 177163 139383
rect 177163 139349 177172 139383
rect 177120 139340 177172 139349
rect 178132 139383 178184 139392
rect 178132 139349 178141 139383
rect 178141 139349 178175 139383
rect 178175 139349 178184 139383
rect 178132 139340 178184 139349
rect 341984 139340 342036 139392
rect 232044 139204 232096 139256
rect 232320 139204 232372 139256
rect 345572 138048 345624 138100
rect 345848 138048 345900 138100
rect 258264 137955 258316 137964
rect 258264 137921 258273 137955
rect 258273 137921 258307 137955
rect 258307 137921 258316 137955
rect 258264 137912 258316 137921
rect 285312 137955 285364 137964
rect 285312 137921 285321 137955
rect 285321 137921 285355 137955
rect 285355 137921 285364 137955
rect 285312 137912 285364 137921
rect 286600 137955 286652 137964
rect 286600 137921 286609 137955
rect 286609 137921 286643 137955
rect 286643 137921 286652 137955
rect 286600 137912 286652 137921
rect 289360 137955 289412 137964
rect 289360 137921 289369 137955
rect 289369 137921 289403 137955
rect 289403 137921 289412 137955
rect 289360 137912 289412 137921
rect 2780 136484 2832 136536
rect 5080 136484 5132 136536
rect 211896 135303 211948 135312
rect 211896 135269 211905 135303
rect 211905 135269 211939 135303
rect 211939 135269 211948 135303
rect 211896 135260 211948 135269
rect 329564 135303 329616 135312
rect 329564 135269 329573 135303
rect 329573 135269 329607 135303
rect 329607 135269 329616 135303
rect 329564 135260 329616 135269
rect 183928 135192 183980 135244
rect 184020 135192 184072 135244
rect 231032 135192 231084 135244
rect 231216 135192 231268 135244
rect 272984 135192 273036 135244
rect 273076 135192 273128 135244
rect 317144 135192 317196 135244
rect 317236 135192 317288 135244
rect 203248 133968 203300 134020
rect 318432 134011 318484 134020
rect 318432 133977 318441 134011
rect 318441 133977 318475 134011
rect 318475 133977 318484 134011
rect 318432 133968 318484 133977
rect 217140 133900 217192 133952
rect 217232 133900 217284 133952
rect 261116 133943 261168 133952
rect 261116 133909 261125 133943
rect 261125 133909 261159 133943
rect 261159 133909 261168 133943
rect 261116 133900 261168 133909
rect 275836 133943 275888 133952
rect 275836 133909 275845 133943
rect 275845 133909 275879 133943
rect 275879 133909 275888 133943
rect 275836 133900 275888 133909
rect 201868 133832 201920 133884
rect 277216 133875 277268 133884
rect 277216 133841 277225 133875
rect 277225 133841 277259 133875
rect 277259 133841 277268 133875
rect 277216 133832 277268 133841
rect 284024 133832 284076 133884
rect 284300 133832 284352 133884
rect 291752 133832 291804 133884
rect 291936 133832 291988 133884
rect 318432 133875 318484 133884
rect 318432 133841 318441 133875
rect 318441 133841 318475 133875
rect 318475 133841 318484 133875
rect 318432 133832 318484 133841
rect 225328 133764 225380 133816
rect 225512 133764 225564 133816
rect 228272 133764 228324 133816
rect 228456 133764 228508 133816
rect 181168 132540 181220 132592
rect 203064 132515 203116 132524
rect 203064 132481 203073 132515
rect 203073 132481 203107 132515
rect 203107 132481 203116 132515
rect 203064 132472 203116 132481
rect 315856 132515 315908 132524
rect 315856 132481 315865 132515
rect 315865 132481 315899 132515
rect 315899 132481 315908 132515
rect 315856 132472 315908 132481
rect 343272 132472 343324 132524
rect 343364 132472 343416 132524
rect 361396 132515 361448 132524
rect 361396 132481 361405 132515
rect 361405 132481 361439 132515
rect 361439 132481 361448 132515
rect 361396 132472 361448 132481
rect 181168 132404 181220 132456
rect 345572 132447 345624 132456
rect 345572 132413 345581 132447
rect 345581 132413 345615 132447
rect 345615 132413 345624 132447
rect 345572 132404 345624 132413
rect 344284 132336 344336 132388
rect 344560 132336 344612 132388
rect 270132 131928 270184 131980
rect 270316 131928 270368 131980
rect 180156 131112 180208 131164
rect 194876 131155 194928 131164
rect 194876 131121 194885 131155
rect 194885 131121 194919 131155
rect 194919 131121 194928 131155
rect 194876 131112 194928 131121
rect 212356 131112 212408 131164
rect 343272 131087 343324 131096
rect 343272 131053 343281 131087
rect 343281 131053 343315 131087
rect 343315 131053 343324 131087
rect 343272 131044 343324 131053
rect 177120 129795 177172 129804
rect 177120 129761 177129 129795
rect 177129 129761 177163 129795
rect 177163 129761 177172 129795
rect 177120 129752 177172 129761
rect 178408 129752 178460 129804
rect 341708 129795 341760 129804
rect 341708 129761 341717 129795
rect 341717 129761 341751 129795
rect 341751 129761 341760 129795
rect 341708 129752 341760 129761
rect 299204 128503 299256 128512
rect 299204 128469 299213 128503
rect 299213 128469 299247 128503
rect 299247 128469 299256 128503
rect 299204 128460 299256 128469
rect 300492 128503 300544 128512
rect 300492 128469 300501 128503
rect 300501 128469 300535 128503
rect 300535 128469 300544 128503
rect 300492 128460 300544 128469
rect 189356 128324 189408 128376
rect 191104 128392 191156 128444
rect 211896 128324 211948 128376
rect 258172 128324 258224 128376
rect 258356 128324 258408 128376
rect 328276 128367 328328 128376
rect 328276 128333 328285 128367
rect 328285 128333 328319 128367
rect 328319 128333 328328 128367
rect 328276 128324 328328 128333
rect 354404 128367 354456 128376
rect 354404 128333 354413 128367
rect 354413 128333 354447 128367
rect 354447 128333 354456 128367
rect 354404 128324 354456 128333
rect 355692 128367 355744 128376
rect 355692 128333 355701 128367
rect 355701 128333 355735 128367
rect 355735 128333 355744 128367
rect 355692 128324 355744 128333
rect 189448 128256 189500 128308
rect 191012 128256 191064 128308
rect 211988 128256 212040 128308
rect 179972 127644 180024 127696
rect 180156 127644 180208 127696
rect 362316 127644 362368 127696
rect 362592 127644 362644 127696
rect 285312 125604 285364 125656
rect 285404 125604 285456 125656
rect 286600 125604 286652 125656
rect 286692 125604 286744 125656
rect 289360 125604 289412 125656
rect 289452 125604 289504 125656
rect 171416 125579 171468 125588
rect 171416 125545 171425 125579
rect 171425 125545 171459 125579
rect 171459 125545 171468 125579
rect 171416 125536 171468 125545
rect 173072 125579 173124 125588
rect 173072 125545 173081 125579
rect 173081 125545 173115 125579
rect 173115 125545 173124 125579
rect 173072 125536 173124 125545
rect 183928 125536 183980 125588
rect 184112 125536 184164 125588
rect 191012 125536 191064 125588
rect 191196 125536 191248 125588
rect 211988 125536 212040 125588
rect 235080 125536 235132 125588
rect 258264 125579 258316 125588
rect 258264 125545 258273 125579
rect 258273 125545 258307 125579
rect 258307 125545 258316 125579
rect 258264 125536 258316 125545
rect 318432 125579 318484 125588
rect 318432 125545 318441 125579
rect 318441 125545 318475 125579
rect 318475 125545 318484 125579
rect 318432 125536 318484 125545
rect 329564 125579 329616 125588
rect 329564 125545 329573 125579
rect 329573 125545 329607 125579
rect 329607 125545 329616 125579
rect 329564 125536 329616 125545
rect 355784 125536 355836 125588
rect 235172 125468 235224 125520
rect 355784 125400 355836 125452
rect 182180 124219 182232 124228
rect 182180 124185 182189 124219
rect 182189 124185 182223 124219
rect 182223 124185 182232 124219
rect 182180 124176 182232 124185
rect 194876 124176 194928 124228
rect 194968 124176 195020 124228
rect 201776 124219 201828 124228
rect 201776 124185 201785 124219
rect 201785 124185 201819 124219
rect 201819 124185 201828 124219
rect 201776 124176 201828 124185
rect 232228 124176 232280 124228
rect 232320 124176 232372 124228
rect 277216 124219 277268 124228
rect 277216 124185 277225 124219
rect 277225 124185 277259 124219
rect 277259 124185 277268 124219
rect 277216 124176 277268 124185
rect 299204 124219 299256 124228
rect 299204 124185 299213 124219
rect 299213 124185 299247 124219
rect 299247 124185 299256 124219
rect 299204 124176 299256 124185
rect 300492 124219 300544 124228
rect 300492 124185 300501 124219
rect 300501 124185 300535 124219
rect 300535 124185 300544 124219
rect 300492 124176 300544 124185
rect 328276 124219 328328 124228
rect 328276 124185 328285 124219
rect 328285 124185 328319 124219
rect 328319 124185 328328 124219
rect 328276 124176 328328 124185
rect 354404 124219 354456 124228
rect 354404 124185 354413 124219
rect 354413 124185 354447 124219
rect 354447 124185 354456 124219
rect 354404 124176 354456 124185
rect 355692 124219 355744 124228
rect 355692 124185 355701 124219
rect 355701 124185 355735 124219
rect 355735 124185 355744 124219
rect 355692 124176 355744 124185
rect 361304 124176 361356 124228
rect 361396 124176 361448 124228
rect 192208 124108 192260 124160
rect 192300 124108 192352 124160
rect 200304 124151 200356 124160
rect 200304 124117 200313 124151
rect 200313 124117 200347 124151
rect 200347 124117 200356 124151
rect 200304 124108 200356 124117
rect 203064 124151 203116 124160
rect 203064 124117 203073 124151
rect 203073 124117 203107 124151
rect 203107 124117 203116 124151
rect 203064 124108 203116 124117
rect 231124 124108 231176 124160
rect 261116 124151 261168 124160
rect 261116 124117 261125 124151
rect 261125 124117 261159 124151
rect 261159 124117 261168 124151
rect 261116 124108 261168 124117
rect 275928 124108 275980 124160
rect 276020 124108 276072 124160
rect 291936 124151 291988 124160
rect 291936 124117 291945 124151
rect 291945 124117 291979 124151
rect 291979 124117 291988 124151
rect 291936 124108 291988 124117
rect 318524 124151 318576 124160
rect 318524 124117 318533 124151
rect 318533 124117 318567 124151
rect 318567 124117 318576 124151
rect 318524 124108 318576 124117
rect 270132 123496 270184 123548
rect 270316 123496 270368 123548
rect 181076 122859 181128 122868
rect 181076 122825 181085 122859
rect 181085 122825 181119 122859
rect 181119 122825 181128 122859
rect 181076 122816 181128 122825
rect 345572 122859 345624 122868
rect 345572 122825 345581 122859
rect 345581 122825 345615 122859
rect 345615 122825 345624 122859
rect 345572 122816 345624 122825
rect 182180 122791 182232 122800
rect 182180 122757 182189 122791
rect 182189 122757 182223 122791
rect 182223 122757 182232 122791
rect 182180 122748 182232 122757
rect 192300 122791 192352 122800
rect 192300 122757 192309 122791
rect 192309 122757 192343 122791
rect 192343 122757 192352 122791
rect 192300 122748 192352 122757
rect 225236 122748 225288 122800
rect 225328 122748 225380 122800
rect 229284 122748 229336 122800
rect 232320 122748 232372 122800
rect 344468 122748 344520 122800
rect 344560 122748 344612 122800
rect 181076 122680 181128 122732
rect 2780 122272 2832 122324
rect 4988 122272 5040 122324
rect 343272 121499 343324 121508
rect 343272 121465 343281 121499
rect 343281 121465 343315 121499
rect 343315 121465 343324 121499
rect 343272 121456 343324 121465
rect 212356 121388 212408 121440
rect 362316 121431 362368 121440
rect 362316 121397 362325 121431
rect 362325 121397 362359 121431
rect 362359 121397 362368 121431
rect 362316 121388 362368 121397
rect 236276 120683 236328 120692
rect 236276 120649 236285 120683
rect 236285 120649 236319 120683
rect 236319 120649 236328 120683
rect 236276 120640 236328 120649
rect 178316 120071 178368 120080
rect 178316 120037 178325 120071
rect 178325 120037 178359 120071
rect 178359 120037 178368 120071
rect 178316 120028 178368 120037
rect 277216 118779 277268 118788
rect 277216 118745 277225 118779
rect 277225 118745 277259 118779
rect 277259 118745 277268 118779
rect 277216 118736 277268 118745
rect 315856 118779 315908 118788
rect 315856 118745 315865 118779
rect 315865 118745 315899 118779
rect 315899 118745 315908 118779
rect 315856 118736 315908 118745
rect 235264 118711 235316 118720
rect 235264 118677 235273 118711
rect 235273 118677 235307 118711
rect 235307 118677 235316 118711
rect 235264 118668 235316 118677
rect 258264 118643 258316 118652
rect 258264 118609 258273 118643
rect 258273 118609 258307 118643
rect 258307 118609 258316 118643
rect 258264 118600 258316 118609
rect 182180 118031 182232 118040
rect 182180 117997 182189 118031
rect 182189 117997 182223 118031
rect 182223 117997 182232 118031
rect 182180 117988 182232 117997
rect 229284 117988 229336 118040
rect 171416 115991 171468 116000
rect 171416 115957 171425 115991
rect 171425 115957 171459 115991
rect 171459 115957 171468 115991
rect 171416 115948 171468 115957
rect 173072 115991 173124 116000
rect 173072 115957 173081 115991
rect 173081 115957 173115 115991
rect 173115 115957 173124 115991
rect 173072 115948 173124 115957
rect 194968 115948 195020 116000
rect 201776 115948 201828 116000
rect 201868 115948 201920 116000
rect 211896 115991 211948 116000
rect 211896 115957 211905 115991
rect 211905 115957 211939 115991
rect 211939 115957 211948 115991
rect 211896 115948 211948 115957
rect 235264 115991 235316 116000
rect 235264 115957 235273 115991
rect 235273 115957 235307 115991
rect 235307 115957 235316 115991
rect 235264 115948 235316 115957
rect 282828 115948 282880 116000
rect 329564 115991 329616 116000
rect 329564 115957 329573 115991
rect 329573 115957 329607 115991
rect 329607 115957 329616 115991
rect 329564 115948 329616 115957
rect 361212 115948 361264 116000
rect 361304 115948 361356 116000
rect 184020 115923 184072 115932
rect 184020 115889 184029 115923
rect 184029 115889 184063 115923
rect 184063 115889 184072 115923
rect 184020 115880 184072 115889
rect 189356 115880 189408 115932
rect 189448 115880 189500 115932
rect 194876 115880 194928 115932
rect 273076 115923 273128 115932
rect 273076 115889 273085 115923
rect 273085 115889 273119 115923
rect 273119 115889 273128 115923
rect 273076 115880 273128 115889
rect 286416 115880 286468 115932
rect 286692 115880 286744 115932
rect 289176 115880 289228 115932
rect 289452 115880 289504 115932
rect 362316 115923 362368 115932
rect 362316 115889 362325 115923
rect 362325 115889 362359 115923
rect 362359 115889 362368 115923
rect 362316 115880 362368 115889
rect 200580 115812 200632 115864
rect 354404 114588 354456 114640
rect 203248 114520 203300 114572
rect 231032 114563 231084 114572
rect 231032 114529 231041 114563
rect 231041 114529 231075 114563
rect 231075 114529 231084 114563
rect 231032 114520 231084 114529
rect 261116 114563 261168 114572
rect 261116 114529 261125 114563
rect 261125 114529 261159 114563
rect 261159 114529 261168 114563
rect 261116 114520 261168 114529
rect 282736 114563 282788 114572
rect 194876 114495 194928 114504
rect 194876 114461 194885 114495
rect 194885 114461 194919 114495
rect 194919 114461 194928 114495
rect 194876 114452 194928 114461
rect 201868 114495 201920 114504
rect 201868 114461 201877 114495
rect 201877 114461 201911 114495
rect 201911 114461 201920 114495
rect 201868 114452 201920 114461
rect 282736 114529 282745 114563
rect 282745 114529 282779 114563
rect 282779 114529 282788 114563
rect 282736 114520 282788 114529
rect 291936 114563 291988 114572
rect 291936 114529 291945 114563
rect 291945 114529 291979 114563
rect 291979 114529 291988 114563
rect 291936 114520 291988 114529
rect 315856 114563 315908 114572
rect 315856 114529 315865 114563
rect 315865 114529 315899 114563
rect 315899 114529 315908 114563
rect 315856 114520 315908 114529
rect 318524 114563 318576 114572
rect 318524 114529 318533 114563
rect 318533 114529 318567 114563
rect 318567 114529 318576 114563
rect 318524 114520 318576 114529
rect 328184 114520 328236 114572
rect 328276 114520 328328 114572
rect 230756 113840 230808 113892
rect 230940 113840 230992 113892
rect 270132 113840 270184 113892
rect 270316 113840 270368 113892
rect 232228 113203 232280 113212
rect 232228 113169 232237 113203
rect 232237 113169 232271 113203
rect 232271 113169 232280 113203
rect 232228 113160 232280 113169
rect 341800 113160 341852 113212
rect 341892 113160 341944 113212
rect 354220 113203 354272 113212
rect 354220 113169 354229 113203
rect 354229 113169 354263 113203
rect 354263 113169 354272 113203
rect 354220 113160 354272 113169
rect 212356 113092 212408 113144
rect 219900 113092 219952 113144
rect 355600 113135 355652 113144
rect 355600 113101 355609 113135
rect 355609 113101 355643 113135
rect 355643 113101 355652 113135
rect 355600 113092 355652 113101
rect 341892 113067 341944 113076
rect 341892 113033 341901 113067
rect 341901 113033 341935 113067
rect 341935 113033 341944 113067
rect 341892 113024 341944 113033
rect 181076 111868 181128 111920
rect 217048 111800 217100 111852
rect 217232 111800 217284 111852
rect 181076 111775 181128 111784
rect 181076 111741 181085 111775
rect 181085 111741 181119 111775
rect 181119 111741 181128 111775
rect 181076 111732 181128 111741
rect 217048 111707 217100 111716
rect 217048 111673 217057 111707
rect 217057 111673 217091 111707
rect 217091 111673 217100 111707
rect 217048 111664 217100 111673
rect 230756 111052 230808 111104
rect 231032 111052 231084 111104
rect 176936 110440 176988 110492
rect 177120 110440 177172 110492
rect 178500 110440 178552 110492
rect 192392 110372 192444 110424
rect 317236 109735 317288 109744
rect 317236 109701 317245 109735
rect 317245 109701 317279 109735
rect 317279 109701 317288 109735
rect 317236 109692 317288 109701
rect 354220 109692 354272 109744
rect 318524 109352 318576 109404
rect 300492 109191 300544 109200
rect 300492 109157 300501 109191
rect 300501 109157 300535 109191
rect 300535 109157 300544 109191
rect 300492 109148 300544 109157
rect 182180 109012 182232 109064
rect 211896 109012 211948 109064
rect 3332 108944 3384 108996
rect 28264 108944 28316 108996
rect 236368 109080 236420 109132
rect 258172 109012 258224 109064
rect 258356 109012 258408 109064
rect 285404 109080 285456 109132
rect 315856 109123 315908 109132
rect 315856 109089 315865 109123
rect 315865 109089 315899 109123
rect 315899 109089 315908 109123
rect 315856 109080 315908 109089
rect 328276 109012 328328 109064
rect 211988 108944 212040 108996
rect 236276 108944 236328 108996
rect 285312 108944 285364 108996
rect 182180 108876 182232 108928
rect 328276 108876 328328 108928
rect 184112 108808 184164 108860
rect 178132 106904 178184 106956
rect 178500 106904 178552 106956
rect 273076 106335 273128 106344
rect 273076 106301 273085 106335
rect 273085 106301 273119 106335
rect 273119 106301 273128 106335
rect 273076 106292 273128 106301
rect 171416 106267 171468 106276
rect 171416 106233 171425 106267
rect 171425 106233 171459 106267
rect 171459 106233 171468 106267
rect 171416 106224 171468 106233
rect 173072 106267 173124 106276
rect 173072 106233 173081 106267
rect 173081 106233 173115 106267
rect 173115 106233 173124 106267
rect 173072 106224 173124 106233
rect 211988 106224 212040 106276
rect 235080 106224 235132 106276
rect 236276 106267 236328 106276
rect 236276 106233 236285 106267
rect 236285 106233 236319 106267
rect 236319 106233 236328 106267
rect 236276 106224 236328 106233
rect 258264 106267 258316 106276
rect 258264 106233 258273 106267
rect 258273 106233 258307 106267
rect 258307 106233 258316 106267
rect 258264 106224 258316 106233
rect 329564 106267 329616 106276
rect 329564 106233 329573 106267
rect 329573 106233 329607 106267
rect 329607 106233 329616 106267
rect 329564 106224 329616 106233
rect 235172 106156 235224 106208
rect 270132 105408 270184 105460
rect 270316 105408 270368 105460
rect 277216 104975 277268 104984
rect 277216 104941 277225 104975
rect 277225 104941 277259 104975
rect 277259 104941 277268 104975
rect 277216 104932 277268 104941
rect 176936 104864 176988 104916
rect 177028 104864 177080 104916
rect 194968 104864 195020 104916
rect 202052 104864 202104 104916
rect 315856 104907 315908 104916
rect 315856 104873 315865 104907
rect 315865 104873 315899 104907
rect 315899 104873 315908 104907
rect 315856 104864 315908 104873
rect 318340 104907 318392 104916
rect 318340 104873 318349 104907
rect 318349 104873 318383 104907
rect 318383 104873 318392 104907
rect 318340 104864 318392 104873
rect 261116 104839 261168 104848
rect 261116 104805 261125 104839
rect 261125 104805 261159 104839
rect 261159 104805 261168 104839
rect 261116 104796 261168 104805
rect 275928 104796 275980 104848
rect 277216 104796 277268 104848
rect 282736 104839 282788 104848
rect 282736 104805 282745 104839
rect 282745 104805 282779 104839
rect 282779 104805 282788 104839
rect 282736 104796 282788 104805
rect 284024 104796 284076 104848
rect 182180 104771 182232 104780
rect 182180 104737 182189 104771
rect 182189 104737 182223 104771
rect 182223 104737 182232 104771
rect 182180 104728 182232 104737
rect 230756 104184 230808 104236
rect 230940 104184 230992 104236
rect 219808 103615 219860 103624
rect 219808 103581 219817 103615
rect 219817 103581 219851 103615
rect 219851 103581 219860 103615
rect 219808 103572 219860 103581
rect 299204 103547 299256 103556
rect 299204 103513 299213 103547
rect 299213 103513 299247 103547
rect 299247 103513 299256 103547
rect 299204 103504 299256 103513
rect 300492 103547 300544 103556
rect 300492 103513 300501 103547
rect 300501 103513 300535 103547
rect 300535 103513 300544 103547
rect 300492 103504 300544 103513
rect 341984 103504 342036 103556
rect 355692 103504 355744 103556
rect 219808 103436 219860 103488
rect 344560 103436 344612 103488
rect 181076 102255 181128 102264
rect 181076 102221 181085 102255
rect 181085 102221 181119 102255
rect 181119 102221 181128 102255
rect 181076 102212 181128 102221
rect 299204 102255 299256 102264
rect 299204 102221 299213 102255
rect 299213 102221 299247 102255
rect 299247 102221 299256 102255
rect 299204 102212 299256 102221
rect 217232 102144 217284 102196
rect 177028 102119 177080 102128
rect 177028 102085 177037 102119
rect 177037 102085 177071 102119
rect 177071 102085 177080 102119
rect 177028 102076 177080 102085
rect 179972 102119 180024 102128
rect 179972 102085 179981 102119
rect 179981 102085 180015 102119
rect 180015 102085 180024 102119
rect 179972 102076 180024 102085
rect 181076 102076 181128 102128
rect 181444 102076 181496 102128
rect 298928 102076 298980 102128
rect 299204 102076 299256 102128
rect 177948 102008 178000 102060
rect 178132 102008 178184 102060
rect 211988 100036 212040 100088
rect 225328 99671 225380 99680
rect 225328 99637 225337 99671
rect 225337 99637 225371 99671
rect 225371 99637 225380 99671
rect 225328 99628 225380 99637
rect 224040 99535 224092 99544
rect 224040 99501 224049 99535
rect 224049 99501 224083 99535
rect 224083 99501 224092 99535
rect 224040 99492 224092 99501
rect 235264 99399 235316 99408
rect 235264 99365 235273 99399
rect 235273 99365 235307 99399
rect 235307 99365 235316 99399
rect 235264 99356 235316 99365
rect 182272 99288 182324 99340
rect 258264 99331 258316 99340
rect 258264 99297 258273 99331
rect 258273 99297 258307 99331
rect 258307 99297 258316 99331
rect 258264 99288 258316 99297
rect 315764 96951 315816 96960
rect 315764 96917 315773 96951
rect 315773 96917 315807 96951
rect 315807 96917 315816 96951
rect 315764 96908 315816 96917
rect 171416 96679 171468 96688
rect 171416 96645 171425 96679
rect 171425 96645 171459 96679
rect 171459 96645 171468 96679
rect 171416 96636 171468 96645
rect 173072 96679 173124 96688
rect 173072 96645 173081 96679
rect 173081 96645 173115 96679
rect 173115 96645 173124 96679
rect 173072 96636 173124 96645
rect 235264 96679 235316 96688
rect 235264 96645 235273 96679
rect 235273 96645 235307 96679
rect 235307 96645 235316 96679
rect 235264 96636 235316 96645
rect 236368 96636 236420 96688
rect 291936 96636 291988 96688
rect 292028 96636 292080 96688
rect 317236 96679 317288 96688
rect 317236 96645 317245 96679
rect 317245 96645 317279 96679
rect 317279 96645 317288 96679
rect 317236 96636 317288 96645
rect 329564 96679 329616 96688
rect 329564 96645 329573 96679
rect 329573 96645 329607 96679
rect 329607 96645 329616 96679
rect 329564 96636 329616 96645
rect 354404 96679 354456 96688
rect 354404 96645 354413 96679
rect 354413 96645 354447 96679
rect 354447 96645 354456 96679
rect 354404 96636 354456 96645
rect 232044 96568 232096 96620
rect 232228 96568 232280 96620
rect 235172 96568 235224 96620
rect 235356 96568 235408 96620
rect 217232 95387 217284 95396
rect 217232 95353 217241 95387
rect 217241 95353 217275 95387
rect 217275 95353 217284 95387
rect 217232 95344 217284 95353
rect 191012 95208 191064 95260
rect 191196 95208 191248 95260
rect 192392 95208 192444 95260
rect 224132 95208 224184 95260
rect 225328 95251 225380 95260
rect 225328 95217 225337 95251
rect 225337 95217 225371 95251
rect 225371 95217 225380 95251
rect 225328 95208 225380 95217
rect 261116 95251 261168 95260
rect 261116 95217 261125 95251
rect 261125 95217 261159 95251
rect 261159 95217 261168 95251
rect 261116 95208 261168 95217
rect 275836 95251 275888 95260
rect 275836 95217 275845 95251
rect 275845 95217 275879 95251
rect 275879 95217 275888 95251
rect 275836 95208 275888 95217
rect 277124 95251 277176 95260
rect 277124 95217 277133 95251
rect 277133 95217 277167 95251
rect 277167 95217 277176 95251
rect 277124 95208 277176 95217
rect 282736 95251 282788 95260
rect 282736 95217 282745 95251
rect 282745 95217 282779 95251
rect 282779 95217 282788 95251
rect 282736 95208 282788 95217
rect 283932 95251 283984 95260
rect 283932 95217 283941 95251
rect 283941 95217 283975 95251
rect 283975 95217 283984 95251
rect 283932 95208 283984 95217
rect 194968 95140 195020 95192
rect 178040 95115 178092 95124
rect 178040 95081 178049 95115
rect 178049 95081 178083 95115
rect 178083 95081 178092 95115
rect 178040 95072 178092 95081
rect 192392 95072 192444 95124
rect 230756 94528 230808 94580
rect 230940 94528 230992 94580
rect 270132 94528 270184 94580
rect 270316 94528 270368 94580
rect 219716 93891 219768 93900
rect 219716 93857 219725 93891
rect 219725 93857 219759 93891
rect 219759 93857 219768 93891
rect 219716 93848 219768 93857
rect 343088 93848 343140 93900
rect 343180 93848 343232 93900
rect 344468 93891 344520 93900
rect 344468 93857 344477 93891
rect 344477 93857 344511 93891
rect 344511 93857 344520 93891
rect 344468 93848 344520 93857
rect 182272 93780 182324 93832
rect 355692 93823 355744 93832
rect 355692 93789 355701 93823
rect 355701 93789 355735 93823
rect 355735 93789 355744 93823
rect 355692 93780 355744 93789
rect 361212 93823 361264 93832
rect 361212 93789 361221 93823
rect 361221 93789 361255 93823
rect 361255 93789 361264 93823
rect 361212 93780 361264 93789
rect 177120 92488 177172 92540
rect 179972 92531 180024 92540
rect 179972 92497 179981 92531
rect 179981 92497 180015 92531
rect 180015 92497 180024 92531
rect 179972 92488 180024 92497
rect 178132 91060 178184 91112
rect 192116 90380 192168 90432
rect 192392 90380 192444 90432
rect 236368 89768 236420 89820
rect 258172 89700 258224 89752
rect 258356 89700 258408 89752
rect 236368 89632 236420 89684
rect 191196 86980 191248 87032
rect 315764 87023 315816 87032
rect 315764 86989 315773 87023
rect 315773 86989 315807 87023
rect 315807 86989 315816 87023
rect 315764 86980 315816 86989
rect 171416 86955 171468 86964
rect 171416 86921 171425 86955
rect 171425 86921 171459 86955
rect 171459 86921 171468 86955
rect 171416 86912 171468 86921
rect 173072 86955 173124 86964
rect 173072 86921 173081 86955
rect 173081 86921 173115 86955
rect 173115 86921 173124 86955
rect 173072 86912 173124 86921
rect 191104 86912 191156 86964
rect 201868 86955 201920 86964
rect 201868 86921 201877 86955
rect 201877 86921 201911 86955
rect 201911 86921 201920 86955
rect 201868 86912 201920 86921
rect 211896 86912 211948 86964
rect 211988 86912 212040 86964
rect 225236 86912 225288 86964
rect 225328 86912 225380 86964
rect 228180 86912 228232 86964
rect 228272 86912 228324 86964
rect 229284 86912 229336 86964
rect 235080 86912 235132 86964
rect 236276 86955 236328 86964
rect 236276 86921 236285 86955
rect 236285 86921 236319 86955
rect 236319 86921 236328 86955
rect 236276 86912 236328 86921
rect 258264 86955 258316 86964
rect 258264 86921 258273 86955
rect 258273 86921 258307 86955
rect 258307 86921 258316 86955
rect 258264 86912 258316 86921
rect 262404 86912 262456 86964
rect 229376 86844 229428 86896
rect 235172 86844 235224 86896
rect 270132 86096 270184 86148
rect 270316 86096 270368 86148
rect 200396 85620 200448 85672
rect 177028 85552 177080 85604
rect 177120 85552 177172 85604
rect 194876 85595 194928 85604
rect 194876 85561 194885 85595
rect 194885 85561 194919 85595
rect 194919 85561 194928 85595
rect 194876 85552 194928 85561
rect 200304 85552 200356 85604
rect 224040 85552 224092 85604
rect 224132 85552 224184 85604
rect 362316 85552 362368 85604
rect 362500 85552 362552 85604
rect 212264 85484 212316 85536
rect 212448 85484 212500 85536
rect 228180 85484 228232 85536
rect 228272 85484 228324 85536
rect 261116 85484 261168 85536
rect 283932 85527 283984 85536
rect 283932 85493 283941 85527
rect 283941 85493 283975 85527
rect 283975 85493 283984 85527
rect 283932 85484 283984 85493
rect 289360 85484 289412 85536
rect 361212 85527 361264 85536
rect 361212 85493 361221 85527
rect 361221 85493 361255 85527
rect 361255 85493 361264 85527
rect 361212 85484 361264 85493
rect 230756 84872 230808 84924
rect 230940 84872 230992 84924
rect 341984 84328 342036 84380
rect 182180 84235 182232 84244
rect 182180 84201 182189 84235
rect 182189 84201 182223 84235
rect 182223 84201 182232 84235
rect 182180 84192 182232 84201
rect 217232 84235 217284 84244
rect 217232 84201 217241 84235
rect 217241 84201 217275 84235
rect 217275 84201 217284 84235
rect 217232 84192 217284 84201
rect 219532 84192 219584 84244
rect 219808 84192 219860 84244
rect 341984 84192 342036 84244
rect 355692 84235 355744 84244
rect 355692 84201 355701 84235
rect 355701 84201 355735 84235
rect 355735 84201 355744 84235
rect 355692 84192 355744 84201
rect 191104 84167 191156 84176
rect 191104 84133 191113 84167
rect 191113 84133 191147 84167
rect 191147 84133 191156 84167
rect 191104 84124 191156 84133
rect 192208 84124 192260 84176
rect 275744 84124 275796 84176
rect 275928 84124 275980 84176
rect 343272 84167 343324 84176
rect 343272 84133 343281 84167
rect 343281 84133 343315 84167
rect 343315 84133 343324 84167
rect 343272 84124 343324 84133
rect 345572 84167 345624 84176
rect 345572 84133 345581 84167
rect 345581 84133 345615 84167
rect 345615 84133 345624 84167
rect 345572 84124 345624 84133
rect 361304 84167 361356 84176
rect 361304 84133 361313 84167
rect 361313 84133 361347 84167
rect 361347 84133 361356 84167
rect 361304 84124 361356 84133
rect 362500 84124 362552 84176
rect 179972 82807 180024 82816
rect 179972 82773 179981 82807
rect 179981 82773 180015 82807
rect 180015 82773 180024 82807
rect 179972 82764 180024 82773
rect 178132 81379 178184 81388
rect 178132 81345 178141 81379
rect 178141 81345 178175 81379
rect 178175 81345 178184 81379
rect 178132 81336 178184 81345
rect 203064 80699 203116 80708
rect 203064 80665 203073 80699
rect 203073 80665 203107 80699
rect 203107 80665 203116 80699
rect 203064 80656 203116 80665
rect 235264 80087 235316 80096
rect 235264 80053 235273 80087
rect 235273 80053 235307 80087
rect 235307 80053 235316 80087
rect 235264 80044 235316 80053
rect 291936 80044 291988 80096
rect 291844 79976 291896 80028
rect 344560 79339 344612 79348
rect 344560 79305 344569 79339
rect 344569 79305 344603 79339
rect 344603 79305 344612 79339
rect 344560 79296 344612 79305
rect 361396 79296 361448 79348
rect 318524 77528 318576 77580
rect 229376 77460 229428 77512
rect 171416 77299 171468 77308
rect 171416 77265 171425 77299
rect 171425 77265 171459 77299
rect 171459 77265 171468 77299
rect 171416 77256 171468 77265
rect 173072 77299 173124 77308
rect 173072 77265 173081 77299
rect 173081 77265 173115 77299
rect 173115 77265 173124 77299
rect 173072 77256 173124 77265
rect 200304 77256 200356 77308
rect 200396 77256 200448 77308
rect 201868 77299 201920 77308
rect 201868 77265 201877 77299
rect 201877 77265 201911 77299
rect 201911 77265 201920 77299
rect 201868 77256 201920 77265
rect 224040 77324 224092 77376
rect 229376 77324 229428 77376
rect 282828 77324 282880 77376
rect 232228 77299 232280 77308
rect 232228 77265 232237 77299
rect 232237 77265 232271 77299
rect 232271 77265 232280 77299
rect 232228 77256 232280 77265
rect 235264 77299 235316 77308
rect 235264 77265 235273 77299
rect 235273 77265 235307 77299
rect 235307 77265 235316 77299
rect 235264 77256 235316 77265
rect 258356 77256 258408 77308
rect 262312 77299 262364 77308
rect 262312 77265 262321 77299
rect 262321 77265 262355 77299
rect 262355 77265 262364 77299
rect 262312 77256 262364 77265
rect 182364 77188 182416 77240
rect 194876 77231 194928 77240
rect 194876 77197 194885 77231
rect 194885 77197 194919 77231
rect 194919 77197 194928 77231
rect 194876 77188 194928 77197
rect 223948 77188 224000 77240
rect 182364 77052 182416 77104
rect 189356 75896 189408 75948
rect 189448 75896 189500 75948
rect 217140 75896 217192 75948
rect 217324 75896 217376 75948
rect 232228 75939 232280 75948
rect 232228 75905 232237 75939
rect 232237 75905 232271 75939
rect 232271 75905 232280 75939
rect 232228 75896 232280 75905
rect 236460 75896 236512 75948
rect 260932 75939 260984 75948
rect 260932 75905 260941 75939
rect 260941 75905 260975 75939
rect 260975 75905 260984 75939
rect 260932 75896 260984 75905
rect 282736 75939 282788 75948
rect 282736 75905 282745 75939
rect 282745 75905 282779 75939
rect 282779 75905 282788 75939
rect 282736 75896 282788 75905
rect 284024 75896 284076 75948
rect 289268 75939 289320 75948
rect 289268 75905 289277 75939
rect 289277 75905 289311 75939
rect 289311 75905 289320 75939
rect 289268 75896 289320 75905
rect 318248 75939 318300 75948
rect 318248 75905 318257 75939
rect 318257 75905 318291 75939
rect 318291 75905 318300 75939
rect 318248 75896 318300 75905
rect 184020 75871 184072 75880
rect 184020 75837 184029 75871
rect 184029 75837 184063 75871
rect 184063 75837 184072 75871
rect 184020 75828 184072 75837
rect 355968 75871 356020 75880
rect 355968 75837 355977 75871
rect 355977 75837 356011 75871
rect 356011 75837 356020 75871
rect 355968 75828 356020 75837
rect 217140 75803 217192 75812
rect 217140 75769 217149 75803
rect 217149 75769 217183 75803
rect 217183 75769 217192 75803
rect 217140 75760 217192 75769
rect 355876 75760 355928 75812
rect 355784 75692 355836 75744
rect 355876 75624 355928 75676
rect 355784 75556 355836 75608
rect 230756 75216 230808 75268
rect 230940 75216 230992 75268
rect 270132 75216 270184 75268
rect 270316 75216 270368 75268
rect 277124 74604 277176 74656
rect 277216 74604 277268 74656
rect 341984 74647 342036 74656
rect 341984 74613 341993 74647
rect 341993 74613 342027 74647
rect 342027 74613 342036 74647
rect 341984 74604 342036 74613
rect 191288 74536 191340 74588
rect 343364 74536 343416 74588
rect 345664 74536 345716 74588
rect 181260 74511 181312 74520
rect 181260 74477 181269 74511
rect 181269 74477 181303 74511
rect 181303 74477 181312 74511
rect 181260 74468 181312 74477
rect 341984 73287 342036 73296
rect 341984 73253 341993 73287
rect 341993 73253 342027 73287
rect 342027 73253 342036 73287
rect 341984 73244 342036 73253
rect 179972 73219 180024 73228
rect 179972 73185 179981 73219
rect 179981 73185 180015 73219
rect 180015 73185 180024 73219
rect 179972 73176 180024 73185
rect 203064 71111 203116 71120
rect 203064 71077 203073 71111
rect 203073 71077 203107 71111
rect 203107 71077 203116 71111
rect 203064 71068 203116 71077
rect 211896 70456 211948 70508
rect 219808 70456 219860 70508
rect 258172 70388 258224 70440
rect 211896 70320 211948 70372
rect 258264 70320 258316 70372
rect 329564 67736 329616 67788
rect 235172 67668 235224 67720
rect 225236 67600 225288 67652
rect 225328 67600 225380 67652
rect 232044 67600 232096 67652
rect 232228 67600 232280 67652
rect 235080 67600 235132 67652
rect 236276 67600 236328 67652
rect 236460 67600 236512 67652
rect 282736 67600 282788 67652
rect 282828 67600 282880 67652
rect 285220 67600 285272 67652
rect 285312 67600 285364 67652
rect 286508 67600 286560 67652
rect 286600 67600 286652 67652
rect 289268 67600 289320 67652
rect 289360 67600 289412 67652
rect 317052 67600 317104 67652
rect 317236 67600 317288 67652
rect 329564 67600 329616 67652
rect 344560 67643 344612 67652
rect 344560 67609 344569 67643
rect 344569 67609 344603 67643
rect 344603 67609 344612 67643
rect 344560 67600 344612 67609
rect 362316 67643 362368 67652
rect 362316 67609 362325 67643
rect 362325 67609 362359 67643
rect 362359 67609 362368 67643
rect 362316 67600 362368 67609
rect 171416 67575 171468 67584
rect 171416 67541 171425 67575
rect 171425 67541 171459 67575
rect 171459 67541 171468 67575
rect 171416 67532 171468 67541
rect 173072 67575 173124 67584
rect 173072 67541 173081 67575
rect 173081 67541 173115 67575
rect 173115 67541 173124 67575
rect 173072 67532 173124 67541
rect 223948 67532 224000 67584
rect 229284 67532 229336 67584
rect 224040 67464 224092 67516
rect 229376 67464 229428 67516
rect 362224 67464 362276 67516
rect 362316 67464 362368 67516
rect 355968 67371 356020 67380
rect 355968 67337 355977 67371
rect 355977 67337 356011 67371
rect 356011 67337 356020 67371
rect 355968 67328 356020 67337
rect 184112 66240 184164 66292
rect 192208 66240 192260 66292
rect 194968 66240 195020 66292
rect 217232 66240 217284 66292
rect 219716 66283 219768 66292
rect 219716 66249 219725 66283
rect 219725 66249 219759 66283
rect 219759 66249 219768 66283
rect 219716 66240 219768 66249
rect 203064 66172 203116 66224
rect 203340 66172 203392 66224
rect 212264 66172 212316 66224
rect 212356 66172 212408 66224
rect 235080 66172 235132 66224
rect 275836 66172 275888 66224
rect 284024 66172 284076 66224
rect 285312 66215 285364 66224
rect 285312 66181 285321 66215
rect 285321 66181 285355 66215
rect 285355 66181 285364 66215
rect 285312 66172 285364 66181
rect 286600 66215 286652 66224
rect 286600 66181 286609 66215
rect 286609 66181 286643 66215
rect 286643 66181 286652 66215
rect 286600 66172 286652 66181
rect 289360 66215 289412 66224
rect 289360 66181 289369 66215
rect 289369 66181 289403 66215
rect 289403 66181 289412 66215
rect 289360 66172 289412 66181
rect 291936 66172 291988 66224
rect 329564 66215 329616 66224
rect 235172 66104 235224 66156
rect 329564 66181 329573 66215
rect 329573 66181 329607 66215
rect 329607 66181 329616 66215
rect 329564 66172 329616 66181
rect 276020 66104 276072 66156
rect 292028 66104 292080 66156
rect 230756 65943 230808 65952
rect 230756 65909 230765 65943
rect 230765 65909 230799 65943
rect 230799 65909 230808 65943
rect 230756 65900 230808 65909
rect 234988 65492 235040 65544
rect 235264 65492 235316 65544
rect 270132 65492 270184 65544
rect 270316 65492 270368 65544
rect 181076 64880 181128 64932
rect 341892 64880 341944 64932
rect 203340 64812 203392 64864
rect 344560 64812 344612 64864
rect 355692 64812 355744 64864
rect 341984 64744 342036 64796
rect 178316 63520 178368 63572
rect 177028 63495 177080 63504
rect 177028 63461 177037 63495
rect 177037 63461 177071 63495
rect 177071 63461 177080 63495
rect 177028 63452 177080 63461
rect 179972 63495 180024 63504
rect 179972 63461 179981 63495
rect 179981 63461 180015 63495
rect 180015 63461 180024 63495
rect 179972 63452 180024 63461
rect 275928 63452 275980 63504
rect 277216 63452 277268 63504
rect 341984 63452 342036 63504
rect 343180 63452 343232 63504
rect 343364 63452 343416 63504
rect 341892 63384 341944 63436
rect 200396 61455 200448 61464
rect 200396 61421 200405 61455
rect 200405 61421 200439 61455
rect 200439 61421 200448 61455
rect 200396 61412 200448 61421
rect 201868 61455 201920 61464
rect 201868 61421 201877 61455
rect 201877 61421 201911 61455
rect 201911 61421 201920 61455
rect 201868 61412 201920 61421
rect 262404 60664 262456 60716
rect 262588 60664 262640 60716
rect 234988 60596 235040 60648
rect 235264 60596 235316 60648
rect 345572 59984 345624 60036
rect 181076 58667 181128 58676
rect 181076 58633 181085 58667
rect 181085 58633 181119 58667
rect 181119 58633 181128 58667
rect 181076 58624 181128 58633
rect 354404 58148 354456 58200
rect 354404 58012 354456 58064
rect 171416 57987 171468 57996
rect 171416 57953 171425 57987
rect 171425 57953 171459 57987
rect 171459 57953 171468 57987
rect 171416 57944 171468 57953
rect 173072 57987 173124 57996
rect 173072 57953 173081 57987
rect 173081 57953 173115 57987
rect 173115 57953 173124 57987
rect 173072 57944 173124 57953
rect 315764 57944 315816 57996
rect 315856 57944 315908 57996
rect 328184 57944 328236 57996
rect 328276 57944 328328 57996
rect 177120 57876 177172 57928
rect 183928 57876 183980 57928
rect 184112 57876 184164 57928
rect 261024 57876 261076 57928
rect 261116 57876 261168 57928
rect 262588 57876 262640 57928
rect 318340 57876 318392 57928
rect 318524 57876 318576 57928
rect 354404 57876 354456 57928
rect 362316 57919 362368 57928
rect 362316 57885 362325 57919
rect 362325 57885 362359 57919
rect 362359 57885 362368 57919
rect 362316 57876 362368 57885
rect 283932 56695 283984 56704
rect 283932 56661 283941 56695
rect 283941 56661 283975 56695
rect 283975 56661 283984 56695
rect 283932 56652 283984 56661
rect 219716 56584 219768 56636
rect 219808 56584 219860 56636
rect 231032 56584 231084 56636
rect 285404 56584 285456 56636
rect 286692 56584 286744 56636
rect 289452 56584 289504 56636
rect 329564 56627 329616 56636
rect 329564 56593 329573 56627
rect 329573 56593 329607 56627
rect 329607 56593 329616 56627
rect 329564 56584 329616 56593
rect 225236 56516 225288 56568
rect 225512 56516 225564 56568
rect 261024 56516 261076 56568
rect 283932 56559 283984 56568
rect 283932 56525 283941 56559
rect 283941 56525 283975 56559
rect 283975 56525 283984 56559
rect 283932 56516 283984 56525
rect 318340 56559 318392 56568
rect 318340 56525 318349 56559
rect 318349 56525 318383 56559
rect 318383 56525 318392 56559
rect 318340 56516 318392 56525
rect 231032 56448 231084 56500
rect 231400 56448 231452 56500
rect 261208 56448 261260 56500
rect 203064 55267 203116 55276
rect 203064 55233 203073 55267
rect 203073 55233 203107 55267
rect 203107 55233 203116 55267
rect 203064 55224 203116 55233
rect 344468 55267 344520 55276
rect 344468 55233 344477 55267
rect 344477 55233 344511 55267
rect 344511 55233 344520 55267
rect 344468 55224 344520 55233
rect 183928 55199 183980 55208
rect 183928 55165 183937 55199
rect 183937 55165 183971 55199
rect 183971 55165 183980 55199
rect 183928 55156 183980 55165
rect 228180 55199 228232 55208
rect 228180 55165 228189 55199
rect 228189 55165 228223 55199
rect 228223 55165 228232 55199
rect 228180 55156 228232 55165
rect 270132 54612 270184 54664
rect 270316 54612 270368 54664
rect 202052 53932 202104 53984
rect 178040 53796 178092 53848
rect 178132 53796 178184 53848
rect 179972 53839 180024 53848
rect 179972 53805 179981 53839
rect 179981 53805 180015 53839
rect 180015 53805 180024 53839
rect 179972 53796 180024 53805
rect 181168 53796 181220 53848
rect 275744 53839 275796 53848
rect 275744 53805 275753 53839
rect 275753 53805 275787 53839
rect 275787 53805 275796 53839
rect 275744 53796 275796 53805
rect 275744 53116 275796 53168
rect 275928 53116 275980 53168
rect 327908 53116 327960 53168
rect 328276 53116 328328 53168
rect 344468 51756 344520 51808
rect 192208 51076 192260 51128
rect 224040 51076 224092 51128
rect 229376 51076 229428 51128
rect 192116 51008 192168 51060
rect 232136 51076 232188 51128
rect 235264 51076 235316 51128
rect 232044 51008 232096 51060
rect 273076 51076 273128 51128
rect 235356 51008 235408 51060
rect 272984 51008 273036 51060
rect 291844 51008 291896 51060
rect 292028 51008 292080 51060
rect 224040 50940 224092 50992
rect 229376 50940 229428 50992
rect 2780 50124 2832 50176
rect 4896 50124 4948 50176
rect 235172 48356 235224 48408
rect 354312 48399 354364 48408
rect 354312 48365 354321 48399
rect 354321 48365 354355 48399
rect 354355 48365 354364 48399
rect 354312 48356 354364 48365
rect 200488 48288 200540 48340
rect 235080 48288 235132 48340
rect 258264 48288 258316 48340
rect 258356 48288 258408 48340
rect 262496 48331 262548 48340
rect 262496 48297 262505 48331
rect 262505 48297 262539 48331
rect 262539 48297 262548 48331
rect 262496 48288 262548 48297
rect 277216 48288 277268 48340
rect 285312 48288 285364 48340
rect 285404 48288 285456 48340
rect 286600 48288 286652 48340
rect 286692 48288 286744 48340
rect 289360 48288 289412 48340
rect 289452 48288 289504 48340
rect 355600 48331 355652 48340
rect 355600 48297 355609 48331
rect 355609 48297 355643 48331
rect 355643 48297 355652 48331
rect 355600 48288 355652 48297
rect 362500 48288 362552 48340
rect 171416 48263 171468 48272
rect 171416 48229 171425 48263
rect 171425 48229 171459 48263
rect 171459 48229 171468 48263
rect 171416 48220 171468 48229
rect 189448 48220 189500 48272
rect 189540 48220 189592 48272
rect 211896 48220 211948 48272
rect 211988 48220 212040 48272
rect 212448 48263 212500 48272
rect 212448 48229 212457 48263
rect 212457 48229 212491 48263
rect 212491 48229 212500 48263
rect 212448 48220 212500 48229
rect 275836 48220 275888 48272
rect 275928 48220 275980 48272
rect 282736 48220 282788 48272
rect 282828 48220 282880 48272
rect 354312 48263 354364 48272
rect 354312 48229 354321 48263
rect 354321 48229 354355 48263
rect 354355 48229 354364 48263
rect 354312 48220 354364 48229
rect 291752 48152 291804 48204
rect 291844 48152 291896 48204
rect 270132 47404 270184 47456
rect 270316 47404 270368 47456
rect 284024 46928 284076 46980
rect 318432 46928 318484 46980
rect 345664 46971 345716 46980
rect 345664 46937 345673 46971
rect 345673 46937 345707 46971
rect 345707 46937 345716 46971
rect 345664 46928 345716 46937
rect 194968 46860 195020 46912
rect 195152 46860 195204 46912
rect 228272 46860 228324 46912
rect 232044 46903 232096 46912
rect 232044 46869 232053 46903
rect 232053 46869 232087 46903
rect 232087 46869 232096 46903
rect 232044 46860 232096 46869
rect 261208 46860 261260 46912
rect 261300 46860 261352 46912
rect 317144 46903 317196 46912
rect 317144 46869 317153 46903
rect 317153 46869 317187 46903
rect 317187 46869 317196 46903
rect 317144 46860 317196 46869
rect 179972 45636 180024 45688
rect 181168 45636 181220 45688
rect 181076 45568 181128 45620
rect 183928 45611 183980 45620
rect 183928 45577 183937 45611
rect 183937 45577 183971 45611
rect 183971 45577 183980 45611
rect 183928 45568 183980 45577
rect 341892 45568 341944 45620
rect 201960 45500 202012 45552
rect 228180 45500 228232 45552
rect 228272 45500 228324 45552
rect 231216 45500 231268 45552
rect 231308 45500 231360 45552
rect 272984 45500 273036 45552
rect 341892 45432 341944 45484
rect 190920 44140 190972 44192
rect 191104 44140 191156 44192
rect 181352 44072 181404 44124
rect 219808 42483 219860 42492
rect 219808 42449 219817 42483
rect 219817 42449 219851 42483
rect 219851 42449 219860 42483
rect 219808 42440 219860 42449
rect 329472 42100 329524 42152
rect 182180 41463 182232 41472
rect 182180 41429 182189 41463
rect 182189 41429 182223 41463
rect 182223 41429 182232 41463
rect 182180 41420 182232 41429
rect 234804 41420 234856 41472
rect 235080 41420 235132 41472
rect 236276 41420 236328 41472
rect 262404 41352 262456 41404
rect 262588 41352 262640 41404
rect 236276 41284 236328 41336
rect 344560 41123 344612 41132
rect 344560 41089 344569 41123
rect 344569 41089 344603 41123
rect 344603 41089 344612 41123
rect 344560 41080 344612 41089
rect 354312 41123 354364 41132
rect 354312 41089 354321 41123
rect 354321 41089 354355 41123
rect 354355 41089 354364 41123
rect 354312 41080 354364 41089
rect 189540 40715 189592 40724
rect 189540 40681 189549 40715
rect 189549 40681 189583 40715
rect 189583 40681 189592 40715
rect 189540 40672 189592 40681
rect 367100 40264 367152 40316
rect 369952 40264 370004 40316
rect 270500 40196 270552 40248
rect 275744 40196 275796 40248
rect 398748 40196 398800 40248
rect 405648 40196 405700 40248
rect 212448 40060 212500 40112
rect 220728 40060 220780 40112
rect 201500 39924 201552 39976
rect 201868 39924 201920 39976
rect 284116 38700 284168 38752
rect 284208 38700 284260 38752
rect 171416 38675 171468 38684
rect 171416 38641 171425 38675
rect 171425 38641 171459 38675
rect 171459 38641 171468 38675
rect 171416 38632 171468 38641
rect 191196 38632 191248 38684
rect 230756 38632 230808 38684
rect 230940 38632 230992 38684
rect 191104 38564 191156 38616
rect 211896 38564 211948 38616
rect 211988 38564 212040 38616
rect 229284 38564 229336 38616
rect 229376 38564 229428 38616
rect 235080 38564 235132 38616
rect 235264 38564 235316 38616
rect 258356 38564 258408 38616
rect 275836 38607 275888 38616
rect 275836 38573 275845 38607
rect 275845 38573 275879 38607
rect 275879 38573 275888 38607
rect 275836 38564 275888 38573
rect 284116 38564 284168 38616
rect 284208 38564 284260 38616
rect 344652 38607 344704 38616
rect 344652 38573 344661 38607
rect 344661 38573 344695 38607
rect 344695 38573 344704 38607
rect 344652 38564 344704 38573
rect 283932 38496 283984 38548
rect 284300 38496 284352 38548
rect 328276 37408 328328 37460
rect 200396 37272 200448 37324
rect 200488 37272 200540 37324
rect 212356 37272 212408 37324
rect 217140 37272 217192 37324
rect 217232 37272 217284 37324
rect 225236 37272 225288 37324
rect 225512 37272 225564 37324
rect 232044 37315 232096 37324
rect 232044 37281 232053 37315
rect 232053 37281 232087 37315
rect 232087 37281 232096 37315
rect 232044 37272 232096 37281
rect 282736 37272 282788 37324
rect 282828 37272 282880 37324
rect 317236 37272 317288 37324
rect 328276 37272 328328 37324
rect 329380 37315 329432 37324
rect 329380 37281 329389 37315
rect 329389 37281 329423 37315
rect 329423 37281 329432 37315
rect 329380 37272 329432 37281
rect 343364 37315 343416 37324
rect 343364 37281 343373 37315
rect 343373 37281 343407 37315
rect 343407 37281 343416 37315
rect 343364 37272 343416 37281
rect 272984 37136 273036 37188
rect 178132 35912 178184 35964
rect 178224 35912 178276 35964
rect 180064 35912 180116 35964
rect 219992 35912 220044 35964
rect 2780 35844 2832 35896
rect 4804 35844 4856 35896
rect 270132 35300 270184 35352
rect 270316 35300 270368 35352
rect 284116 33804 284168 33856
rect 318432 33804 318484 33856
rect 318524 33736 318576 33788
rect 284116 33668 284168 33720
rect 275928 33192 275980 33244
rect 196072 31832 196124 31884
rect 266544 31832 266596 31884
rect 362592 31832 362644 31884
rect 178224 31764 178276 31816
rect 180064 31764 180116 31816
rect 234804 31764 234856 31816
rect 285404 31764 285456 31816
rect 286692 31764 286744 31816
rect 291844 31764 291896 31816
rect 328184 31764 328236 31816
rect 361396 31764 361448 31816
rect 178132 31696 178184 31748
rect 179972 31696 180024 31748
rect 196072 31696 196124 31748
rect 234712 31696 234764 31748
rect 258264 31739 258316 31748
rect 258264 31705 258273 31739
rect 258273 31705 258307 31739
rect 258307 31705 258316 31739
rect 258264 31696 258316 31705
rect 266544 31696 266596 31748
rect 285312 31696 285364 31748
rect 286600 31696 286652 31748
rect 291936 31696 291988 31748
rect 370504 30268 370556 30320
rect 580264 30268 580316 30320
rect 231308 29044 231360 29096
rect 232044 28976 232096 29028
rect 232136 28976 232188 29028
rect 261116 28976 261168 29028
rect 261208 28976 261260 29028
rect 284024 28976 284076 29028
rect 284300 28976 284352 29028
rect 289268 28976 289320 29028
rect 289452 28976 289504 29028
rect 317144 28976 317196 29028
rect 317236 28976 317288 29028
rect 344652 29019 344704 29028
rect 344652 28985 344661 29019
rect 344661 28985 344695 29019
rect 344695 28985 344704 29019
rect 344652 28976 344704 28985
rect 361304 29019 361356 29028
rect 361304 28985 361313 29019
rect 361313 28985 361347 29019
rect 361347 28985 361356 29019
rect 361304 28976 361356 28985
rect 362408 29019 362460 29028
rect 362408 28985 362417 29019
rect 362417 28985 362451 29019
rect 362451 28985 362460 29019
rect 362408 28976 362460 28985
rect 171416 28908 171468 28960
rect 173072 28908 173124 28960
rect 173164 28908 173216 28960
rect 184020 28908 184072 28960
rect 184112 28908 184164 28960
rect 203156 28908 203208 28960
rect 203248 28908 203300 28960
rect 231124 28908 231176 28960
rect 236368 28951 236420 28960
rect 236368 28917 236377 28951
rect 236377 28917 236411 28951
rect 236411 28917 236420 28951
rect 236368 28908 236420 28917
rect 329472 28951 329524 28960
rect 329472 28917 329481 28951
rect 329481 28917 329515 28951
rect 329515 28917 329524 28951
rect 329472 28908 329524 28917
rect 317144 28883 317196 28892
rect 317144 28849 317153 28883
rect 317153 28849 317187 28883
rect 317187 28849 317196 28883
rect 317144 28840 317196 28849
rect 343364 28475 343416 28484
rect 343364 28441 343373 28475
rect 343373 28441 343407 28475
rect 343407 28441 343416 28475
rect 343364 28432 343416 28441
rect 272984 27684 273036 27736
rect 182180 27659 182232 27668
rect 182180 27625 182189 27659
rect 182189 27625 182223 27659
rect 182223 27625 182232 27659
rect 189540 27659 189592 27668
rect 182180 27616 182232 27625
rect 189540 27625 189549 27659
rect 189549 27625 189583 27659
rect 189583 27625 189592 27659
rect 189540 27616 189592 27625
rect 200396 27659 200448 27668
rect 200396 27625 200405 27659
rect 200405 27625 200439 27659
rect 200439 27625 200448 27659
rect 200396 27616 200448 27625
rect 201868 27659 201920 27668
rect 201868 27625 201877 27659
rect 201877 27625 201911 27659
rect 201911 27625 201920 27659
rect 201868 27616 201920 27625
rect 219808 27616 219860 27668
rect 219992 27616 220044 27668
rect 273076 27616 273128 27668
rect 328092 27659 328144 27668
rect 328092 27625 328101 27659
rect 328101 27625 328135 27659
rect 328135 27625 328144 27659
rect 328092 27616 328144 27625
rect 212080 27548 212132 27600
rect 212172 27548 212224 27600
rect 212264 27591 212316 27600
rect 212264 27557 212273 27591
rect 212273 27557 212307 27591
rect 212307 27557 212316 27591
rect 261116 27591 261168 27600
rect 212264 27548 212316 27557
rect 261116 27557 261125 27591
rect 261125 27557 261159 27591
rect 261159 27557 261168 27591
rect 261116 27548 261168 27557
rect 268752 27591 268804 27600
rect 268752 27557 268761 27591
rect 268761 27557 268795 27591
rect 268795 27557 268804 27591
rect 268752 27548 268804 27557
rect 275928 27591 275980 27600
rect 275928 27557 275937 27591
rect 275937 27557 275971 27591
rect 275971 27557 275980 27591
rect 275928 27548 275980 27557
rect 277216 27548 277268 27600
rect 343364 27548 343416 27600
rect 344652 27548 344704 27600
rect 345664 27591 345716 27600
rect 345664 27557 345673 27591
rect 345673 27557 345707 27591
rect 345707 27557 345716 27591
rect 345664 27548 345716 27557
rect 354404 27548 354456 27600
rect 355692 27548 355744 27600
rect 361304 27548 361356 27600
rect 270132 26868 270184 26920
rect 270316 26868 270368 26920
rect 230940 26596 230992 26648
rect 231124 26596 231176 26648
rect 181076 26299 181128 26308
rect 181076 26265 181085 26299
rect 181085 26265 181119 26299
rect 181119 26265 181128 26299
rect 181076 26256 181128 26265
rect 200396 26299 200448 26308
rect 200396 26265 200405 26299
rect 200405 26265 200439 26299
rect 200439 26265 200448 26299
rect 200396 26256 200448 26265
rect 178132 26231 178184 26240
rect 178132 26197 178141 26231
rect 178141 26197 178175 26231
rect 178175 26197 178184 26231
rect 178132 26188 178184 26197
rect 179972 26231 180024 26240
rect 179972 26197 179981 26231
rect 179981 26197 180015 26231
rect 180015 26197 180024 26231
rect 179972 26188 180024 26197
rect 182180 26188 182232 26240
rect 182456 26188 182508 26240
rect 194876 26231 194928 26240
rect 194876 26197 194885 26231
rect 194885 26197 194919 26231
rect 194919 26197 194928 26231
rect 194876 26188 194928 26197
rect 181168 26120 181220 26172
rect 181352 26120 181404 26172
rect 234712 25100 234764 25152
rect 235172 25100 235224 25152
rect 266544 23604 266596 23656
rect 266820 23604 266872 23656
rect 200396 22108 200448 22160
rect 217140 22108 217192 22160
rect 291936 22108 291988 22160
rect 214104 22040 214156 22092
rect 214288 22040 214340 22092
rect 262404 22040 262456 22092
rect 262588 22040 262640 22092
rect 200396 21972 200448 22024
rect 217140 21972 217192 22024
rect 291936 21972 291988 22024
rect 171324 19363 171376 19372
rect 171324 19329 171333 19363
rect 171333 19329 171367 19363
rect 171367 19329 171376 19363
rect 171324 19320 171376 19329
rect 223948 19320 224000 19372
rect 224040 19320 224092 19372
rect 229284 19320 229336 19372
rect 229376 19320 229428 19372
rect 236368 19363 236420 19372
rect 236368 19329 236377 19363
rect 236377 19329 236411 19363
rect 236411 19329 236420 19363
rect 236368 19320 236420 19329
rect 317236 19320 317288 19372
rect 329564 19320 329616 19372
rect 192208 19252 192260 19304
rect 212264 19295 212316 19304
rect 212264 19261 212273 19295
rect 212273 19261 212307 19295
rect 212307 19261 212316 19295
rect 212264 19252 212316 19261
rect 214288 19295 214340 19304
rect 214288 19261 214297 19295
rect 214297 19261 214331 19295
rect 214331 19261 214340 19295
rect 214288 19252 214340 19261
rect 291936 19252 291988 19304
rect 328276 19252 328328 19304
rect 352932 19295 352984 19304
rect 352932 19261 352941 19295
rect 352941 19261 352975 19295
rect 352975 19261 352984 19295
rect 352932 19252 352984 19261
rect 362592 19252 362644 19304
rect 341892 18411 341944 18420
rect 341892 18377 341901 18411
rect 341901 18377 341935 18411
rect 341935 18377 341944 18411
rect 341892 18368 341944 18377
rect 219716 18028 219768 18080
rect 182364 18003 182416 18012
rect 182364 17969 182373 18003
rect 182373 17969 182407 18003
rect 182407 17969 182416 18003
rect 182364 17960 182416 17969
rect 219808 17960 219860 18012
rect 261116 18003 261168 18012
rect 261116 17969 261125 18003
rect 261125 17969 261159 18003
rect 261159 17969 261168 18003
rect 261116 17960 261168 17969
rect 268752 18003 268804 18012
rect 268752 17969 268761 18003
rect 268761 17969 268795 18003
rect 268795 17969 268804 18003
rect 268752 17960 268804 17969
rect 272800 17960 272852 18012
rect 272892 17960 272944 18012
rect 275928 18003 275980 18012
rect 275928 17969 275937 18003
rect 275937 17969 275971 18003
rect 275971 17969 275980 18003
rect 275928 17960 275980 17969
rect 345664 18003 345716 18012
rect 345664 17969 345673 18003
rect 345673 17969 345707 18003
rect 345707 17969 345716 18003
rect 345664 17960 345716 17969
rect 354312 18003 354364 18012
rect 354312 17969 354321 18003
rect 354321 17969 354355 18003
rect 354355 17969 354364 18003
rect 354312 17960 354364 17969
rect 355508 18003 355560 18012
rect 355508 17969 355517 18003
rect 355517 17969 355551 18003
rect 355551 17969 355560 18003
rect 355508 17960 355560 17969
rect 361212 18003 361264 18012
rect 361212 17969 361221 18003
rect 361221 17969 361255 18003
rect 361255 17969 361264 18003
rect 361212 17960 361264 17969
rect 169760 17892 169812 17944
rect 579620 17892 579672 17944
rect 182364 17799 182416 17808
rect 182364 17765 182373 17799
rect 182373 17765 182407 17799
rect 182407 17765 182416 17799
rect 182364 17756 182416 17765
rect 270132 17212 270184 17264
rect 270316 17212 270368 17264
rect 230572 16736 230624 16788
rect 230756 16736 230808 16788
rect 177120 16668 177172 16720
rect 177028 16600 177080 16652
rect 178132 16643 178184 16652
rect 178132 16609 178141 16643
rect 178141 16609 178175 16643
rect 178175 16609 178184 16643
rect 178132 16600 178184 16609
rect 179972 16643 180024 16652
rect 179972 16609 179981 16643
rect 179981 16609 180015 16643
rect 180015 16609 180024 16643
rect 179972 16600 180024 16609
rect 194968 16600 195020 16652
rect 296444 14696 296496 14748
rect 367100 14696 367152 14748
rect 297732 14628 297784 14680
rect 371240 14628 371292 14680
rect 299112 14560 299164 14612
rect 375196 14560 375248 14612
rect 300400 14492 300452 14544
rect 378140 14492 378192 14544
rect 358544 14424 358596 14476
rect 546500 14424 546552 14476
rect 499580 13744 499632 13796
rect 502340 13676 502392 13728
rect 506480 13608 506532 13660
rect 346124 13540 346176 13592
rect 510620 13540 510672 13592
rect 347412 13472 347464 13524
rect 517520 13472 517572 13524
rect 348884 13404 348936 13456
rect 520280 13404 520332 13456
rect 350264 13336 350316 13388
rect 524420 13336 524472 13388
rect 351552 13268 351604 13320
rect 528560 13268 528612 13320
rect 354312 13200 354364 13252
rect 535460 13200 535512 13252
rect 355508 13132 355560 13184
rect 538220 13132 538272 13184
rect 289268 13107 289320 13116
rect 289268 13073 289277 13107
rect 289277 13073 289311 13107
rect 289311 13073 289320 13107
rect 289268 13064 289320 13073
rect 357164 13064 357216 13116
rect 542360 13064 542412 13116
rect 340512 12996 340564 13048
rect 495440 12996 495492 13048
rect 339224 12928 339276 12980
rect 492680 12928 492732 12980
rect 337844 12860 337896 12912
rect 488540 12860 488592 12912
rect 337752 12792 337804 12844
rect 485780 12792 485832 12844
rect 335176 12724 335228 12776
rect 480260 12724 480312 12776
rect 333612 12656 333664 12708
rect 477592 12656 477644 12708
rect 212264 12563 212316 12572
rect 212264 12529 212273 12563
rect 212273 12529 212307 12563
rect 212307 12529 212316 12563
rect 212264 12520 212316 12529
rect 234712 12452 234764 12504
rect 235172 12452 235224 12504
rect 285404 12452 285456 12504
rect 286692 12452 286744 12504
rect 329472 12495 329524 12504
rect 329472 12461 329481 12495
rect 329481 12461 329515 12495
rect 329515 12461 329524 12495
rect 329472 12452 329524 12461
rect 171140 12384 171192 12436
rect 171324 12384 171376 12436
rect 211896 12384 211948 12436
rect 212172 12384 212224 12436
rect 265256 12384 265308 12436
rect 265808 12384 265860 12436
rect 285312 12384 285364 12436
rect 286600 12384 286652 12436
rect 332416 12384 332468 12436
rect 469220 12384 469272 12436
rect 333704 12316 333756 12368
rect 473360 12316 473412 12368
rect 335268 12248 335320 12300
rect 478880 12248 478932 12300
rect 336464 12180 336516 12232
rect 484400 12180 484452 12232
rect 337936 12112 337988 12164
rect 487160 12112 487212 12164
rect 339316 12044 339368 12096
rect 491300 12044 491352 12096
rect 340604 11976 340656 12028
rect 494060 11976 494112 12028
rect 342076 11908 342128 11960
rect 498200 11908 498252 11960
rect 125508 11840 125560 11892
rect 212724 11840 212776 11892
rect 343456 11840 343508 11892
rect 502432 11840 502484 11892
rect 121368 11772 121420 11824
rect 211252 11772 211304 11824
rect 344744 11772 344796 11824
rect 505100 11772 505152 11824
rect 31668 11704 31720 11756
rect 180984 11704 181036 11756
rect 531320 11704 531372 11756
rect 304816 11636 304868 11688
rect 390560 11636 390612 11688
rect 303436 11568 303488 11620
rect 387800 11568 387852 11620
rect 302056 11500 302108 11552
rect 383660 11500 383712 11552
rect 300676 11432 300728 11484
rect 380900 11432 380952 11484
rect 300584 11364 300636 11416
rect 376760 11364 376812 11416
rect 299296 11296 299348 11348
rect 374092 11296 374144 11348
rect 297824 11228 297876 11280
rect 369860 11228 369912 11280
rect 366732 11024 366784 11076
rect 367008 11024 367060 11076
rect 103428 10956 103480 11008
rect 204352 10956 204404 11008
rect 307576 10956 307628 11008
rect 397460 10956 397512 11008
rect 99288 10888 99340 10940
rect 202972 10888 203024 10940
rect 308864 10888 308916 10940
rect 400312 10888 400364 10940
rect 96528 10820 96580 10872
rect 201684 10820 201736 10872
rect 336556 10820 336608 10872
rect 483020 10820 483072 10872
rect 92388 10752 92440 10804
rect 201592 10752 201644 10804
rect 338028 10752 338080 10804
rect 485872 10752 485924 10804
rect 89628 10684 89680 10736
rect 200212 10684 200264 10736
rect 339408 10684 339460 10736
rect 489920 10684 489972 10736
rect 85488 10616 85540 10668
rect 198924 10616 198976 10668
rect 340788 10616 340840 10668
rect 494152 10616 494204 10668
rect 82728 10548 82780 10600
rect 197452 10548 197504 10600
rect 340696 10548 340748 10600
rect 496820 10548 496872 10600
rect 78588 10480 78640 10532
rect 195980 10480 196032 10532
rect 342168 10480 342220 10532
rect 500960 10480 501012 10532
rect 74448 10412 74500 10464
rect 194876 10412 194928 10464
rect 343548 10412 343600 10464
rect 503720 10412 503772 10464
rect 71688 10344 71740 10396
rect 193312 10344 193364 10396
rect 344836 10344 344888 10396
rect 507860 10344 507912 10396
rect 28908 10276 28960 10328
rect 179604 10276 179656 10328
rect 347504 10276 347556 10328
rect 513380 10276 513432 10328
rect 107568 10208 107620 10260
rect 205732 10208 205784 10260
rect 306196 10208 306248 10260
rect 393320 10208 393372 10260
rect 110328 10140 110380 10192
rect 207112 10140 207164 10192
rect 304908 10140 304960 10192
rect 390652 10140 390704 10192
rect 114468 10072 114520 10124
rect 208492 10072 208544 10124
rect 303528 10072 303580 10124
rect 386420 10072 386472 10124
rect 150348 10004 150400 10056
rect 221096 10004 221148 10056
rect 302148 10004 302200 10056
rect 382372 10004 382424 10056
rect 153108 9936 153160 9988
rect 222384 9936 222436 9988
rect 300768 9936 300820 9988
rect 379520 9936 379572 9988
rect 157248 9868 157300 9920
rect 223856 9868 223908 9920
rect 299388 9868 299440 9920
rect 375380 9868 375432 9920
rect 284024 9732 284076 9784
rect 189264 9664 189316 9716
rect 189540 9664 189592 9716
rect 192116 9707 192168 9716
rect 192116 9673 192125 9707
rect 192125 9673 192159 9707
rect 192159 9673 192168 9707
rect 192116 9664 192168 9673
rect 212264 9707 212316 9716
rect 212264 9673 212273 9707
rect 212273 9673 212307 9707
rect 212307 9673 212316 9707
rect 212264 9664 212316 9673
rect 214288 9707 214340 9716
rect 214288 9673 214297 9707
rect 214297 9673 214331 9707
rect 214331 9673 214340 9707
rect 214288 9664 214340 9673
rect 277216 9664 277268 9716
rect 291844 9707 291896 9716
rect 291844 9673 291853 9707
rect 291853 9673 291887 9707
rect 291887 9673 291896 9707
rect 291844 9664 291896 9673
rect 328184 9707 328236 9716
rect 328184 9673 328193 9707
rect 328193 9673 328227 9707
rect 328227 9673 328236 9707
rect 328184 9664 328236 9673
rect 329472 9707 329524 9716
rect 329472 9673 329481 9707
rect 329481 9673 329515 9707
rect 329515 9673 329524 9707
rect 329472 9664 329524 9673
rect 362500 9707 362552 9716
rect 362500 9673 362509 9707
rect 362509 9673 362543 9707
rect 362543 9673 362552 9707
rect 362500 9664 362552 9673
rect 138480 9596 138532 9648
rect 216956 9596 217008 9648
rect 317052 9596 317104 9648
rect 427544 9596 427596 9648
rect 137284 9528 137336 9580
rect 134892 9460 134944 9512
rect 215392 9460 215444 9512
rect 216864 9528 216916 9580
rect 318340 9528 318392 9580
rect 431132 9528 431184 9580
rect 319996 9460 320048 9512
rect 434628 9460 434680 9512
rect 131396 9392 131448 9444
rect 214012 9392 214064 9444
rect 321376 9392 321428 9444
rect 438216 9392 438268 9444
rect 133788 9324 133840 9376
rect 215576 9324 215628 9376
rect 322664 9324 322716 9376
rect 441804 9324 441856 9376
rect 130200 9256 130252 9308
rect 214288 9256 214340 9308
rect 322756 9256 322808 9308
rect 445392 9256 445444 9308
rect 126612 9188 126664 9240
rect 212908 9188 212960 9240
rect 324136 9188 324188 9240
rect 448980 9188 449032 9240
rect 67180 9120 67232 9172
rect 192024 9120 192076 9172
rect 325516 9120 325568 9172
rect 452476 9120 452528 9172
rect 23112 9052 23164 9104
rect 177028 9052 177080 9104
rect 180156 9052 180208 9104
rect 230940 9052 230992 9104
rect 326804 9052 326856 9104
rect 456064 9052 456116 9104
rect 18328 8984 18380 9036
rect 175372 8984 175424 9036
rect 177764 8984 177816 9036
rect 230664 8984 230716 9036
rect 328184 8984 328236 9036
rect 459652 8984 459704 9036
rect 13636 8916 13688 8968
rect 173992 8916 174044 8968
rect 176568 8916 176620 8968
rect 230572 8916 230624 8968
rect 329472 8916 329524 8968
rect 463240 8916 463292 8968
rect 140872 8848 140924 8900
rect 218152 8848 218204 8900
rect 315856 8848 315908 8900
rect 423956 8848 424008 8900
rect 142068 8780 142120 8832
rect 218244 8780 218296 8832
rect 314476 8780 314528 8832
rect 420368 8780 420420 8832
rect 145656 8712 145708 8764
rect 219624 8712 219676 8764
rect 313096 8712 313148 8764
rect 416872 8712 416924 8764
rect 117136 8644 117188 8696
rect 179972 8644 180024 8696
rect 311716 8644 311768 8696
rect 413284 8644 413336 8696
rect 162308 8576 162360 8628
rect 225236 8576 225288 8628
rect 311624 8576 311676 8628
rect 409696 8576 409748 8628
rect 165896 8508 165948 8560
rect 226616 8508 226668 8560
rect 310336 8508 310388 8560
rect 406108 8508 406160 8560
rect 169392 8440 169444 8492
rect 227996 8440 228048 8492
rect 308956 8440 309008 8492
rect 402520 8440 402572 8492
rect 172980 8372 173032 8424
rect 229376 8372 229428 8424
rect 307668 8372 307720 8424
rect 399024 8372 399076 8424
rect 181076 8304 181128 8356
rect 181260 8304 181312 8356
rect 182180 8304 182232 8356
rect 182456 8304 182508 8356
rect 283932 8347 283984 8356
rect 283932 8313 283941 8347
rect 283941 8313 283975 8347
rect 283975 8313 283984 8347
rect 283932 8304 283984 8313
rect 306288 8304 306340 8356
rect 395436 8304 395488 8356
rect 101588 8236 101640 8288
rect 204536 8236 204588 8288
rect 355784 8236 355836 8288
rect 541716 8236 541768 8288
rect 98092 8168 98144 8220
rect 203156 8168 203208 8220
rect 357256 8168 357308 8220
rect 545304 8168 545356 8220
rect 94504 8100 94556 8152
rect 201868 8100 201920 8152
rect 358636 8100 358688 8152
rect 548892 8100 548944 8152
rect 90916 8032 90968 8084
rect 200396 8032 200448 8084
rect 346676 8032 346728 8084
rect 359924 8032 359976 8084
rect 552388 8032 552440 8084
rect 87328 7964 87380 8016
rect 198832 7964 198884 8016
rect 289544 7964 289596 8016
rect 349068 7964 349120 8016
rect 361304 7964 361356 8016
rect 555976 7964 556028 8016
rect 83832 7896 83884 7948
rect 198740 7896 198792 7948
rect 290924 7896 290976 7948
rect 352564 7896 352616 7948
rect 363604 7896 363656 7948
rect 559564 7896 559616 7948
rect 80244 7828 80296 7880
rect 197544 7828 197596 7880
rect 292304 7828 292356 7880
rect 356152 7828 356204 7880
rect 364156 7828 364208 7880
rect 563152 7828 563204 7880
rect 76656 7760 76708 7812
rect 196164 7760 196216 7812
rect 293684 7760 293736 7812
rect 359740 7760 359792 7812
rect 365444 7760 365496 7812
rect 566740 7760 566792 7812
rect 63592 7692 63644 7744
rect 191932 7692 191984 7744
rect 294972 7692 295024 7744
rect 363328 7692 363380 7744
rect 366824 7692 366876 7744
rect 570236 7692 570288 7744
rect 60004 7624 60056 7676
rect 190552 7624 190604 7676
rect 296536 7624 296588 7676
rect 366916 7624 366968 7676
rect 367008 7624 367060 7676
rect 573824 7624 573876 7676
rect 56416 7556 56468 7608
rect 189172 7556 189224 7608
rect 295156 7556 295208 7608
rect 364524 7556 364576 7608
rect 368204 7556 368256 7608
rect 577412 7556 577464 7608
rect 105176 7488 105228 7540
rect 205824 7488 205876 7540
rect 355876 7488 355928 7540
rect 538128 7488 538180 7540
rect 108764 7420 108816 7472
rect 207204 7420 207256 7472
rect 354496 7420 354548 7472
rect 534540 7420 534592 7472
rect 112352 7352 112404 7404
rect 208584 7352 208636 7404
rect 353116 7352 353168 7404
rect 531044 7352 531096 7404
rect 115940 7284 115992 7336
rect 209780 7284 209832 7336
rect 351644 7284 351696 7336
rect 527456 7284 527508 7336
rect 119436 7216 119488 7268
rect 209872 7216 209924 7268
rect 350356 7216 350408 7268
rect 523868 7216 523920 7268
rect 123024 7148 123076 7200
rect 211344 7148 211396 7200
rect 348792 7148 348844 7200
rect 520372 7148 520424 7200
rect 153936 7080 153988 7132
rect 222292 7080 222344 7132
rect 347596 7080 347648 7132
rect 516784 7080 516836 7132
rect 157524 7012 157576 7064
rect 223764 7012 223816 7064
rect 346216 7012 346268 7064
rect 513196 7012 513248 7064
rect 161112 6944 161164 6996
rect 225052 6944 225104 6996
rect 344928 6944 344980 6996
rect 509608 6944 509660 6996
rect 129004 6808 129056 6860
rect 213920 6808 213972 6860
rect 320088 6808 320140 6860
rect 437020 6808 437072 6860
rect 73068 6740 73120 6792
rect 194784 6740 194836 6792
rect 321468 6740 321520 6792
rect 440608 6740 440660 6792
rect 49332 6672 49384 6724
rect 186412 6672 186464 6724
rect 322848 6672 322900 6724
rect 444196 6672 444248 6724
rect 44548 6604 44600 6656
rect 185124 6604 185176 6656
rect 324228 6604 324280 6656
rect 447784 6604 447836 6656
rect 40960 6536 41012 6588
rect 183744 6536 183796 6588
rect 325608 6536 325660 6588
rect 451280 6536 451332 6588
rect 37372 6468 37424 6520
rect 182272 6468 182324 6520
rect 326988 6468 327040 6520
rect 454868 6468 454920 6520
rect 33876 6400 33928 6452
rect 180892 6400 180944 6452
rect 186044 6400 186096 6452
rect 233516 6400 233568 6452
rect 328368 6400 328420 6452
rect 458456 6400 458508 6452
rect 30288 6332 30340 6384
rect 179512 6332 179564 6384
rect 182548 6332 182600 6384
rect 232136 6332 232188 6384
rect 329656 6332 329708 6384
rect 462044 6332 462096 6384
rect 26700 6264 26752 6316
rect 178132 6264 178184 6316
rect 178960 6264 179012 6316
rect 230480 6264 230532 6316
rect 329748 6264 329800 6316
rect 465632 6264 465684 6316
rect 8852 6196 8904 6248
rect 172796 6196 172848 6248
rect 175372 6196 175424 6248
rect 229192 6196 229244 6248
rect 331128 6196 331180 6248
rect 469128 6196 469180 6248
rect 4068 6128 4120 6180
rect 171232 6128 171284 6180
rect 171784 6128 171836 6180
rect 227904 6128 227956 6180
rect 332508 6128 332560 6180
rect 472716 6128 472768 6180
rect 132592 6060 132644 6112
rect 215300 6060 215352 6112
rect 318708 6060 318760 6112
rect 433524 6060 433576 6112
rect 136088 5992 136140 6044
rect 216772 5992 216824 6044
rect 318616 5992 318668 6044
rect 429936 5992 429988 6044
rect 139676 5924 139728 5976
rect 217140 5924 217192 5976
rect 317328 5924 317380 5976
rect 426348 5924 426400 5976
rect 143264 5856 143316 5908
rect 218060 5856 218112 5908
rect 315948 5856 316000 5908
rect 422760 5856 422812 5908
rect 146852 5788 146904 5840
rect 219808 5788 219860 5840
rect 314568 5788 314620 5840
rect 419172 5788 419224 5840
rect 150440 5720 150492 5772
rect 221004 5720 221056 5772
rect 313188 5720 313240 5772
rect 415676 5720 415728 5772
rect 159916 5652 159968 5704
rect 224040 5652 224092 5704
rect 311808 5652 311860 5704
rect 412088 5652 412140 5704
rect 164700 5584 164752 5636
rect 226432 5584 226484 5636
rect 310428 5584 310480 5636
rect 408500 5584 408552 5636
rect 168196 5516 168248 5568
rect 227812 5516 227864 5568
rect 309048 5516 309100 5568
rect 404912 5516 404964 5568
rect 65984 5448 66036 5500
rect 192116 5448 192168 5500
rect 288256 5448 288308 5500
rect 341892 5448 341944 5500
rect 357348 5448 357400 5500
rect 544108 5448 544160 5500
rect 62396 5380 62448 5432
rect 190644 5380 190696 5432
rect 286784 5380 286836 5432
rect 340696 5380 340748 5432
rect 358728 5380 358780 5432
rect 547696 5380 547748 5432
rect 58808 5312 58860 5364
rect 189356 5312 189408 5364
rect 208676 5312 208728 5364
rect 241704 5312 241756 5364
rect 289636 5312 289688 5364
rect 345480 5312 345532 5364
rect 360016 5312 360068 5364
rect 551192 5312 551244 5364
rect 55220 5244 55272 5296
rect 187976 5244 188028 5296
rect 205088 5244 205140 5296
rect 240324 5244 240376 5296
rect 288164 5244 288216 5296
rect 344284 5244 344336 5296
rect 361488 5244 361540 5296
rect 554780 5244 554832 5296
rect 51632 5176 51684 5228
rect 187792 5176 187844 5228
rect 201500 5176 201552 5228
rect 238944 5176 238996 5228
rect 289728 5176 289780 5228
rect 347872 5176 347924 5228
rect 362776 5176 362828 5228
rect 558368 5176 558420 5228
rect 48136 5108 48188 5160
rect 186504 5108 186556 5160
rect 198004 5108 198056 5160
rect 237656 5108 237708 5160
rect 291016 5108 291068 5160
rect 351368 5108 351420 5160
rect 362684 5108 362736 5160
rect 561956 5108 562008 5160
rect 17316 5040 17368 5092
rect 175556 5040 175608 5092
rect 194416 5040 194468 5092
rect 236368 5040 236420 5092
rect 292396 5040 292448 5092
rect 354956 5040 355008 5092
rect 364248 5040 364300 5092
rect 565544 5040 565596 5092
rect 12440 4972 12492 5024
rect 174084 4972 174136 5024
rect 190828 4972 190880 5024
rect 234896 4972 234948 5024
rect 293776 4972 293828 5024
rect 358544 4972 358596 5024
rect 365536 4972 365588 5024
rect 569040 4972 569092 5024
rect 7656 4904 7708 4956
rect 172704 4904 172756 4956
rect 187240 4904 187292 4956
rect 233332 4904 233384 4956
rect 295248 4904 295300 4956
rect 362132 4904 362184 4956
rect 366732 4904 366784 4956
rect 572628 4904 572680 4956
rect 2872 4836 2924 4888
rect 169944 4836 169996 4888
rect 174176 4836 174228 4888
rect 229100 4836 229152 4888
rect 296628 4836 296680 4888
rect 365720 4836 365772 4888
rect 368296 4836 368348 4888
rect 576216 4836 576268 4888
rect 1676 4768 1728 4820
rect 169852 4768 169904 4820
rect 170588 4768 170640 4820
rect 228180 4768 228232 4820
rect 298008 4768 298060 4820
rect 369216 4768 369268 4820
rect 369676 4768 369728 4820
rect 579804 4768 579856 4820
rect 69480 4700 69532 4752
rect 193496 4700 193548 4752
rect 286600 4700 286652 4752
rect 338304 4700 338356 4752
rect 355968 4700 356020 4752
rect 540520 4700 540572 4752
rect 127808 4632 127860 4684
rect 212816 4632 212868 4684
rect 286876 4632 286928 4684
rect 337108 4632 337160 4684
rect 354588 4632 354640 4684
rect 536932 4632 536984 4684
rect 144460 4564 144512 4616
rect 219440 4564 219492 4616
rect 285312 4564 285364 4616
rect 334716 4564 334768 4616
rect 353208 4564 353260 4616
rect 533436 4564 533488 4616
rect 148048 4496 148100 4548
rect 220820 4496 220872 4548
rect 283932 4496 283984 4548
rect 331220 4496 331272 4548
rect 351736 4496 351788 4548
rect 529848 4496 529900 4548
rect 151544 4428 151596 4480
rect 220912 4428 220964 4480
rect 285496 4428 285548 4480
rect 333612 4428 333664 4480
rect 351828 4428 351880 4480
rect 526260 4428 526312 4480
rect 155132 4360 155184 4412
rect 222200 4360 222252 4412
rect 284116 4360 284168 4412
rect 330024 4360 330076 4412
rect 350448 4360 350500 4412
rect 522672 4360 522724 4412
rect 158720 4292 158772 4344
rect 223580 4292 223632 4344
rect 282736 4292 282788 4344
rect 327632 4292 327684 4344
rect 348976 4292 349028 4344
rect 519084 4292 519136 4344
rect 163504 4224 163556 4276
rect 224960 4224 225012 4276
rect 281356 4224 281408 4276
rect 324044 4224 324096 4276
rect 347688 4224 347740 4276
rect 515588 4224 515640 4276
rect 167092 4156 167144 4208
rect 226340 4156 226392 4208
rect 277216 4156 277268 4208
rect 61200 4088 61252 4140
rect 186964 4088 187016 4140
rect 199200 4088 199252 4140
rect 203524 4088 203576 4140
rect 211068 4088 211120 4140
rect 211804 4088 211856 4140
rect 214656 4088 214708 4140
rect 215208 4088 215260 4140
rect 217048 4088 217100 4140
rect 218704 4088 218756 4140
rect 221740 4088 221792 4140
rect 245016 4088 245068 4140
rect 257436 4088 257488 4140
rect 257988 4088 258040 4140
rect 258172 4088 258224 4140
rect 258632 4088 258684 4140
rect 259368 4088 259420 4140
rect 259828 4088 259880 4140
rect 261484 4088 261536 4140
rect 262220 4088 262272 4140
rect 54024 4020 54076 4072
rect 185584 4020 185636 4072
rect 206284 4020 206336 4072
rect 211896 4020 211948 4072
rect 215852 4020 215904 4072
rect 240784 4020 240836 4072
rect 241428 4020 241480 4072
rect 261576 4020 261628 4072
rect 264612 4088 264664 4140
rect 269764 4088 269816 4140
rect 272892 4088 272944 4140
rect 263508 4020 263560 4072
rect 270500 4020 270552 4072
rect 14832 3952 14884 4004
rect 17224 3952 17276 4004
rect 43352 3952 43404 4004
rect 183836 3952 183888 4004
rect 213460 3952 213512 4004
rect 234804 3952 234856 4004
rect 247776 3952 247828 4004
rect 267556 3952 267608 4004
rect 276480 4020 276532 4072
rect 276664 4088 276716 4140
rect 277676 4088 277728 4140
rect 279976 4156 280028 4208
rect 320456 4156 320508 4208
rect 346308 4156 346360 4208
rect 512000 4156 512052 4208
rect 279424 4088 279476 4140
rect 282460 4088 282512 4140
rect 283656 4088 283708 4140
rect 272800 3952 272852 4004
rect 42156 3884 42208 3936
rect 183928 3884 183980 3936
rect 195612 3884 195664 3936
rect 225328 3884 225380 3936
rect 226248 3884 226300 3936
rect 233240 3884 233292 3936
rect 233700 3884 233752 3936
rect 240692 3884 240744 3936
rect 241980 3884 242032 3936
rect 249156 3884 249208 3936
rect 268752 3884 268804 3936
rect 285956 3952 286008 4004
rect 286968 4088 287020 4140
rect 306380 4088 306432 4140
rect 352472 4088 352524 4140
rect 460848 4088 460900 4140
rect 469864 4088 469916 4140
rect 550088 4088 550140 4140
rect 310980 4020 311032 4072
rect 311072 4020 311124 4072
rect 316960 4020 317012 4072
rect 345664 4020 345716 4072
rect 453672 4020 453724 4072
rect 474004 4020 474056 4072
rect 557172 4020 557224 4072
rect 314568 3952 314620 4004
rect 316684 3952 316736 4004
rect 328828 3952 328880 4004
rect 330484 3952 330536 4004
rect 439412 3952 439464 4004
rect 475384 3952 475436 4004
rect 564348 3952 564400 4004
rect 283656 3884 283708 3936
rect 285588 3884 285640 3936
rect 287612 3884 287664 3936
rect 24308 3816 24360 3868
rect 31024 3816 31076 3868
rect 36176 3816 36228 3868
rect 182364 3816 182416 3868
rect 192024 3816 192076 3868
rect 235264 3816 235316 3868
rect 242992 3816 243044 3868
rect 265624 3816 265676 3868
rect 25504 3748 25556 3800
rect 32404 3748 32456 3800
rect 34980 3748 35032 3800
rect 181076 3748 181128 3800
rect 193220 3748 193272 3800
rect 236000 3748 236052 3800
rect 246764 3748 246816 3800
rect 254124 3748 254176 3800
rect 267648 3748 267700 3800
rect 287152 3816 287204 3868
rect 278872 3748 278924 3800
rect 280068 3748 280120 3800
rect 318064 3884 318116 3936
rect 337384 3884 337436 3936
rect 467932 3884 467984 3936
rect 478144 3884 478196 3936
rect 571432 3884 571484 3936
rect 16028 3680 16080 3732
rect 24124 3680 24176 3732
rect 29092 3680 29144 3732
rect 179420 3680 179472 3732
rect 189632 3680 189684 3732
rect 234620 3680 234672 3732
rect 243084 3680 243136 3732
rect 243176 3680 243228 3732
rect 251824 3680 251876 3732
rect 262128 3680 262180 3732
rect 268108 3680 268160 3732
rect 270408 3680 270460 3732
rect 278688 3680 278740 3732
rect 20720 3612 20772 3664
rect 176752 3612 176804 3664
rect 188436 3612 188488 3664
rect 234712 3612 234764 3664
rect 239588 3612 239640 3664
rect 250444 3612 250496 3664
rect 266176 3612 266228 3664
rect 281264 3612 281316 3664
rect 281448 3612 281500 3664
rect 321652 3816 321704 3868
rect 333888 3816 333940 3868
rect 475108 3816 475160 3868
rect 477500 3816 477552 3868
rect 478696 3816 478748 3868
rect 480904 3816 480956 3868
rect 578608 3816 578660 3868
rect 287980 3748 288032 3800
rect 335912 3748 335964 3800
rect 336648 3748 336700 3800
rect 482284 3748 482336 3800
rect 520280 3748 520332 3800
rect 521476 3748 521528 3800
rect 339500 3680 339552 3732
rect 360108 3680 360160 3732
rect 553584 3680 553636 3732
rect 288348 3612 288400 3664
rect 343088 3612 343140 3664
rect 362868 3612 362920 3664
rect 560760 3612 560812 3664
rect 19524 3544 19576 3596
rect 176660 3544 176712 3596
rect 183744 3544 183796 3596
rect 231860 3544 231912 3596
rect 6460 3476 6512 3528
rect 10324 3476 10376 3528
rect 11244 3476 11296 3528
rect 173164 3476 173216 3528
rect 184848 3476 184900 3528
rect 236092 3544 236144 3596
rect 244372 3544 244424 3596
rect 245568 3544 245620 3596
rect 263416 3544 263468 3596
rect 269304 3544 269356 3596
rect 270132 3544 270184 3596
rect 290740 3544 290792 3596
rect 291108 3544 291160 3596
rect 350264 3544 350316 3596
rect 365628 3544 365680 3596
rect 567844 3544 567896 3596
rect 236000 3476 236052 3528
rect 249984 3476 250036 3528
rect 251456 3476 251508 3528
rect 252468 3476 252520 3528
rect 266268 3476 266320 3528
rect 10048 3408 10100 3460
rect 172888 3408 172940 3460
rect 181352 3408 181404 3460
rect 27896 3340 27948 3392
rect 28908 3340 28960 3392
rect 32680 3340 32732 3392
rect 35164 3340 35216 3392
rect 39764 3340 39816 3392
rect 42064 3340 42116 3392
rect 70676 3340 70728 3392
rect 71688 3340 71740 3392
rect 38568 3272 38620 3324
rect 68284 3272 68336 3324
rect 188344 3340 188396 3392
rect 77852 3272 77904 3324
rect 78588 3272 78640 3324
rect 81440 3272 81492 3324
rect 82728 3272 82780 3324
rect 191012 3272 191064 3324
rect 45744 3204 45796 3256
rect 71044 3204 71096 3256
rect 84936 3204 84988 3256
rect 85488 3204 85540 3256
rect 57612 3136 57664 3188
rect 82636 3136 82688 3188
rect 192576 3204 192628 3256
rect 196808 3204 196860 3256
rect 204904 3204 204956 3256
rect 209872 3204 209924 3256
rect 226524 3408 226576 3460
rect 227628 3408 227680 3460
rect 232412 3408 232464 3460
rect 232504 3408 232556 3460
rect 249064 3408 249116 3460
rect 249156 3408 249208 3460
rect 251916 3408 251968 3460
rect 263324 3408 263376 3460
rect 271696 3408 271748 3460
rect 272524 3476 272576 3528
rect 275284 3476 275336 3528
rect 291936 3476 291988 3528
rect 292488 3476 292540 3528
rect 353760 3476 353812 3528
rect 368388 3476 368440 3528
rect 575020 3476 575072 3528
rect 231952 3340 232004 3392
rect 245568 3340 245620 3392
rect 250536 3340 250588 3392
rect 267004 3340 267056 3392
rect 274088 3340 274140 3392
rect 274180 3340 274232 3392
rect 293132 3408 293184 3460
rect 293868 3408 293920 3460
rect 297364 3408 297416 3460
rect 301412 3408 301464 3460
rect 357348 3408 357400 3460
rect 358084 3408 358136 3460
rect 369768 3408 369820 3460
rect 582196 3408 582248 3460
rect 88524 3136 88576 3188
rect 89628 3136 89680 3188
rect 50528 3068 50580 3120
rect 77944 3068 77996 3120
rect 79048 3068 79100 3120
rect 86132 3068 86184 3120
rect 192484 3136 192536 3188
rect 207480 3136 207532 3188
rect 208308 3136 208360 3188
rect 218152 3136 218204 3188
rect 239404 3272 239456 3324
rect 250352 3272 250404 3324
rect 255596 3272 255648 3324
rect 268844 3272 268896 3324
rect 280068 3340 280120 3392
rect 277216 3272 277268 3324
rect 277308 3272 277360 3324
rect 309784 3340 309836 3392
rect 312544 3340 312596 3392
rect 313372 3340 313424 3392
rect 93308 3068 93360 3120
rect 193864 3068 193916 3120
rect 200396 3068 200448 3120
rect 201408 3068 201460 3120
rect 202696 3068 202748 3120
rect 209044 3068 209096 3120
rect 224132 3068 224184 3120
rect 243544 3204 243596 3256
rect 253848 3204 253900 3256
rect 256884 3204 256936 3256
rect 275928 3204 275980 3256
rect 307392 3272 307444 3324
rect 309692 3272 309744 3324
rect 325240 3340 325292 3392
rect 341524 3340 341576 3392
rect 446588 3340 446640 3392
rect 494060 3340 494112 3392
rect 495348 3340 495400 3392
rect 502340 3340 502392 3392
rect 503628 3340 503680 3392
rect 326436 3272 326488 3324
rect 327724 3272 327776 3324
rect 417976 3272 418028 3324
rect 302976 3204 303028 3256
rect 306196 3204 306248 3256
rect 322848 3204 322900 3256
rect 340144 3204 340196 3256
rect 425152 3204 425204 3256
rect 228916 3136 228968 3188
rect 247684 3136 247736 3188
rect 271788 3136 271840 3188
rect 95700 3000 95752 3052
rect 96528 3000 96580 3052
rect 96896 3000 96948 3052
rect 102600 3000 102652 3052
rect 102784 3000 102836 3052
rect 103428 3000 103480 3052
rect 103980 3000 104032 3052
rect 104808 3000 104860 3052
rect 106372 3000 106424 3052
rect 107568 3000 107620 3052
rect 111156 3000 111208 3052
rect 111708 3000 111760 3052
rect 46940 2932 46992 2984
rect 71872 2932 71924 2984
rect 84844 2932 84896 2984
rect 88984 2932 89036 2984
rect 89720 2932 89772 2984
rect 95884 2932 95936 2984
rect 100484 2932 100536 2984
rect 195336 3000 195388 3052
rect 222936 3000 222988 3052
rect 229744 3000 229796 3052
rect 113548 2932 113600 2984
rect 114468 2932 114520 2984
rect 120632 2932 120684 2984
rect 121368 2932 121420 2984
rect 64788 2864 64840 2916
rect 106924 2864 106976 2916
rect 114744 2864 114796 2916
rect 75184 2796 75236 2848
rect 75460 2796 75512 2848
rect 86224 2796 86276 2848
rect 97264 2796 97316 2848
rect 107568 2796 107620 2848
rect 195244 2932 195296 2984
rect 195428 2864 195480 2916
rect 220544 2864 220596 2916
rect 238024 3068 238076 3120
rect 273168 3068 273220 3120
rect 300308 3136 300360 3188
rect 301504 3136 301556 3188
rect 299112 3068 299164 3120
rect 300124 3068 300176 3120
rect 305000 3068 305052 3120
rect 231308 3000 231360 3052
rect 248604 3000 248656 3052
rect 252652 3000 252704 3052
rect 254584 3000 254636 3052
rect 274548 3000 274600 3052
rect 280436 3000 280488 3052
rect 295524 3000 295576 3052
rect 298744 3000 298796 3052
rect 302608 3000 302660 3052
rect 326344 3136 326396 3188
rect 410892 3136 410944 3188
rect 305644 3068 305696 3120
rect 308404 3068 308456 3120
rect 323584 3068 323636 3120
rect 403716 3068 403768 3120
rect 308588 3000 308640 3052
rect 319444 3000 319496 3052
rect 360936 3000 360988 3052
rect 432328 3000 432380 3052
rect 121828 2796 121880 2848
rect 122748 2796 122800 2848
rect 124220 2796 124272 2848
rect 125508 2796 125560 2848
rect 125416 2728 125468 2780
rect 196624 2796 196676 2848
rect 227720 2796 227772 2848
rect 244924 2932 244976 2984
rect 270224 2932 270276 2984
rect 289544 2932 289596 2984
rect 303804 2932 303856 2984
rect 305736 2932 305788 2984
rect 319260 2932 319312 2984
rect 322204 2932 322256 2984
rect 396632 2932 396684 2984
rect 269028 2864 269080 2916
rect 288348 2864 288400 2916
rect 290464 2864 290516 2916
rect 297916 2864 297968 2916
rect 304264 2864 304316 2916
rect 315764 2864 315816 2916
rect 334624 2864 334676 2916
rect 382280 2864 382332 2916
rect 382372 2864 382424 2916
rect 383568 2864 383620 2916
rect 390560 2864 390612 2916
rect 391848 2864 391900 2916
rect 268936 2796 268988 2848
rect 284760 2796 284812 2848
rect 283564 2728 283616 2780
rect 294328 2796 294380 2848
rect 302884 2796 302936 2848
rect 312176 2796 312228 2848
rect 345756 2796 345808 2848
rect 389456 2796 389508 2848
rect 291844 892 291896 944
rect 296720 892 296772 944
rect 367100 484 367152 536
rect 368020 484 368072 536
rect 375380 484 375432 536
rect 376392 484 376444 536
rect 376760 484 376812 536
rect 377588 484 377640 536
rect 383660 484 383712 536
rect 384672 484 384724 536
rect 385040 484 385092 536
rect 385868 484 385920 536
rect 391940 484 391992 536
rect 393044 484 393096 536
rect 463700 484 463752 536
rect 464436 484 464488 536
rect 478880 484 478932 536
rect 479892 484 479944 536
rect 485872 484 485924 536
rect 486976 484 487028 536
rect 487160 484 487212 536
rect 488172 484 488224 536
rect 489920 484 489972 536
rect 490564 484 490616 536
rect 495440 484 495492 536
rect 496544 484 496596 536
rect 496820 484 496872 536
rect 497740 484 497792 536
rect 538220 484 538272 536
rect 539324 484 539376 536
<< metal2 >>
rect 8086 703600 8198 704800
rect 24278 703600 24390 704800
rect 40470 703600 40582 704800
rect 56754 703600 56866 704800
rect 72946 703600 73058 704800
rect 89138 703600 89250 704800
rect 105422 703600 105534 704800
rect 121614 703600 121726 704800
rect 137806 703600 137918 704800
rect 154090 703600 154202 704800
rect 170282 703600 170394 704800
rect 186474 703600 186586 704800
rect 202758 703600 202870 704800
rect 218950 703600 219062 704800
rect 235142 703600 235254 704800
rect 251426 703600 251538 704800
rect 267618 703600 267730 704800
rect 283810 703600 283922 704800
rect 300094 703600 300206 704800
rect 316286 703600 316398 704800
rect 332478 703600 332590 704800
rect 348762 703600 348874 704800
rect 364954 703600 365066 704800
rect 381146 703600 381258 704800
rect 397430 703600 397542 704800
rect 413622 703600 413734 704800
rect 429814 703600 429926 704800
rect 446098 703600 446210 704800
rect 462290 703600 462402 704800
rect 478482 703600 478594 704800
rect 494766 703610 494878 704800
rect 494766 703600 494928 703610
rect 510958 703600 511070 704800
rect 527150 703600 527262 704800
rect 543434 703600 543546 704800
rect 559626 703600 559738 704800
rect 575818 703600 575930 704800
rect 8128 700330 8156 703600
rect 24320 700466 24348 703600
rect 40512 700534 40540 703600
rect 72988 700670 73016 703600
rect 89180 700806 89208 703600
rect 105464 700874 105492 703600
rect 137848 701010 137876 703600
rect 137836 701004 137888 701010
rect 137836 700946 137888 700952
rect 105452 700868 105504 700874
rect 105452 700810 105504 700816
rect 89168 700800 89220 700806
rect 89168 700742 89220 700748
rect 72976 700664 73028 700670
rect 72976 700606 73028 700612
rect 40500 700528 40552 700534
rect 40500 700470 40552 700476
rect 24308 700460 24360 700466
rect 24308 700402 24360 700408
rect 8116 700324 8168 700330
rect 8116 700266 8168 700272
rect 154132 700194 154160 703600
rect 154120 700188 154172 700194
rect 154120 700130 154172 700136
rect 170324 700126 170352 703600
rect 170312 700120 170364 700126
rect 170312 700062 170364 700068
rect 202800 699990 202828 703600
rect 202788 699984 202840 699990
rect 202788 699926 202840 699932
rect 218992 699854 219020 703600
rect 218980 699848 219032 699854
rect 218980 699790 219032 699796
rect 235184 699786 235212 703600
rect 262128 700936 262180 700942
rect 262128 700878 262180 700884
rect 255228 700732 255280 700738
rect 255228 700674 255280 700680
rect 249708 700392 249760 700398
rect 249708 700334 249760 700340
rect 252374 700360 252430 700369
rect 235172 699780 235224 699786
rect 235172 699722 235224 699728
rect 245568 696992 245620 696998
rect 245568 696934 245620 696940
rect 3514 682272 3570 682281
rect 3514 682207 3570 682216
rect 3528 681766 3556 682207
rect 3516 681760 3568 681766
rect 3516 681702 3568 681708
rect 242808 673532 242860 673538
rect 242808 673474 242860 673480
rect 3422 667992 3478 668001
rect 3422 667927 3424 667936
rect 3476 667927 3478 667936
rect 3424 667898 3476 667904
rect 3054 653576 3110 653585
rect 3054 653511 3110 653520
rect 3068 652798 3096 653511
rect 3056 652792 3108 652798
rect 3056 652734 3108 652740
rect 240048 650072 240100 650078
rect 240048 650014 240100 650020
rect 238668 626612 238720 626618
rect 238668 626554 238720 626560
rect 3422 624880 3478 624889
rect 3422 624815 3478 624824
rect 3436 623830 3464 624815
rect 3424 623824 3476 623830
rect 3424 623766 3476 623772
rect 3422 610464 3478 610473
rect 3422 610399 3478 610408
rect 3436 610026 3464 610399
rect 3424 610020 3476 610026
rect 3424 609962 3476 609968
rect 234528 603152 234580 603158
rect 234528 603094 234580 603100
rect 3238 596048 3294 596057
rect 3238 595983 3294 595992
rect 3252 594862 3280 595983
rect 3240 594856 3292 594862
rect 3240 594798 3292 594804
rect 233148 579692 233200 579698
rect 233148 579634 233200 579640
rect 3422 567352 3478 567361
rect 3422 567287 3478 567296
rect 3436 567254 3464 567287
rect 3424 567248 3476 567254
rect 3424 567190 3476 567196
rect 229008 556232 229060 556238
rect 229008 556174 229060 556180
rect 3146 553072 3202 553081
rect 3146 553007 3202 553016
rect 3160 552090 3188 553007
rect 3148 552084 3200 552090
rect 3148 552026 3200 552032
rect 3422 538656 3478 538665
rect 3422 538591 3478 538600
rect 3436 538286 3464 538591
rect 3424 538280 3476 538286
rect 3424 538222 3476 538228
rect 227628 532772 227680 532778
rect 227628 532714 227680 532720
rect 196806 523016 196862 523025
rect 196806 522951 196862 522960
rect 209686 523016 209742 523025
rect 222014 523016 222070 523025
rect 209686 522951 209742 522960
rect 219072 522980 219124 522986
rect 190000 522844 190052 522850
rect 190000 522786 190052 522792
rect 2964 522776 3016 522782
rect 2964 522718 3016 522724
rect 184846 522744 184902 522753
rect 2976 509969 3004 522718
rect 4712 522708 4764 522714
rect 184846 522679 184902 522688
rect 4712 522650 4764 522656
rect 3056 522640 3108 522646
rect 3056 522582 3108 522588
rect 2962 509960 3018 509969
rect 2962 509895 3018 509904
rect 2780 495576 2832 495582
rect 2778 495544 2780 495553
rect 2832 495544 2834 495553
rect 2778 495479 2834 495488
rect 3068 481137 3096 522582
rect 3148 522572 3200 522578
rect 3148 522514 3200 522520
rect 3054 481128 3110 481137
rect 3054 481063 3110 481072
rect 3056 452464 3108 452470
rect 3054 452432 3056 452441
rect 3108 452432 3110 452441
rect 3054 452367 3110 452376
rect 3160 438025 3188 522514
rect 3240 522504 3292 522510
rect 3240 522446 3292 522452
rect 3146 438016 3202 438025
rect 3146 437951 3202 437960
rect 3148 424108 3200 424114
rect 3148 424050 3200 424056
rect 3160 423745 3188 424050
rect 3146 423736 3202 423745
rect 3146 423671 3202 423680
rect 3252 395049 3280 522446
rect 4068 522300 4120 522306
rect 4068 522242 4120 522248
rect 3884 521892 3936 521898
rect 3884 521834 3936 521840
rect 3792 521824 3844 521830
rect 3792 521766 3844 521772
rect 3332 519376 3384 519382
rect 3332 519318 3384 519324
rect 3238 395040 3294 395049
rect 3238 394975 3294 394984
rect 2780 380656 2832 380662
rect 2778 380624 2780 380633
rect 2832 380624 2834 380633
rect 2778 380559 2834 380568
rect 2780 366988 2832 366994
rect 2780 366930 2832 366936
rect 2792 366217 2820 366930
rect 2778 366208 2834 366217
rect 2778 366143 2834 366152
rect 3344 337521 3372 519318
rect 3700 519240 3752 519246
rect 3700 519182 3752 519188
rect 3424 519036 3476 519042
rect 3424 518978 3476 518984
rect 3330 337512 3386 337521
rect 3330 337447 3386 337456
rect 3148 324216 3200 324222
rect 3148 324158 3200 324164
rect 3160 323105 3188 324158
rect 3146 323096 3202 323105
rect 3146 323031 3202 323040
rect 3332 280152 3384 280158
rect 3330 280120 3332 280129
rect 3384 280120 3386 280129
rect 3330 280055 3386 280064
rect 2780 266076 2832 266082
rect 2780 266018 2832 266024
rect 2792 265713 2820 266018
rect 2778 265704 2834 265713
rect 2778 265639 2834 265648
rect 3332 237380 3384 237386
rect 3332 237322 3384 237328
rect 3344 237017 3372 237322
rect 3330 237008 3386 237017
rect 3330 236943 3386 236952
rect 3148 194540 3200 194546
rect 3148 194482 3200 194488
rect 3160 193905 3188 194482
rect 3146 193896 3202 193905
rect 3146 193831 3202 193840
rect 2780 165504 2832 165510
rect 2780 165446 2832 165452
rect 2792 165073 2820 165446
rect 2778 165064 2834 165073
rect 2778 164999 2834 165008
rect 3332 151768 3384 151774
rect 3332 151710 3384 151716
rect 3344 150793 3372 151710
rect 3330 150784 3386 150793
rect 3330 150719 3386 150728
rect 2780 136536 2832 136542
rect 2780 136478 2832 136484
rect 2792 136377 2820 136478
rect 2778 136368 2834 136377
rect 2778 136303 2834 136312
rect 2780 122324 2832 122330
rect 2780 122266 2832 122272
rect 2792 122097 2820 122266
rect 2778 122088 2834 122097
rect 2778 122023 2834 122032
rect 3332 108996 3384 109002
rect 3332 108938 3384 108944
rect 3344 107681 3372 108938
rect 3330 107672 3386 107681
rect 3330 107607 3386 107616
rect 3436 78985 3464 518978
rect 3606 518800 3662 518809
rect 3606 518735 3662 518744
rect 3516 518288 3568 518294
rect 3516 518230 3568 518236
rect 3528 93265 3556 518230
rect 3620 179489 3648 518735
rect 3712 208185 3740 519182
rect 3804 222601 3832 521766
rect 3896 251297 3924 521834
rect 3976 519308 4028 519314
rect 3976 519250 4028 519256
rect 3988 294409 4016 519250
rect 4080 308825 4108 522242
rect 4724 495582 4752 522650
rect 174542 522608 174598 522617
rect 174542 522543 174598 522552
rect 28262 522472 28318 522481
rect 5448 522436 5500 522442
rect 28262 522407 28318 522416
rect 5448 522378 5500 522384
rect 4894 522336 4950 522345
rect 4894 522271 4950 522280
rect 4804 518968 4856 518974
rect 4804 518910 4856 518916
rect 4712 495576 4764 495582
rect 4712 495518 4764 495524
rect 4066 308816 4122 308825
rect 4066 308751 4122 308760
rect 3974 294400 4030 294409
rect 3974 294335 4030 294344
rect 3882 251288 3938 251297
rect 3882 251223 3938 251232
rect 3790 222592 3846 222601
rect 3790 222527 3846 222536
rect 3698 208176 3754 208185
rect 3698 208111 3754 208120
rect 3606 179480 3662 179489
rect 3606 179415 3662 179424
rect 3514 93256 3570 93265
rect 3514 93191 3570 93200
rect 3422 78976 3478 78985
rect 3422 78911 3478 78920
rect 754 64832 810 64841
rect 754 64767 810 64776
rect 768 64569 796 64767
rect 754 64560 810 64569
rect 754 64495 810 64504
rect 2780 50176 2832 50182
rect 2778 50144 2780 50153
rect 2832 50144 2834 50153
rect 2778 50079 2834 50088
rect 4816 35902 4844 518910
rect 4908 50182 4936 522271
rect 5264 522028 5316 522034
rect 5264 521970 5316 521976
rect 5080 521756 5132 521762
rect 5080 521698 5132 521704
rect 4988 519104 5040 519110
rect 4988 519046 5040 519052
rect 5000 122330 5028 519046
rect 5092 136542 5120 521698
rect 5172 519172 5224 519178
rect 5172 519114 5224 519120
rect 5184 165510 5212 519114
rect 5276 266082 5304 521970
rect 5356 519444 5408 519450
rect 5356 519386 5408 519392
rect 5368 366994 5396 519386
rect 5460 380662 5488 522378
rect 6184 522368 6236 522374
rect 6184 522310 6236 522316
rect 5448 380656 5500 380662
rect 5448 380598 5500 380604
rect 5356 366988 5408 366994
rect 5356 366930 5408 366936
rect 6196 324222 6224 522310
rect 19984 522232 20036 522238
rect 19984 522174 20036 522180
rect 10324 522164 10376 522170
rect 10324 522106 10376 522112
rect 6368 519512 6420 519518
rect 6368 519454 6420 519460
rect 6274 517576 6330 517585
rect 6274 517511 6330 517520
rect 6288 424114 6316 517511
rect 6380 452470 6408 519454
rect 6368 452464 6420 452470
rect 6368 452406 6420 452412
rect 6276 424108 6328 424114
rect 6276 424050 6328 424056
rect 6184 324216 6236 324222
rect 6184 324158 6236 324164
rect 10336 280158 10364 522106
rect 13084 522096 13136 522102
rect 13084 522038 13136 522044
rect 12530 517712 12586 517721
rect 12360 517670 12530 517698
rect 12360 517585 12388 517670
rect 12530 517647 12586 517656
rect 12346 517576 12402 517585
rect 12346 517511 12402 517520
rect 10324 280152 10376 280158
rect 10324 280094 10376 280100
rect 5264 266076 5316 266082
rect 5264 266018 5316 266024
rect 13096 237386 13124 522038
rect 13084 237380 13136 237386
rect 13084 237322 13136 237328
rect 17224 217320 17276 217326
rect 10322 217288 10378 217297
rect 17224 217262 17276 217268
rect 10322 217223 10378 217232
rect 5172 165504 5224 165510
rect 5172 165446 5224 165452
rect 5080 136536 5132 136542
rect 5080 136478 5132 136484
rect 4988 122324 5040 122330
rect 4988 122266 5040 122272
rect 4896 50176 4948 50182
rect 4896 50118 4948 50124
rect 2780 35896 2832 35902
rect 2778 35864 2780 35873
rect 4804 35896 4856 35902
rect 2832 35864 2834 35873
rect 4804 35838 4856 35844
rect 2778 35799 2834 35808
rect 478 21992 534 22001
rect 478 21927 534 21936
rect 492 21457 520 21927
rect 478 21448 534 21457
rect 478 21383 534 21392
rect 2962 10296 3018 10305
rect 2962 10231 3018 10240
rect 2976 7177 3004 10231
rect 2962 7168 3018 7177
rect 2962 7103 3018 7112
rect 8852 6248 8904 6254
rect 8852 6190 8904 6196
rect 4068 6180 4120 6186
rect 4068 6122 4120 6128
rect 2872 4888 2924 4894
rect 570 4856 626 4865
rect 2872 4830 2924 4836
rect 570 4791 626 4800
rect 1676 4820 1728 4826
rect 584 400 612 4791
rect 1676 4762 1728 4768
rect 1688 400 1716 4762
rect 2884 400 2912 4830
rect 4080 400 4108 6122
rect 7656 4956 7708 4962
rect 7656 4898 7708 4904
rect 6460 3528 6512 3534
rect 6460 3470 6512 3476
rect 5262 3360 5318 3369
rect 5262 3295 5318 3304
rect 5276 400 5304 3295
rect 6472 400 6500 3470
rect 7668 400 7696 4898
rect 8864 400 8892 6190
rect 10336 3534 10364 217223
rect 13636 8968 13688 8974
rect 13636 8910 13688 8916
rect 12440 5024 12492 5030
rect 12440 4966 12492 4972
rect 10324 3528 10376 3534
rect 10324 3470 10376 3476
rect 11244 3528 11296 3534
rect 11244 3470 11296 3476
rect 10048 3460 10100 3466
rect 10048 3402 10100 3408
rect 10060 400 10088 3402
rect 11256 400 11284 3470
rect 12452 400 12480 4966
rect 13648 400 13676 8910
rect 17236 4010 17264 217262
rect 19996 194546 20024 522174
rect 21364 521960 21416 521966
rect 21364 521902 21416 521908
rect 19984 194540 20036 194546
rect 19984 194482 20036 194488
rect 21376 151774 21404 521902
rect 22006 517712 22062 517721
rect 22062 517670 22232 517698
rect 22006 517647 22062 517656
rect 22204 517585 22232 517670
rect 27620 517608 27672 517614
rect 22190 517576 22246 517585
rect 22190 517511 22246 517520
rect 27618 517576 27620 517585
rect 27672 517576 27674 517585
rect 27618 517511 27674 517520
rect 24124 217388 24176 217394
rect 24124 217330 24176 217336
rect 21364 151768 21416 151774
rect 21364 151710 21416 151716
rect 23112 9104 23164 9110
rect 23112 9046 23164 9052
rect 18328 9036 18380 9042
rect 18328 8978 18380 8984
rect 17316 5092 17368 5098
rect 17316 5034 17368 5040
rect 14832 4004 14884 4010
rect 14832 3946 14884 3952
rect 17224 4004 17276 4010
rect 17224 3946 17276 3952
rect 14844 400 14872 3946
rect 16028 3732 16080 3738
rect 16028 3674 16080 3680
rect 16040 400 16068 3674
rect 17328 2530 17356 5034
rect 17236 2502 17356 2530
rect 17236 400 17264 2502
rect 18340 400 18368 8978
rect 21914 6216 21970 6225
rect 21914 6151 21970 6160
rect 20720 3664 20772 3670
rect 20720 3606 20772 3612
rect 19524 3596 19576 3602
rect 19524 3538 19576 3544
rect 19536 400 19564 3538
rect 20732 400 20760 3606
rect 21928 400 21956 6151
rect 23124 400 23152 9046
rect 24136 3738 24164 217330
rect 28276 109002 28304 522407
rect 174556 519874 174584 522543
rect 181350 522064 181406 522073
rect 181350 521999 181406 522008
rect 177946 521928 178002 521937
rect 177946 521863 178002 521872
rect 176198 521792 176254 521801
rect 176198 521727 176254 521736
rect 176212 519874 176240 521727
rect 177960 519874 177988 521863
rect 181364 519874 181392 521999
rect 183192 520328 183244 520334
rect 183192 520270 183244 520276
rect 183204 519874 183232 520270
rect 184860 519874 184888 522679
rect 186136 521688 186188 521694
rect 186136 521630 186188 521636
rect 186148 520010 186176 521630
rect 188160 520396 188212 520402
rect 188160 520338 188212 520344
rect 186148 519982 186254 520010
rect 188172 519874 188200 520338
rect 190012 519874 190040 522786
rect 190642 522744 190698 522753
rect 190642 522679 190698 522688
rect 190656 522209 190684 522679
rect 190642 522200 190698 522209
rect 190642 522135 190698 522144
rect 191654 520296 191710 520305
rect 191654 520231 191710 520240
rect 191668 519874 191696 520231
rect 196820 519874 196848 522951
rect 201958 522880 202014 522889
rect 201958 522815 202014 522824
rect 201972 519874 202000 522815
rect 209700 522753 209728 522951
rect 222014 522951 222070 522960
rect 219072 522922 219124 522928
rect 213828 522912 213880 522918
rect 213828 522854 213880 522860
rect 209686 522744 209742 522753
rect 209686 522679 209742 522688
rect 212080 520668 212132 520674
rect 212080 520610 212132 520616
rect 208768 520600 208820 520606
rect 208768 520542 208820 520548
rect 206928 520532 206980 520538
rect 206928 520474 206980 520480
rect 203616 520464 203668 520470
rect 203616 520406 203668 520412
rect 203628 519874 203656 520406
rect 206940 519874 206968 520474
rect 208780 519874 208808 520542
rect 212092 519874 212120 520610
rect 213840 519874 213868 522854
rect 217232 520736 217284 520742
rect 217232 520678 217284 520684
rect 217244 519874 217272 520678
rect 219084 519874 219112 522922
rect 220728 520804 220780 520810
rect 220728 520746 220780 520752
rect 220740 519874 220768 520746
rect 222028 520010 222056 522951
rect 224224 520872 224276 520878
rect 224224 520814 224276 520820
rect 222028 519982 222134 520010
rect 224236 519874 224264 520814
rect 227640 519874 227668 532714
rect 229020 519874 229048 556174
rect 231768 545148 231820 545154
rect 231768 545090 231820 545096
rect 231780 526522 231808 545090
rect 233160 526522 233188 579634
rect 234540 526522 234568 603094
rect 235908 592068 235960 592074
rect 235908 592010 235960 592016
rect 235920 526522 235948 592010
rect 238680 526522 238708 626554
rect 230480 526516 230532 526522
rect 230480 526458 230532 526464
rect 231768 526516 231820 526522
rect 231768 526458 231820 526464
rect 231860 526516 231912 526522
rect 231860 526458 231912 526464
rect 233148 526516 233200 526522
rect 233148 526458 233200 526464
rect 233240 526516 233292 526522
rect 233240 526458 233292 526464
rect 234528 526516 234580 526522
rect 234528 526458 234580 526464
rect 234620 526516 234672 526522
rect 234620 526458 234672 526464
rect 235908 526516 235960 526522
rect 235908 526458 235960 526464
rect 237380 526516 237432 526522
rect 237380 526458 237432 526464
rect 238668 526516 238720 526522
rect 238668 526458 238720 526464
rect 230492 520010 230520 526458
rect 230492 519982 230690 520010
rect 174294 519846 174584 519874
rect 175950 519846 176240 519874
rect 177698 519846 177988 519874
rect 181102 519846 181392 519874
rect 182850 519846 183232 519874
rect 184506 519846 184888 519874
rect 187910 519846 188200 519874
rect 189658 519846 190040 519874
rect 191314 519846 191696 519874
rect 196466 519846 196848 519874
rect 201618 519846 202000 519874
rect 203366 519846 203656 519874
rect 206770 519846 206968 519874
rect 208426 519846 208808 519874
rect 211830 519846 212120 519874
rect 213578 519846 213868 519874
rect 216982 519846 217272 519874
rect 218730 519846 219112 519874
rect 220386 519846 220768 519874
rect 223882 519846 224264 519874
rect 227286 519846 227668 519874
rect 228942 519846 229048 519874
rect 231872 519874 231900 526458
rect 233252 519874 233280 526458
rect 234632 520282 234660 526458
rect 234632 520254 235488 520282
rect 235460 520010 235488 520254
rect 237392 520010 237420 526458
rect 240060 520146 240088 650014
rect 241428 638988 241480 638994
rect 241428 638930 241480 638936
rect 241440 520146 241468 638930
rect 239600 520118 240088 520146
rect 241256 520118 241468 520146
rect 235460 519982 235842 520010
rect 237392 519982 237498 520010
rect 239600 519874 239628 520118
rect 241256 519874 241284 520118
rect 242820 519874 242848 673474
rect 245580 520146 245608 696934
rect 246948 685908 247000 685914
rect 246948 685850 247000 685856
rect 246960 520146 246988 685850
rect 248144 523728 248196 523734
rect 248144 523670 248196 523676
rect 244660 520118 245608 520146
rect 246316 520118 246988 520146
rect 244660 519874 244688 520118
rect 246316 519874 246344 520118
rect 248156 519874 248184 523670
rect 249720 519874 249748 700334
rect 252374 700295 252430 700304
rect 252388 688650 252416 700295
rect 252296 688634 252416 688650
rect 252284 688628 252416 688634
rect 252336 688622 252416 688628
rect 252468 688628 252520 688634
rect 252284 688570 252336 688576
rect 252468 688570 252520 688576
rect 252296 688539 252324 688570
rect 252480 685846 252508 688570
rect 252468 685840 252520 685846
rect 252468 685782 252520 685788
rect 252376 676252 252428 676258
rect 252376 676194 252428 676200
rect 252388 669338 252416 676194
rect 252296 669322 252416 669338
rect 252284 669316 252416 669322
rect 252336 669310 252416 669316
rect 252468 669316 252520 669322
rect 252284 669258 252336 669264
rect 252468 669258 252520 669264
rect 252296 669227 252324 669258
rect 252480 666534 252508 669258
rect 252468 666528 252520 666534
rect 252468 666470 252520 666476
rect 252376 656940 252428 656946
rect 252376 656882 252428 656888
rect 252388 650026 252416 656882
rect 252296 650010 252416 650026
rect 252284 650004 252416 650010
rect 252336 649998 252416 650004
rect 252468 650004 252520 650010
rect 252284 649946 252336 649952
rect 252468 649946 252520 649952
rect 252296 649915 252324 649946
rect 252480 647222 252508 649946
rect 252468 647216 252520 647222
rect 252468 647158 252520 647164
rect 252376 637628 252428 637634
rect 252376 637570 252428 637576
rect 252388 630714 252416 637570
rect 252296 630686 252416 630714
rect 252296 630578 252324 630686
rect 252296 630550 252416 630578
rect 252388 621058 252416 630550
rect 252388 621030 252508 621058
rect 252480 620922 252508 621030
rect 252388 620894 252508 620922
rect 252388 611402 252416 620894
rect 252296 611374 252416 611402
rect 252296 611266 252324 611374
rect 252296 611238 252416 611266
rect 252388 601746 252416 611238
rect 252388 601718 252508 601746
rect 252480 601610 252508 601718
rect 252388 601582 252508 601610
rect 252388 592090 252416 601582
rect 252296 592062 252416 592090
rect 252296 591954 252324 592062
rect 252296 591926 252416 591954
rect 252388 582434 252416 591926
rect 252388 582406 252508 582434
rect 252480 582298 252508 582406
rect 252388 582270 252508 582298
rect 252388 572778 252416 582270
rect 252296 572750 252416 572778
rect 252296 572642 252324 572750
rect 252296 572614 252416 572642
rect 252388 563122 252416 572614
rect 252388 563094 252508 563122
rect 252480 562986 252508 563094
rect 252388 562958 252508 562986
rect 252388 553466 252416 562958
rect 252296 553438 252416 553466
rect 252296 553330 252324 553438
rect 252296 553302 252416 553330
rect 252388 543810 252416 553302
rect 252388 543782 252508 543810
rect 252480 543674 252508 543782
rect 252388 543646 252508 543674
rect 252388 534138 252416 543646
rect 251824 534132 251876 534138
rect 251824 534074 251876 534080
rect 252376 534132 252428 534138
rect 252376 534074 252428 534080
rect 251836 528578 251864 534074
rect 251744 528550 251864 528578
rect 251744 520146 251772 528550
rect 253112 523796 253164 523802
rect 253112 523738 253164 523744
rect 251468 520118 251772 520146
rect 251468 519874 251496 520118
rect 253124 519874 253152 523738
rect 255240 520146 255268 700674
rect 256608 700596 256660 700602
rect 256608 700538 256660 700544
rect 254964 520118 255268 520146
rect 254964 519874 254992 520118
rect 256620 519874 256648 700538
rect 260748 700256 260800 700262
rect 260748 700198 260800 700204
rect 257988 617568 258040 617574
rect 257988 617510 258040 617516
rect 258000 520146 258028 617510
rect 260760 520146 260788 700198
rect 262140 520146 262168 700878
rect 267660 700058 267688 703600
rect 280160 701004 280212 701010
rect 280160 700946 280212 700952
rect 277400 700120 277452 700126
rect 277400 700062 277452 700068
rect 279424 700120 279476 700126
rect 279424 700062 279476 700068
rect 267648 700052 267700 700058
rect 267648 699994 267700 700000
rect 269120 700052 269172 700058
rect 269120 699994 269172 700000
rect 264888 699916 264940 699922
rect 264888 699858 264940 699864
rect 263324 523932 263376 523938
rect 263324 523874 263376 523880
rect 258000 520118 258120 520146
rect 258092 519874 258120 520118
rect 260116 520118 260788 520146
rect 261772 520118 262168 520146
rect 260116 519874 260144 520118
rect 261772 519874 261800 520118
rect 263336 519874 263364 523874
rect 264900 519874 264928 699858
rect 267648 699712 267700 699718
rect 267648 699654 267700 699660
rect 267660 688770 267688 699654
rect 269132 698306 269160 699994
rect 274640 699984 274692 699990
rect 274640 699926 274692 699932
rect 273260 699780 273312 699786
rect 273260 699722 273312 699728
rect 271788 699712 271840 699718
rect 271788 699654 271840 699660
rect 269132 698278 269344 698306
rect 269316 695502 269344 698278
rect 269304 695496 269356 695502
rect 269304 695438 269356 695444
rect 267648 688764 267700 688770
rect 267648 688706 267700 688712
rect 267556 685976 267608 685982
rect 267556 685918 267608 685924
rect 269212 685976 269264 685982
rect 269212 685918 269264 685924
rect 267568 684486 267596 685918
rect 269224 684486 269252 685918
rect 267556 684480 267608 684486
rect 267556 684422 267608 684428
rect 269212 684480 269264 684486
rect 269212 684422 269264 684428
rect 267648 682984 267700 682990
rect 267648 682926 267700 682932
rect 267660 674830 267688 682926
rect 269304 676252 269356 676258
rect 269304 676194 269356 676200
rect 267648 674824 267700 674830
rect 267648 674766 267700 674772
rect 269316 669390 269344 676194
rect 269304 669384 269356 669390
rect 269304 669326 269356 669332
rect 269396 669248 269448 669254
rect 269396 669190 269448 669196
rect 267372 665304 267424 665310
rect 267372 665246 267424 665252
rect 267384 665174 267412 665246
rect 267372 665168 267424 665174
rect 267372 665110 267424 665116
rect 269408 663746 269436 669190
rect 269396 663740 269448 663746
rect 269396 663682 269448 663688
rect 267556 659592 267608 659598
rect 267556 659534 267608 659540
rect 267568 650214 267596 659534
rect 267556 650208 267608 650214
rect 267556 650150 267608 650156
rect 269396 649936 269448 649942
rect 269396 649878 269448 649884
rect 267464 645924 267516 645930
rect 267464 645866 267516 645872
rect 267476 645833 267504 645866
rect 267462 645824 267518 645833
rect 267462 645759 267518 645768
rect 269408 640422 269436 649878
rect 269396 640416 269448 640422
rect 269396 640358 269448 640364
rect 269304 640280 269356 640286
rect 267554 640248 267610 640257
rect 269304 640222 269356 640228
rect 267554 640183 267610 640192
rect 267568 630902 267596 640183
rect 267556 630896 267608 630902
rect 267556 630838 267608 630844
rect 267464 626680 267516 626686
rect 267464 626622 267516 626628
rect 267476 623150 267504 626622
rect 267464 623144 267516 623150
rect 267464 623086 267516 623092
rect 267556 623144 267608 623150
rect 267556 623086 267608 623092
rect 267568 611402 267596 623086
rect 269316 611454 269344 640222
rect 269304 611448 269356 611454
rect 267568 611374 267688 611402
rect 269304 611390 269356 611396
rect 267660 611266 267688 611374
rect 267476 611238 267688 611266
rect 269304 611312 269356 611318
rect 269304 611254 269356 611260
rect 267476 601746 267504 611238
rect 267384 601718 267504 601746
rect 269316 601730 269344 611254
rect 269120 601724 269172 601730
rect 267384 592142 267412 601718
rect 269120 601666 269172 601672
rect 269304 601724 269356 601730
rect 269304 601666 269356 601672
rect 269132 598942 269160 601666
rect 269120 598936 269172 598942
rect 269120 598878 269172 598884
rect 267372 592136 267424 592142
rect 267372 592078 267424 592084
rect 267280 589416 267332 589422
rect 267280 589358 267332 589364
rect 267292 582418 267320 589358
rect 269212 589348 269264 589354
rect 269212 589290 269264 589296
rect 269224 587858 269252 589290
rect 269212 587852 269264 587858
rect 269212 587794 269264 587800
rect 267280 582412 267332 582418
rect 267280 582354 267332 582360
rect 269304 582412 269356 582418
rect 269304 582354 269356 582360
rect 267372 582276 267424 582282
rect 267372 582218 267424 582224
rect 267384 578241 267412 582218
rect 269316 578241 269344 582354
rect 267370 578232 267426 578241
rect 267370 578167 267426 578176
rect 267554 578232 267610 578241
rect 267554 578167 267610 578176
rect 269118 578232 269174 578241
rect 269118 578167 269174 578176
rect 269302 578232 269358 578241
rect 269302 578167 269358 578176
rect 267568 568596 267596 578167
rect 269132 568614 269160 578167
rect 267384 568585 267596 568596
rect 269120 568608 269172 568614
rect 267370 568576 267610 568585
rect 267426 568568 267554 568576
rect 267370 568511 267426 568520
rect 269120 568550 269172 568556
rect 269396 568608 269448 568614
rect 269396 568550 269448 568556
rect 267554 568511 267610 568520
rect 267568 562970 267596 568511
rect 269408 563174 269436 568550
rect 269396 563168 269448 563174
rect 269396 563110 269448 563116
rect 269304 563032 269356 563038
rect 269304 562974 269356 562980
rect 267372 562964 267424 562970
rect 267372 562906 267424 562912
rect 267556 562964 267608 562970
rect 267556 562906 267608 562912
rect 267384 553330 267412 562906
rect 269316 553330 269344 562974
rect 267384 553302 267504 553330
rect 267476 543810 267504 553302
rect 269224 553302 269344 553330
rect 269224 548894 269252 553302
rect 269212 548888 269264 548894
rect 269212 548830 269264 548836
rect 269488 548888 269540 548894
rect 269488 548830 269540 548836
rect 267476 543782 267596 543810
rect 267568 531350 267596 543782
rect 269500 540977 269528 548830
rect 269302 540968 269358 540977
rect 269302 540903 269358 540912
rect 269486 540968 269542 540977
rect 269486 540903 269542 540912
rect 269316 531350 269344 540903
rect 267188 531344 267240 531350
rect 267002 531312 267058 531321
rect 267002 531247 267058 531256
rect 267186 531312 267188 531321
rect 267556 531344 267608 531350
rect 267240 531312 267242 531321
rect 267556 531286 267608 531292
rect 269304 531344 269356 531350
rect 269304 531286 269356 531292
rect 269580 531344 269632 531350
rect 269580 531286 269632 531292
rect 267186 531247 267242 531256
rect 267016 519874 267044 531247
rect 269592 526402 269620 531286
rect 269408 526374 269620 526402
rect 268568 523864 268620 523870
rect 268568 523806 268620 523812
rect 268580 519874 268608 523806
rect 269408 520010 269436 526374
rect 269408 519982 269974 520010
rect 271800 519874 271828 699654
rect 273272 520010 273300 699722
rect 274652 520010 274680 699926
rect 276020 699848 276072 699854
rect 276020 699790 276072 699796
rect 276032 692730 276060 699790
rect 276032 692702 276244 692730
rect 276216 683194 276244 692702
rect 276020 683188 276072 683194
rect 276020 683130 276072 683136
rect 276204 683188 276256 683194
rect 276204 683130 276256 683136
rect 276032 669322 276060 683130
rect 276020 669316 276072 669322
rect 276020 669258 276072 669264
rect 276204 669316 276256 669322
rect 276204 669258 276256 669264
rect 276216 666534 276244 669258
rect 276204 666528 276256 666534
rect 276204 666470 276256 666476
rect 276112 656940 276164 656946
rect 276112 656882 276164 656888
rect 276124 650026 276152 656882
rect 276124 649998 276244 650026
rect 276216 644502 276244 649998
rect 276020 644496 276072 644502
rect 276020 644438 276072 644444
rect 276204 644496 276256 644502
rect 276204 644438 276256 644444
rect 276032 640234 276060 644438
rect 276032 640206 276152 640234
rect 276124 630714 276152 640206
rect 276124 630686 276244 630714
rect 276216 611386 276244 630686
rect 276020 611380 276072 611386
rect 276020 611322 276072 611328
rect 276204 611380 276256 611386
rect 276204 611322 276256 611328
rect 276032 611266 276060 611322
rect 276032 611238 276152 611266
rect 276124 601798 276152 611238
rect 276112 601792 276164 601798
rect 276112 601734 276164 601740
rect 276204 601724 276256 601730
rect 276204 601666 276256 601672
rect 276216 598942 276244 601666
rect 276204 598936 276256 598942
rect 276204 598878 276256 598884
rect 276204 592000 276256 592006
rect 276204 591942 276256 591948
rect 276216 589286 276244 591942
rect 276204 589280 276256 589286
rect 276204 589222 276256 589228
rect 276204 582276 276256 582282
rect 276204 582218 276256 582224
rect 276216 572762 276244 582218
rect 276020 572756 276072 572762
rect 276020 572698 276072 572704
rect 276204 572756 276256 572762
rect 276204 572698 276256 572704
rect 276032 572642 276060 572698
rect 276032 572614 276152 572642
rect 276124 563122 276152 572614
rect 276124 563094 276244 563122
rect 276216 560266 276244 563094
rect 276124 560238 276244 560266
rect 276124 550662 276152 560238
rect 276020 550656 276072 550662
rect 276018 550624 276020 550633
rect 276112 550656 276164 550662
rect 276072 550624 276074 550633
rect 276112 550598 276164 550604
rect 276478 550624 276534 550633
rect 276018 550559 276074 550568
rect 276478 550559 276534 550568
rect 276492 549250 276520 550559
rect 276400 549222 276520 549250
rect 276400 539646 276428 549222
rect 276296 539640 276348 539646
rect 276296 539582 276348 539588
rect 276388 539640 276440 539646
rect 276388 539582 276440 539588
rect 276308 531350 276336 539582
rect 276296 531344 276348 531350
rect 276296 531286 276348 531292
rect 276572 531344 276624 531350
rect 276572 531286 276624 531292
rect 276584 526386 276612 531286
rect 276388 526380 276440 526386
rect 276388 526322 276440 526328
rect 276572 526380 276624 526386
rect 276572 526322 276624 526328
rect 276400 520146 276428 526322
rect 277412 520146 277440 700062
rect 279436 523938 279464 700062
rect 279424 523932 279476 523938
rect 279424 523874 279476 523880
rect 276400 520118 276612 520146
rect 277412 520118 278268 520146
rect 276584 520010 276612 520118
rect 278240 520010 278268 520118
rect 280172 520010 280200 700946
rect 283012 700868 283064 700874
rect 283012 700810 283064 700816
rect 281540 700188 281592 700194
rect 281540 700130 281592 700136
rect 281552 520010 281580 700130
rect 283024 520010 283052 700810
rect 283852 699718 283880 703600
rect 287244 700800 287296 700806
rect 287244 700742 287296 700748
rect 284300 700664 284352 700670
rect 284300 700606 284352 700612
rect 283840 699712 283892 699718
rect 283840 699654 283892 699660
rect 284312 520146 284340 700606
rect 287256 695502 287284 700742
rect 288440 700528 288492 700534
rect 288440 700470 288492 700476
rect 287244 695496 287296 695502
rect 287244 695438 287296 695444
rect 287152 688356 287204 688362
rect 287152 688298 287204 688304
rect 287164 678994 287192 688298
rect 287164 678966 287284 678994
rect 287256 676190 287284 678966
rect 287244 676184 287296 676190
rect 287244 676126 287296 676132
rect 287152 666596 287204 666602
rect 287152 666538 287204 666544
rect 287164 659682 287192 666538
rect 287164 659654 287284 659682
rect 287256 649942 287284 659654
rect 287244 649936 287296 649942
rect 287244 649878 287296 649884
rect 287244 649800 287296 649806
rect 287244 649742 287296 649748
rect 287256 630698 287284 649742
rect 287060 630692 287112 630698
rect 287060 630634 287112 630640
rect 287244 630692 287296 630698
rect 287244 630634 287296 630640
rect 287072 630578 287100 630634
rect 287072 630550 287192 630578
rect 287164 621058 287192 630550
rect 287164 621030 287284 621058
rect 287256 611386 287284 621030
rect 287060 611380 287112 611386
rect 287060 611322 287112 611328
rect 287244 611380 287296 611386
rect 287244 611322 287296 611328
rect 287072 611266 287100 611322
rect 287072 611238 287192 611266
rect 287164 608598 287192 611238
rect 287152 608592 287204 608598
rect 287152 608534 287204 608540
rect 287244 599004 287296 599010
rect 287244 598946 287296 598952
rect 287256 572762 287284 598946
rect 287060 572756 287112 572762
rect 287060 572698 287112 572704
rect 287244 572756 287296 572762
rect 287244 572698 287296 572704
rect 287072 572642 287100 572698
rect 287072 572614 287192 572642
rect 287164 563122 287192 572614
rect 287164 563094 287284 563122
rect 287256 560266 287284 563094
rect 287164 560238 287284 560266
rect 287164 550662 287192 560238
rect 287060 550656 287112 550662
rect 287058 550624 287060 550633
rect 287152 550656 287204 550662
rect 287112 550624 287114 550633
rect 287152 550598 287204 550604
rect 287242 550624 287298 550633
rect 287058 550559 287114 550568
rect 287242 550559 287298 550568
rect 287256 549273 287284 550559
rect 287058 549264 287114 549273
rect 287058 549199 287114 549208
rect 287242 549264 287298 549273
rect 287242 549199 287298 549208
rect 287072 540938 287100 549199
rect 287060 540932 287112 540938
rect 287060 540874 287112 540880
rect 287244 540932 287296 540938
rect 287244 540874 287296 540880
rect 287256 539594 287284 540874
rect 287256 539566 287376 539594
rect 287348 534138 287376 539566
rect 287336 534132 287388 534138
rect 287336 534074 287388 534080
rect 287152 531344 287204 531350
rect 287152 531286 287204 531292
rect 287164 524498 287192 531286
rect 287072 524470 287192 524498
rect 287072 524362 287100 524470
rect 287072 524334 287192 524362
rect 284312 520118 284984 520146
rect 284956 520010 284984 520118
rect 273272 519982 273378 520010
rect 274652 519982 275126 520010
rect 276584 519982 276874 520010
rect 278240 519982 278530 520010
rect 280172 519982 280278 520010
rect 281552 519982 281934 520010
rect 283024 519982 283682 520010
rect 284956 519982 285338 520010
rect 287164 519874 287192 524334
rect 288452 520010 288480 700470
rect 290004 700324 290056 700330
rect 290004 700266 290056 700272
rect 290016 695502 290044 700266
rect 291384 698216 291436 698222
rect 291384 698158 291436 698164
rect 291396 695502 291424 698158
rect 290004 695496 290056 695502
rect 290004 695438 290056 695444
rect 291384 695496 291436 695502
rect 291384 695438 291436 695444
rect 300136 688634 300164 703600
rect 332520 699922 332548 703600
rect 336004 700324 336056 700330
rect 336004 700266 336056 700272
rect 332508 699916 332560 699922
rect 332508 699858 332560 699864
rect 289912 688628 289964 688634
rect 289912 688570 289964 688576
rect 291384 688628 291436 688634
rect 291384 688570 291436 688576
rect 299664 688628 299716 688634
rect 299664 688570 299716 688576
rect 300124 688628 300176 688634
rect 300124 688570 300176 688576
rect 289924 678994 289952 688570
rect 291396 685930 291424 688570
rect 299676 685930 299704 688570
rect 291396 685902 291516 685930
rect 291488 679046 291516 685902
rect 299584 685902 299704 685930
rect 299584 684486 299612 685902
rect 299572 684480 299624 684486
rect 299572 684422 299624 684428
rect 292580 681760 292632 681766
rect 292580 681702 292632 681708
rect 291476 679040 291528 679046
rect 289924 678966 290044 678994
rect 291476 678982 291528 678988
rect 290016 669338 290044 678966
rect 291384 678972 291436 678978
rect 291384 678914 291436 678920
rect 289832 669310 290044 669338
rect 289832 666534 289860 669310
rect 289820 666528 289872 666534
rect 289820 666470 289872 666476
rect 289820 656940 289872 656946
rect 289820 656882 289872 656888
rect 289832 647222 289860 656882
rect 289820 647216 289872 647222
rect 289820 647158 289872 647164
rect 289820 637628 289872 637634
rect 289820 637570 289872 637576
rect 289832 630578 289860 637570
rect 291396 637566 291424 678914
rect 291384 637560 291436 637566
rect 291384 637502 291436 637508
rect 289832 630550 289952 630578
rect 289924 627910 289952 630550
rect 291292 627972 291344 627978
rect 291292 627914 291344 627920
rect 289912 627904 289964 627910
rect 289912 627846 289964 627852
rect 291304 627858 291332 627914
rect 291304 627830 291424 627858
rect 290004 618316 290056 618322
rect 290004 618258 290056 618264
rect 290016 611386 290044 618258
rect 291396 618254 291424 627830
rect 291384 618248 291436 618254
rect 291384 618190 291436 618196
rect 289820 611380 289872 611386
rect 289820 611322 289872 611328
rect 290004 611380 290056 611386
rect 290004 611322 290056 611328
rect 289832 591954 289860 611322
rect 291292 608660 291344 608666
rect 291292 608602 291344 608608
rect 291304 607170 291332 608602
rect 291292 607164 291344 607170
rect 291292 607106 291344 607112
rect 291384 597576 291436 597582
rect 291384 597518 291436 597524
rect 289832 591926 290044 591954
rect 290016 572762 290044 591926
rect 291396 579630 291424 597518
rect 291384 579624 291436 579630
rect 291384 579566 291436 579572
rect 289820 572756 289872 572762
rect 289820 572698 289872 572704
rect 290004 572756 290056 572762
rect 290004 572698 290056 572704
rect 289832 572642 289860 572698
rect 289832 572614 289952 572642
rect 289924 563122 289952 572614
rect 291476 569968 291528 569974
rect 291476 569910 291528 569916
rect 291488 563174 291516 569910
rect 291476 563168 291528 563174
rect 289924 563094 290044 563122
rect 291476 563110 291528 563116
rect 290016 553450 290044 563094
rect 291384 563032 291436 563038
rect 291384 562974 291436 562980
rect 291396 560266 291424 562974
rect 291304 560238 291424 560266
rect 289820 553444 289872 553450
rect 289820 553386 289872 553392
rect 290004 553444 290056 553450
rect 290004 553386 290056 553392
rect 289832 543674 289860 553386
rect 291304 553382 291332 560238
rect 291292 553376 291344 553382
rect 291292 553318 291344 553324
rect 291292 553240 291344 553246
rect 291292 553182 291344 553188
rect 291304 549273 291332 553182
rect 291106 549264 291162 549273
rect 291106 549199 291162 549208
rect 291290 549264 291346 549273
rect 291290 549199 291346 549208
rect 289832 543646 289952 543674
rect 289924 534154 289952 543646
rect 291120 540682 291148 549199
rect 292592 548078 292620 681702
rect 296720 667956 296772 667962
rect 296720 667898 296772 667904
rect 295340 652792 295392 652798
rect 295340 652734 295392 652740
rect 292580 548072 292632 548078
rect 292580 548014 292632 548020
rect 293316 548072 293368 548078
rect 293316 548014 293368 548020
rect 291120 540654 291332 540682
rect 289924 534126 290044 534154
rect 290016 520010 290044 534126
rect 291304 531350 291332 540654
rect 293328 531350 293356 548014
rect 291292 531344 291344 531350
rect 291292 531286 291344 531292
rect 291844 531344 291896 531350
rect 293316 531344 293368 531350
rect 291844 531286 291896 531292
rect 293314 531312 293316 531321
rect 293500 531344 293552 531350
rect 293368 531312 293370 531321
rect 291856 526402 291884 531286
rect 293314 531247 293370 531256
rect 293498 531312 293500 531321
rect 293552 531312 293554 531321
rect 293498 531247 293554 531256
rect 291672 526374 291884 526402
rect 291672 520010 291700 526374
rect 293328 520010 293356 531247
rect 295352 520010 295380 652734
rect 296732 520282 296760 667898
rect 299940 666596 299992 666602
rect 299940 666538 299992 666544
rect 299952 659682 299980 666538
rect 299768 659654 299980 659682
rect 299768 647290 299796 659654
rect 299664 647284 299716 647290
rect 299664 647226 299716 647232
rect 299756 647284 299808 647290
rect 299756 647226 299808 647232
rect 299676 640422 299704 647226
rect 299664 640416 299716 640422
rect 299664 640358 299716 640364
rect 299756 640416 299808 640422
rect 299756 640358 299808 640364
rect 299768 630698 299796 640358
rect 299572 630692 299624 630698
rect 299572 630634 299624 630640
rect 299756 630692 299808 630698
rect 299756 630634 299808 630640
rect 299584 630578 299612 630634
rect 299584 630550 299704 630578
rect 298100 623824 298152 623830
rect 298100 623766 298152 623772
rect 296732 520254 296944 520282
rect 296916 520010 296944 520254
rect 298112 520146 298140 623766
rect 299676 621058 299704 630550
rect 299676 621030 299796 621058
rect 299768 611386 299796 621030
rect 336016 617574 336044 700266
rect 348804 700058 348832 703600
rect 364996 700126 365024 703600
rect 397472 700262 397500 703600
rect 413664 700942 413692 703600
rect 413652 700936 413704 700942
rect 413652 700878 413704 700884
rect 429856 700330 429884 703600
rect 462332 700738 462360 703600
rect 462320 700732 462372 700738
rect 462320 700674 462372 700680
rect 478524 700602 478552 703600
rect 494808 703582 494928 703600
rect 478512 700596 478564 700602
rect 478512 700538 478564 700544
rect 429844 700324 429896 700330
rect 429844 700266 429896 700272
rect 397460 700256 397512 700262
rect 397460 700198 397512 700204
rect 364984 700120 365036 700126
rect 364984 700062 365036 700068
rect 348792 700052 348844 700058
rect 348792 699994 348844 700000
rect 494900 686089 494928 703582
rect 527192 700398 527220 703600
rect 527180 700392 527232 700398
rect 543476 700369 543504 703600
rect 527180 700334 527232 700340
rect 543462 700360 543518 700369
rect 543462 700295 543518 700304
rect 559668 688634 559696 703600
rect 579894 698048 579950 698057
rect 579894 697983 579950 697992
rect 579908 696998 579936 697983
rect 579896 696992 579948 696998
rect 579896 696934 579948 696940
rect 559104 688628 559156 688634
rect 559104 688570 559156 688576
rect 559656 688628 559708 688634
rect 559656 688570 559708 688576
rect 494886 686080 494942 686089
rect 494886 686015 494942 686024
rect 494242 685944 494298 685953
rect 559116 685930 559144 688570
rect 580078 686352 580134 686361
rect 580078 686287 580134 686296
rect 494242 685879 494298 685888
rect 559024 685902 559144 685930
rect 580092 685914 580120 686287
rect 580080 685908 580132 685914
rect 494256 678994 494284 685879
rect 559024 684486 559052 685902
rect 580080 685850 580132 685856
rect 559012 684480 559064 684486
rect 559012 684422 559064 684428
rect 494072 678966 494284 678994
rect 494072 676190 494100 678966
rect 494060 676184 494112 676190
rect 494060 676126 494112 676132
rect 580262 674656 580318 674665
rect 580262 674591 580318 674600
rect 580276 673538 580304 674591
rect 580264 673532 580316 673538
rect 580264 673474 580316 673480
rect 494152 666596 494204 666602
rect 494152 666538 494204 666544
rect 559380 666596 559432 666602
rect 559380 666538 559432 666544
rect 494164 659682 494192 666538
rect 559392 659682 559420 666538
rect 494164 659654 494284 659682
rect 494256 654158 494284 659654
rect 559208 659654 559420 659682
rect 494060 654152 494112 654158
rect 494060 654094 494112 654100
rect 494244 654152 494296 654158
rect 494244 654094 494296 654100
rect 494072 644450 494100 654094
rect 559208 647290 559236 659654
rect 579894 651128 579950 651137
rect 579894 651063 579950 651072
rect 579908 650078 579936 651063
rect 579896 650072 579948 650078
rect 579896 650014 579948 650020
rect 559104 647284 559156 647290
rect 559104 647226 559156 647232
rect 559196 647284 559248 647290
rect 559196 647226 559248 647232
rect 494072 644422 494284 644450
rect 494256 634846 494284 644422
rect 559116 640422 559144 647226
rect 559104 640416 559156 640422
rect 559104 640358 559156 640364
rect 559196 640416 559248 640422
rect 559196 640358 559248 640364
rect 494060 634840 494112 634846
rect 494060 634782 494112 634788
rect 494244 634840 494296 634846
rect 494244 634782 494296 634788
rect 494072 625138 494100 634782
rect 559208 630698 559236 640358
rect 580078 639432 580134 639441
rect 580078 639367 580134 639376
rect 580092 638994 580120 639367
rect 580080 638988 580132 638994
rect 580080 638930 580132 638936
rect 559012 630692 559064 630698
rect 559012 630634 559064 630640
rect 559196 630692 559248 630698
rect 559196 630634 559248 630640
rect 559024 630578 559052 630634
rect 559024 630550 559144 630578
rect 494072 625110 494284 625138
rect 336004 617568 336056 617574
rect 336004 617510 336056 617516
rect 494256 615534 494284 625110
rect 559116 621058 559144 630550
rect 580262 627736 580318 627745
rect 580262 627671 580318 627680
rect 580276 626618 580304 627671
rect 580264 626612 580316 626618
rect 580264 626554 580316 626560
rect 559116 621030 559236 621058
rect 494060 615528 494112 615534
rect 494060 615470 494112 615476
rect 494244 615528 494296 615534
rect 494244 615470 494296 615476
rect 299572 611380 299624 611386
rect 299572 611322 299624 611328
rect 299756 611380 299808 611386
rect 299756 611322 299808 611328
rect 299584 611266 299612 611322
rect 299584 611238 299704 611266
rect 299676 608598 299704 611238
rect 302240 610020 302292 610026
rect 302240 609962 302292 609968
rect 299664 608592 299716 608598
rect 299664 608534 299716 608540
rect 299848 601724 299900 601730
rect 299848 601666 299900 601672
rect 299860 598942 299888 601666
rect 299848 598936 299900 598942
rect 299848 598878 299900 598884
rect 299572 594856 299624 594862
rect 299572 594798 299624 594804
rect 299480 572756 299532 572762
rect 299480 572698 299532 572704
rect 299492 553382 299520 572698
rect 299480 553376 299532 553382
rect 299480 553318 299532 553324
rect 299584 520282 299612 594798
rect 299756 589348 299808 589354
rect 299756 589290 299808 589296
rect 299768 582418 299796 589290
rect 299756 582412 299808 582418
rect 299756 582354 299808 582360
rect 299848 582276 299900 582282
rect 299848 582218 299900 582224
rect 299860 572762 299888 582218
rect 299848 572756 299900 572762
rect 299848 572698 299900 572704
rect 299940 553376 299992 553382
rect 299940 553318 299992 553324
rect 299952 543862 299980 553318
rect 299940 543856 299992 543862
rect 299940 543798 299992 543804
rect 299848 543720 299900 543726
rect 299848 543662 299900 543668
rect 299860 540977 299888 543662
rect 299662 540968 299718 540977
rect 299662 540903 299718 540912
rect 299846 540968 299902 540977
rect 299846 540903 299902 540912
rect 299676 531350 299704 540903
rect 299664 531344 299716 531350
rect 299664 531286 299716 531292
rect 299940 531344 299992 531350
rect 299940 531286 299992 531292
rect 299952 523870 299980 531286
rect 299940 523864 299992 523870
rect 299940 523806 299992 523812
rect 299584 520254 300440 520282
rect 298112 520118 298600 520146
rect 298572 520010 298600 520118
rect 300412 520010 300440 520254
rect 302252 520010 302280 609962
rect 494072 605826 494100 615470
rect 559208 611386 559236 621030
rect 559012 611380 559064 611386
rect 559012 611322 559064 611328
rect 559196 611380 559248 611386
rect 559196 611322 559248 611328
rect 559024 611266 559052 611322
rect 559024 611238 559144 611266
rect 559116 608598 559144 611238
rect 559104 608592 559156 608598
rect 559104 608534 559156 608540
rect 494072 605798 494284 605826
rect 494256 596222 494284 605798
rect 579894 604208 579950 604217
rect 579894 604143 579950 604152
rect 579908 603158 579936 604143
rect 579896 603152 579948 603158
rect 579896 603094 579948 603100
rect 559288 601724 559340 601730
rect 559288 601666 559340 601672
rect 559300 598942 559328 601666
rect 559288 598936 559340 598942
rect 559288 598878 559340 598884
rect 494060 596216 494112 596222
rect 494244 596216 494296 596222
rect 494112 596164 494192 596170
rect 494060 596158 494192 596164
rect 494244 596158 494296 596164
rect 494072 596142 494192 596158
rect 494164 596034 494192 596142
rect 494164 596006 494284 596034
rect 494256 591954 494284 596006
rect 580078 592512 580134 592521
rect 580078 592447 580134 592456
rect 580092 592074 580120 592447
rect 580080 592068 580132 592074
rect 580080 592010 580132 592016
rect 494164 591926 494284 591954
rect 494164 589286 494192 591926
rect 559380 589348 559432 589354
rect 559380 589290 559432 589296
rect 493876 589280 493928 589286
rect 493876 589222 493928 589228
rect 494152 589280 494204 589286
rect 494152 589222 494204 589228
rect 493888 579737 493916 589222
rect 559392 582486 559420 589290
rect 559380 582480 559432 582486
rect 559380 582422 559432 582428
rect 559288 582344 559340 582350
rect 559288 582286 559340 582292
rect 493874 579728 493930 579737
rect 493874 579663 493930 579672
rect 494058 579728 494114 579737
rect 494058 579663 494114 579672
rect 494072 572642 494100 579663
rect 559300 572642 559328 582286
rect 580262 580816 580318 580825
rect 580262 580751 580318 580760
rect 580276 579698 580304 580751
rect 580264 579692 580316 579698
rect 580264 579634 580316 579640
rect 494072 572614 494192 572642
rect 494164 569906 494192 572614
rect 559116 572614 559328 572642
rect 559116 569922 559144 572614
rect 494152 569900 494204 569906
rect 494152 569842 494204 569848
rect 559024 569894 559144 569922
rect 303620 567248 303672 567254
rect 303620 567190 303672 567196
rect 303632 520010 303660 567190
rect 559024 563174 559052 569894
rect 559012 563168 559064 563174
rect 559012 563110 559064 563116
rect 494336 563100 494388 563106
rect 494336 563042 494388 563048
rect 494348 560289 494376 563042
rect 559012 563032 559064 563038
rect 559012 562974 559064 562980
rect 494150 560280 494206 560289
rect 494150 560215 494206 560224
rect 494334 560280 494390 560289
rect 559024 560250 559052 562974
rect 494334 560215 494390 560224
rect 559012 560244 559064 560250
rect 306380 552084 306432 552090
rect 306380 552026 306432 552032
rect 305000 538280 305052 538286
rect 305000 538222 305052 538228
rect 305012 520146 305040 538222
rect 306392 520146 306420 552026
rect 494164 550662 494192 560215
rect 559012 560186 559064 560192
rect 579894 557288 579950 557297
rect 579894 557223 579950 557232
rect 579908 556238 579936 557223
rect 579896 556232 579948 556238
rect 579896 556174 579948 556180
rect 494152 550656 494204 550662
rect 494152 550598 494204 550604
rect 494428 550656 494480 550662
rect 494428 550598 494480 550604
rect 559196 550656 559248 550662
rect 559196 550598 559248 550604
rect 494440 543862 494468 550598
rect 494428 543856 494480 543862
rect 494428 543798 494480 543804
rect 494336 543720 494388 543726
rect 494336 543662 494388 543668
rect 494348 540977 494376 543662
rect 559208 543658 559236 550598
rect 580078 545592 580134 545601
rect 580078 545527 580134 545536
rect 580092 545154 580120 545527
rect 580080 545148 580132 545154
rect 580080 545090 580132 545096
rect 559012 543652 559064 543658
rect 559012 543594 559064 543600
rect 559196 543652 559248 543658
rect 559196 543594 559248 543600
rect 494150 540968 494206 540977
rect 494150 540903 494206 540912
rect 494334 540968 494390 540977
rect 494334 540903 494390 540912
rect 494164 531350 494192 540903
rect 559024 534018 559052 543594
rect 559024 533990 559144 534018
rect 494152 531344 494204 531350
rect 494152 531286 494204 531292
rect 494428 531344 494480 531350
rect 494428 531286 494480 531292
rect 494440 523802 494468 531286
rect 559116 524498 559144 533990
rect 580262 533896 580318 533905
rect 580262 533831 580318 533840
rect 580276 532778 580304 533831
rect 580264 532772 580316 532778
rect 580264 532714 580316 532720
rect 559116 524470 559236 524498
rect 494428 523796 494480 523802
rect 494428 523738 494480 523744
rect 559208 523734 559236 524470
rect 559196 523728 559248 523734
rect 559196 523670 559248 523676
rect 371056 522980 371108 522986
rect 371056 522922 371108 522928
rect 370780 522912 370832 522918
rect 370780 522854 370832 522860
rect 309140 522776 309192 522782
rect 309140 522718 309192 522724
rect 305012 520118 305224 520146
rect 306392 520118 307064 520146
rect 305196 520010 305224 520118
rect 307036 520010 307064 520118
rect 309152 520010 309180 522718
rect 312452 522708 312504 522714
rect 312452 522650 312504 522656
rect 310612 522640 310664 522646
rect 310612 522582 310664 522588
rect 310624 520010 310652 522582
rect 311806 522200 311862 522209
rect 311806 522135 311862 522144
rect 311990 522200 312046 522209
rect 311990 522135 312046 522144
rect 311820 521626 311848 522135
rect 312004 521626 312032 522135
rect 311808 521620 311860 521626
rect 311808 521562 311860 521568
rect 311992 521620 312044 521626
rect 311992 521562 312044 521568
rect 312464 520010 312492 522650
rect 370502 522608 370558 522617
rect 317420 522572 317472 522578
rect 370502 522543 370558 522552
rect 317420 522514 317472 522520
rect 317432 520010 317460 522514
rect 319260 522504 319312 522510
rect 319260 522446 319312 522452
rect 353482 522472 353538 522481
rect 319272 520010 319300 522446
rect 323032 522436 323084 522442
rect 323032 522378 323084 522384
rect 325700 522436 325752 522442
rect 325700 522378 325752 522384
rect 335268 522436 335320 522442
rect 353482 522407 353538 522416
rect 335268 522378 335320 522384
rect 288452 519982 288834 520010
rect 290016 519982 290490 520010
rect 291672 519982 292238 520010
rect 293328 519982 293894 520010
rect 295352 519982 295642 520010
rect 296916 519982 297390 520010
rect 298572 519982 299046 520010
rect 300412 519982 300794 520010
rect 302252 519982 302450 520010
rect 303632 519982 304198 520010
rect 305196 519982 305854 520010
rect 307036 519982 307602 520010
rect 309152 519982 309350 520010
rect 310624 519982 311006 520010
rect 312464 519982 312754 520010
rect 317432 519982 317814 520010
rect 319272 519982 319562 520010
rect 323044 519874 323072 522378
rect 325712 522209 325740 522378
rect 327724 522368 327776 522374
rect 327724 522310 327776 522316
rect 326068 522300 326120 522306
rect 326068 522242 326120 522248
rect 325698 522200 325754 522209
rect 325698 522135 325754 522144
rect 326080 520010 326108 522242
rect 327736 520010 327764 522310
rect 335280 522209 335308 522378
rect 343180 522232 343232 522238
rect 335266 522200 335322 522209
rect 332876 522164 332928 522170
rect 345020 522232 345072 522238
rect 343180 522174 343232 522180
rect 345018 522200 345020 522209
rect 345072 522200 345074 522209
rect 335266 522135 335322 522144
rect 332876 522106 332928 522112
rect 331220 522028 331272 522034
rect 331220 521970 331272 521976
rect 331232 520010 331260 521970
rect 332888 520010 332916 522106
rect 338120 522096 338172 522102
rect 338120 522038 338172 522044
rect 334532 521892 334584 521898
rect 334532 521834 334584 521840
rect 334544 520010 334572 521834
rect 336372 521824 336424 521830
rect 336372 521766 336424 521772
rect 336384 520010 336412 521766
rect 338132 520010 338160 522038
rect 343192 520010 343220 522174
rect 345018 522135 345074 522144
rect 348332 521960 348384 521966
rect 348332 521902 348384 521908
rect 346492 521756 346544 521762
rect 346492 521698 346544 521704
rect 346504 520010 346532 521698
rect 348344 520010 348372 521902
rect 353496 520010 353524 522407
rect 356794 522336 356850 522345
rect 356794 522271 356850 522280
rect 354588 522232 354640 522238
rect 354586 522200 354588 522209
rect 354640 522200 354642 522209
rect 354586 522135 354642 522144
rect 356808 520010 356836 522271
rect 369768 520872 369820 520878
rect 369768 520814 369820 520820
rect 369676 520600 369728 520606
rect 369676 520542 369728 520548
rect 369584 520532 369636 520538
rect 369584 520474 369636 520480
rect 369492 520464 369544 520470
rect 369492 520406 369544 520412
rect 326080 519982 326370 520010
rect 327736 519982 328118 520010
rect 331232 519982 331522 520010
rect 332888 519982 333270 520010
rect 334544 519982 334926 520010
rect 336384 519982 336674 520010
rect 338132 519982 338330 520010
rect 343192 519982 343482 520010
rect 346504 519982 346886 520010
rect 348344 519982 348634 520010
rect 353496 519982 353786 520010
rect 356808 519982 357190 520010
rect 231872 519846 232346 519874
rect 233252 519846 234094 519874
rect 239246 519846 239628 519874
rect 240902 519846 241284 519874
rect 242650 519846 242848 519874
rect 244306 519846 244688 519874
rect 246054 519846 246344 519874
rect 247802 519846 248184 519874
rect 249458 519846 249748 519874
rect 251206 519846 251496 519874
rect 252862 519846 253152 519874
rect 254610 519846 254992 519874
rect 256358 519846 256648 519874
rect 258014 519846 258120 519874
rect 259762 519846 260144 519874
rect 261418 519846 261800 519874
rect 263166 519846 263364 519874
rect 264822 519846 264928 519874
rect 266570 519846 267044 519874
rect 268318 519846 268608 519874
rect 271722 519846 271828 519874
rect 287086 519846 287192 519874
rect 322966 519846 323072 519874
rect 179354 519586 179460 519602
rect 215326 519586 215616 519602
rect 179354 519580 179472 519586
rect 179354 519574 179420 519580
rect 215326 519580 215628 519586
rect 215326 519574 215576 519580
rect 179420 519522 179472 519528
rect 215576 519522 215628 519528
rect 314108 519512 314160 519518
rect 314160 519460 314410 519466
rect 314108 519454 314410 519460
rect 314120 519438 314410 519454
rect 320928 519450 321310 519466
rect 320916 519444 321310 519450
rect 320968 519438 321310 519444
rect 320916 519386 320968 519392
rect 324412 519376 324464 519382
rect 172886 519344 172942 519353
rect 169772 519302 170890 519330
rect 172546 519302 172886 519330
rect 37186 517984 37242 517993
rect 37186 517919 37242 517928
rect 57886 517984 57942 517993
rect 57886 517919 57942 517928
rect 77206 517984 77262 517993
rect 77206 517919 77262 517928
rect 96526 517984 96582 517993
rect 96526 517919 96582 517928
rect 115846 517984 115902 517993
rect 115846 517919 115902 517928
rect 135166 517984 135222 517993
rect 135166 517919 135222 517928
rect 154486 517984 154542 517993
rect 154486 517919 154542 517928
rect 166998 517984 167054 517993
rect 166998 517919 167054 517928
rect 37200 517614 37228 517919
rect 57900 517886 57928 517919
rect 77220 517886 77248 517919
rect 96540 517886 96568 517919
rect 115860 517886 115888 517919
rect 135180 517886 135208 517919
rect 154500 517886 154528 517919
rect 50988 517880 51040 517886
rect 50986 517848 50988 517857
rect 57888 517880 57940 517886
rect 51040 517848 51042 517857
rect 70308 517880 70360 517886
rect 57888 517822 57940 517828
rect 70306 517848 70308 517857
rect 77208 517880 77260 517886
rect 70360 517848 70362 517857
rect 50986 517783 51042 517792
rect 89628 517880 89680 517886
rect 77208 517822 77260 517828
rect 89626 517848 89628 517857
rect 96528 517880 96580 517886
rect 89680 517848 89682 517857
rect 70306 517783 70362 517792
rect 108948 517880 109000 517886
rect 96528 517822 96580 517828
rect 108946 517848 108948 517857
rect 115848 517880 115900 517886
rect 109000 517848 109002 517857
rect 89626 517783 89682 517792
rect 128268 517880 128320 517886
rect 115848 517822 115900 517828
rect 128266 517848 128268 517857
rect 135168 517880 135220 517886
rect 128320 517848 128322 517857
rect 108946 517783 109002 517792
rect 147588 517880 147640 517886
rect 135168 517822 135220 517828
rect 147586 517848 147588 517857
rect 154488 517880 154540 517886
rect 147640 517848 147642 517857
rect 128266 517783 128322 517792
rect 154488 517822 154540 517828
rect 166906 517848 166962 517857
rect 147586 517783 147642 517792
rect 167012 517834 167040 517919
rect 166962 517806 167040 517834
rect 166906 517783 166962 517792
rect 37188 517608 37240 517614
rect 37188 517550 37240 517556
rect 88984 218000 89036 218006
rect 88984 217942 89036 217948
rect 86224 217932 86276 217938
rect 86224 217874 86276 217880
rect 77944 217864 77996 217870
rect 77944 217806 77996 217812
rect 75184 217796 75236 217802
rect 75184 217738 75236 217744
rect 71044 217728 71096 217734
rect 71044 217670 71096 217676
rect 42064 217660 42116 217666
rect 42064 217602 42116 217608
rect 35164 217592 35216 217598
rect 35164 217534 35216 217540
rect 32404 217524 32456 217530
rect 32404 217466 32456 217472
rect 31024 217456 31076 217462
rect 31024 217398 31076 217404
rect 28264 108996 28316 109002
rect 28264 108938 28316 108944
rect 28908 10328 28960 10334
rect 28908 10270 28960 10276
rect 26700 6316 26752 6322
rect 26700 6258 26752 6264
rect 24308 3868 24360 3874
rect 24308 3810 24360 3816
rect 24124 3732 24176 3738
rect 24124 3674 24176 3680
rect 24320 400 24348 3810
rect 25504 3800 25556 3806
rect 25504 3742 25556 3748
rect 25516 400 25544 3742
rect 26712 400 26740 6258
rect 28920 3398 28948 10270
rect 30288 6384 30340 6390
rect 30288 6326 30340 6332
rect 29092 3732 29144 3738
rect 29092 3674 29144 3680
rect 27896 3392 27948 3398
rect 27896 3334 27948 3340
rect 28908 3392 28960 3398
rect 28908 3334 28960 3340
rect 27908 400 27936 3334
rect 29104 400 29132 3674
rect 30300 400 30328 6326
rect 31036 3874 31064 217398
rect 31668 11756 31720 11762
rect 31668 11698 31720 11704
rect 31024 3868 31076 3874
rect 31024 3810 31076 3816
rect 31680 3346 31708 11698
rect 32416 3806 32444 217466
rect 33876 6452 33928 6458
rect 33876 6394 33928 6400
rect 32404 3800 32456 3806
rect 32404 3742 32456 3748
rect 31496 3318 31708 3346
rect 32680 3392 32732 3398
rect 32680 3334 32732 3340
rect 31496 400 31524 3318
rect 32692 400 32720 3334
rect 33888 400 33916 6394
rect 34980 3800 35032 3806
rect 34980 3742 35032 3748
rect 34992 400 35020 3742
rect 35176 3398 35204 217534
rect 40960 6588 41012 6594
rect 40960 6530 41012 6536
rect 37372 6520 37424 6526
rect 37372 6462 37424 6468
rect 36176 3868 36228 3874
rect 36176 3810 36228 3816
rect 35164 3392 35216 3398
rect 35164 3334 35216 3340
rect 36188 400 36216 3810
rect 37384 400 37412 6462
rect 39764 3392 39816 3398
rect 39764 3334 39816 3340
rect 38568 3324 38620 3330
rect 38568 3266 38620 3272
rect 38580 400 38608 3266
rect 39776 400 39804 3334
rect 40972 400 41000 6530
rect 42076 3398 42104 217602
rect 67180 9172 67232 9178
rect 67180 9114 67232 9120
rect 63592 7744 63644 7750
rect 63592 7686 63644 7692
rect 60004 7676 60056 7682
rect 60004 7618 60056 7624
rect 56416 7608 56468 7614
rect 52826 7576 52882 7585
rect 56416 7550 56468 7556
rect 52826 7511 52882 7520
rect 49332 6724 49384 6730
rect 49332 6666 49384 6672
rect 44548 6656 44600 6662
rect 44548 6598 44600 6604
rect 43352 4004 43404 4010
rect 43352 3946 43404 3952
rect 42156 3936 42208 3942
rect 42156 3878 42208 3884
rect 42064 3392 42116 3398
rect 42064 3334 42116 3340
rect 42168 400 42196 3878
rect 43364 400 43392 3946
rect 44560 400 44588 6598
rect 48136 5160 48188 5166
rect 48136 5102 48188 5108
rect 45744 3256 45796 3262
rect 45744 3198 45796 3204
rect 45756 400 45784 3198
rect 46940 2984 46992 2990
rect 46940 2926 46992 2932
rect 46952 400 46980 2926
rect 48148 400 48176 5102
rect 49344 400 49372 6666
rect 51632 5228 51684 5234
rect 51632 5170 51684 5176
rect 50528 3120 50580 3126
rect 50528 3062 50580 3068
rect 50540 400 50568 3062
rect 51644 400 51672 5170
rect 52840 400 52868 7511
rect 55220 5296 55272 5302
rect 55220 5238 55272 5244
rect 54024 4072 54076 4078
rect 54024 4014 54076 4020
rect 54036 400 54064 4014
rect 55232 400 55260 5238
rect 56428 400 56456 7550
rect 58808 5364 58860 5370
rect 58808 5306 58860 5312
rect 57612 3188 57664 3194
rect 57612 3130 57664 3136
rect 57624 400 57652 3130
rect 58820 400 58848 5306
rect 60016 400 60044 7618
rect 62396 5432 62448 5438
rect 62396 5374 62448 5380
rect 61200 4140 61252 4146
rect 61200 4082 61252 4088
rect 61212 400 61240 4082
rect 62408 400 62436 5374
rect 63604 400 63632 7686
rect 65984 5500 66036 5506
rect 65984 5442 66036 5448
rect 64788 2916 64840 2922
rect 64788 2858 64840 2864
rect 64800 400 64828 2858
rect 65996 400 66024 5442
rect 67192 400 67220 9114
rect 69480 4752 69532 4758
rect 69480 4694 69532 4700
rect 68284 3324 68336 3330
rect 68284 3266 68336 3272
rect 68296 400 68324 3266
rect 69492 400 69520 4694
rect 70676 3392 70728 3398
rect 70676 3334 70728 3340
rect 70688 400 70716 3334
rect 71056 3262 71084 217670
rect 74448 10464 74500 10470
rect 74448 10406 74500 10412
rect 71688 10396 71740 10402
rect 71688 10338 71740 10344
rect 71700 3398 71728 10338
rect 73068 6792 73120 6798
rect 73068 6734 73120 6740
rect 71688 3392 71740 3398
rect 71688 3334 71740 3340
rect 71044 3256 71096 3262
rect 71044 3198 71096 3204
rect 71872 2984 71924 2990
rect 71872 2926 71924 2932
rect 71884 400 71912 2926
rect 73080 400 73108 6734
rect 74460 3482 74488 10406
rect 74276 3454 74488 3482
rect 74276 400 74304 3454
rect 75196 2854 75224 217738
rect 76656 7812 76708 7818
rect 76656 7754 76708 7760
rect 75184 2848 75236 2854
rect 75184 2790 75236 2796
rect 75460 2848 75512 2854
rect 75460 2790 75512 2796
rect 75472 400 75500 2790
rect 76668 400 76696 7754
rect 77852 3324 77904 3330
rect 77852 3266 77904 3272
rect 77864 400 77892 3266
rect 77956 3126 77984 217806
rect 84844 217252 84896 217258
rect 84844 217194 84896 217200
rect 82728 10600 82780 10606
rect 82728 10542 82780 10548
rect 78588 10532 78640 10538
rect 78588 10474 78640 10480
rect 78600 3330 78628 10474
rect 80244 7880 80296 7886
rect 80244 7822 80296 7828
rect 78588 3324 78640 3330
rect 78588 3266 78640 3272
rect 77944 3120 77996 3126
rect 77944 3062 77996 3068
rect 79048 3120 79100 3126
rect 79048 3062 79100 3068
rect 79060 400 79088 3062
rect 80256 400 80284 7822
rect 82740 3330 82768 10542
rect 83832 7948 83884 7954
rect 83832 7890 83884 7896
rect 81440 3324 81492 3330
rect 81440 3266 81492 3272
rect 82728 3324 82780 3330
rect 82728 3266 82780 3272
rect 81452 400 81480 3266
rect 82636 3188 82688 3194
rect 82636 3130 82688 3136
rect 82648 400 82676 3130
rect 83844 400 83872 7890
rect 84856 2990 84884 217194
rect 85488 10668 85540 10674
rect 85488 10610 85540 10616
rect 85500 3262 85528 10610
rect 84936 3256 84988 3262
rect 84936 3198 84988 3204
rect 85488 3256 85540 3262
rect 85488 3198 85540 3204
rect 84844 2984 84896 2990
rect 84844 2926 84896 2932
rect 84948 400 84976 3198
rect 86132 3120 86184 3126
rect 86132 3062 86184 3068
rect 86144 400 86172 3062
rect 86236 2854 86264 217874
rect 87328 8016 87380 8022
rect 87328 7958 87380 7964
rect 86224 2848 86276 2854
rect 86224 2790 86276 2796
rect 87340 400 87368 7958
rect 88524 3188 88576 3194
rect 88524 3130 88576 3136
rect 88536 400 88564 3130
rect 88996 2990 89024 217942
rect 95884 217184 95936 217190
rect 95884 217126 95936 217132
rect 92388 10804 92440 10810
rect 92388 10746 92440 10752
rect 89628 10736 89680 10742
rect 89628 10678 89680 10684
rect 89640 3194 89668 10678
rect 90916 8084 90968 8090
rect 90916 8026 90968 8032
rect 89628 3188 89680 3194
rect 89628 3130 89680 3136
rect 88984 2984 89036 2990
rect 88984 2926 89036 2932
rect 89720 2984 89772 2990
rect 89720 2926 89772 2932
rect 89732 400 89760 2926
rect 90928 400 90956 8026
rect 92400 3346 92428 10746
rect 94504 8152 94556 8158
rect 94504 8094 94556 8100
rect 92124 3318 92428 3346
rect 92124 400 92152 3318
rect 93308 3120 93360 3126
rect 93308 3062 93360 3068
rect 93320 400 93348 3062
rect 94516 400 94544 8094
rect 95700 3052 95752 3058
rect 95700 2994 95752 3000
rect 95712 400 95740 2994
rect 95896 2990 95924 217126
rect 104808 217116 104860 217122
rect 104808 217058 104860 217064
rect 102784 217048 102836 217054
rect 102784 216990 102836 216996
rect 97264 216776 97316 216782
rect 97264 216718 97316 216724
rect 96528 10872 96580 10878
rect 96528 10814 96580 10820
rect 96540 3058 96568 10814
rect 96528 3052 96580 3058
rect 96528 2994 96580 3000
rect 96896 3052 96948 3058
rect 96896 2994 96948 3000
rect 95884 2984 95936 2990
rect 95884 2926 95936 2932
rect 96908 400 96936 2994
rect 97276 2854 97304 216718
rect 99288 10940 99340 10946
rect 99288 10882 99340 10888
rect 98092 8220 98144 8226
rect 98092 8162 98144 8168
rect 97264 2848 97316 2854
rect 97264 2790 97316 2796
rect 98104 400 98132 8162
rect 99300 400 99328 10882
rect 101588 8288 101640 8294
rect 101588 8230 101640 8236
rect 100484 2984 100536 2990
rect 100484 2926 100536 2932
rect 100496 400 100524 2926
rect 101600 400 101628 8230
rect 102796 3210 102824 216990
rect 103428 11008 103480 11014
rect 103428 10950 103480 10956
rect 102612 3182 102824 3210
rect 102612 3058 102640 3182
rect 103440 3058 103468 10950
rect 104820 3058 104848 217058
rect 111708 216980 111760 216986
rect 111708 216922 111760 216928
rect 106924 216708 106976 216714
rect 106924 216650 106976 216656
rect 105176 7540 105228 7546
rect 105176 7482 105228 7488
rect 102600 3052 102652 3058
rect 102600 2994 102652 3000
rect 102784 3052 102836 3058
rect 102784 2994 102836 3000
rect 103428 3052 103480 3058
rect 103428 2994 103480 3000
rect 103980 3052 104032 3058
rect 103980 2994 104032 3000
rect 104808 3052 104860 3058
rect 104808 2994 104860 3000
rect 102796 400 102824 2994
rect 103992 400 104020 2994
rect 105188 400 105216 7482
rect 106372 3052 106424 3058
rect 106372 2994 106424 3000
rect 106384 400 106412 2994
rect 106936 2922 106964 216650
rect 107568 10260 107620 10266
rect 107568 10202 107620 10208
rect 107580 3058 107608 10202
rect 110328 10192 110380 10198
rect 110328 10134 110380 10140
rect 108764 7472 108816 7478
rect 108764 7414 108816 7420
rect 107568 3052 107620 3058
rect 107568 2994 107620 3000
rect 106924 2916 106976 2922
rect 106924 2858 106976 2864
rect 107568 2848 107620 2854
rect 107568 2790 107620 2796
rect 107580 400 107608 2790
rect 108776 400 108804 7414
rect 110340 3482 110368 10134
rect 109972 3454 110368 3482
rect 109972 400 110000 3454
rect 111720 3058 111748 216922
rect 118608 216912 118660 216918
rect 118608 216854 118660 216860
rect 114468 10124 114520 10130
rect 114468 10066 114520 10072
rect 112352 7404 112404 7410
rect 112352 7346 112404 7352
rect 111156 3052 111208 3058
rect 111156 2994 111208 3000
rect 111708 3052 111760 3058
rect 111708 2994 111760 3000
rect 111168 400 111196 2994
rect 112364 400 112392 7346
rect 114480 2990 114508 10066
rect 117136 8696 117188 8702
rect 117136 8638 117188 8644
rect 115940 7336 115992 7342
rect 115940 7278 115992 7284
rect 113548 2984 113600 2990
rect 113548 2926 113600 2932
rect 114468 2984 114520 2990
rect 114468 2926 114520 2932
rect 113560 400 113588 2926
rect 114744 2916 114796 2922
rect 114744 2858 114796 2864
rect 114756 400 114784 2858
rect 115952 400 115980 7278
rect 117148 400 117176 8638
rect 118620 490 118648 216854
rect 122748 216844 122800 216850
rect 122748 216786 122800 216792
rect 121368 11824 121420 11830
rect 121368 11766 121420 11772
rect 119436 7268 119488 7274
rect 119436 7210 119488 7216
rect 118252 462 118648 490
rect 118252 400 118280 462
rect 119448 400 119476 7210
rect 121380 2990 121408 11766
rect 120632 2984 120684 2990
rect 120632 2926 120684 2932
rect 121368 2984 121420 2990
rect 121368 2926 121420 2932
rect 120644 400 120672 2926
rect 122760 2854 122788 216786
rect 169772 17950 169800 519302
rect 193126 519344 193182 519353
rect 193062 519302 193126 519330
rect 172886 519279 172942 519288
rect 195058 519344 195114 519353
rect 194810 519302 195058 519330
rect 193126 519279 193182 519288
rect 198370 519344 198426 519353
rect 198214 519302 198370 519330
rect 195058 519279 195114 519288
rect 199934 519344 199990 519353
rect 199870 519302 199934 519330
rect 198370 519279 198426 519288
rect 205178 519344 205234 519353
rect 205022 519302 205178 519330
rect 199934 519279 199990 519288
rect 210330 519344 210386 519353
rect 210174 519302 210330 519330
rect 205178 519279 205234 519288
rect 225786 519344 225842 519353
rect 225538 519302 225786 519330
rect 210330 519279 210386 519288
rect 225786 519279 225842 519288
rect 315762 519344 315818 519353
rect 315818 519302 316158 519330
rect 339684 519376 339736 519382
rect 324464 519324 324714 519330
rect 324412 519318 324714 519324
rect 324424 519302 324714 519318
rect 329668 519314 329866 519330
rect 341614 519344 341670 519353
rect 339736 519324 340078 519330
rect 339684 519318 340078 519324
rect 329656 519308 329866 519314
rect 315762 519279 315818 519288
rect 329708 519302 329866 519308
rect 339696 519302 340078 519318
rect 359002 519344 359058 519353
rect 341670 519302 341826 519330
rect 345032 519314 345230 519330
rect 350000 519314 350382 519330
rect 351840 519314 352038 519330
rect 355152 519314 355442 519330
rect 345020 519308 345230 519314
rect 341614 519279 341670 519288
rect 329656 519250 329708 519256
rect 345072 519302 345230 519308
rect 349988 519308 350382 519314
rect 345020 519250 345072 519256
rect 350040 519302 350382 519308
rect 351828 519308 352038 519314
rect 349988 519250 350040 519256
rect 351880 519302 352038 519308
rect 355140 519308 355442 519314
rect 351828 519250 351880 519256
rect 355192 519302 355442 519308
rect 358846 519302 359002 519330
rect 361946 519344 362002 519353
rect 360304 519314 360594 519330
rect 359002 519279 359058 519288
rect 360292 519308 360594 519314
rect 355140 519250 355192 519256
rect 360344 519302 360594 519308
rect 363602 519344 363658 519353
rect 362002 519302 362342 519330
rect 361946 519279 362002 519288
rect 363658 519302 363998 519330
rect 363602 519279 363658 519288
rect 360292 519250 360344 519256
rect 369504 322810 369532 520406
rect 369596 346390 369624 520474
rect 369688 369850 369716 520542
rect 369780 510610 369808 520814
rect 370320 518696 370372 518702
rect 370318 518664 370320 518673
rect 370372 518664 370374 518673
rect 370318 518599 370374 518608
rect 369768 510604 369820 510610
rect 369768 510546 369820 510552
rect 369676 369844 369728 369850
rect 369676 369786 369728 369792
rect 369584 346384 369636 346390
rect 369584 346326 369636 346332
rect 369676 322924 369728 322930
rect 369676 322866 369728 322872
rect 369688 322810 369716 322866
rect 369504 322782 369716 322810
rect 223698 220238 223896 220266
rect 170048 220102 170246 220130
rect 170324 220102 170614 220130
rect 170692 220102 170982 220130
rect 171244 220102 171442 220130
rect 169944 210520 169996 210526
rect 169944 210462 169996 210468
rect 169852 210452 169904 210458
rect 169852 210394 169904 210400
rect 169760 17944 169812 17950
rect 169760 17886 169812 17892
rect 125508 11892 125560 11898
rect 125508 11834 125560 11840
rect 123024 7200 123076 7206
rect 123024 7142 123076 7148
rect 121828 2848 121880 2854
rect 121828 2790 121880 2796
rect 122748 2848 122800 2854
rect 122748 2790 122800 2796
rect 121840 400 121868 2790
rect 123036 400 123064 7142
rect 125520 2854 125548 11834
rect 150348 10056 150400 10062
rect 150348 9998 150400 10004
rect 138480 9648 138532 9654
rect 138480 9590 138532 9596
rect 137284 9580 137336 9586
rect 137284 9522 137336 9528
rect 134892 9512 134944 9518
rect 134892 9454 134944 9460
rect 131396 9444 131448 9450
rect 131396 9386 131448 9392
rect 130200 9308 130252 9314
rect 130200 9250 130252 9256
rect 126612 9240 126664 9246
rect 126612 9182 126664 9188
rect 124220 2848 124272 2854
rect 124220 2790 124272 2796
rect 125508 2848 125560 2854
rect 125508 2790 125560 2796
rect 124232 400 124260 2790
rect 125416 2780 125468 2786
rect 125416 2722 125468 2728
rect 125428 400 125456 2722
rect 126624 400 126652 9182
rect 129004 6860 129056 6866
rect 129004 6802 129056 6808
rect 127808 4684 127860 4690
rect 127808 4626 127860 4632
rect 127820 400 127848 4626
rect 129016 400 129044 6802
rect 130212 400 130240 9250
rect 131408 400 131436 9386
rect 133788 9376 133840 9382
rect 133788 9318 133840 9324
rect 132592 6112 132644 6118
rect 132592 6054 132644 6060
rect 132604 400 132632 6054
rect 133800 400 133828 9318
rect 134904 400 134932 9454
rect 136088 6044 136140 6050
rect 136088 5986 136140 5992
rect 136100 400 136128 5986
rect 137296 400 137324 9522
rect 138492 400 138520 9590
rect 140872 8900 140924 8906
rect 140872 8842 140924 8848
rect 139676 5976 139728 5982
rect 139676 5918 139728 5924
rect 139688 400 139716 5918
rect 140884 400 140912 8842
rect 142068 8832 142120 8838
rect 142068 8774 142120 8780
rect 142080 400 142108 8774
rect 145656 8764 145708 8770
rect 145656 8706 145708 8712
rect 143264 5908 143316 5914
rect 143264 5850 143316 5856
rect 143276 400 143304 5850
rect 144460 4616 144512 4622
rect 144460 4558 144512 4564
rect 144472 400 144500 4558
rect 145668 400 145696 8706
rect 146852 5840 146904 5846
rect 146852 5782 146904 5788
rect 146864 400 146892 5782
rect 148048 4548 148100 4554
rect 148048 4490 148100 4496
rect 148060 400 148088 4490
rect 150360 3346 150388 9998
rect 153108 9988 153160 9994
rect 153108 9930 153160 9936
rect 150440 5772 150492 5778
rect 150440 5714 150492 5720
rect 149256 3318 150388 3346
rect 149256 400 149284 3318
rect 150452 400 150480 5714
rect 151544 4480 151596 4486
rect 151544 4422 151596 4428
rect 151556 400 151584 4422
rect 153120 3482 153148 9930
rect 157248 9920 157300 9926
rect 157248 9862 157300 9868
rect 153936 7132 153988 7138
rect 153936 7074 153988 7080
rect 152752 3454 153148 3482
rect 152752 400 152780 3454
rect 153948 400 153976 7074
rect 155132 4412 155184 4418
rect 155132 4354 155184 4360
rect 155144 400 155172 4354
rect 157260 3482 157288 9862
rect 162308 8628 162360 8634
rect 162308 8570 162360 8576
rect 157524 7064 157576 7070
rect 157524 7006 157576 7012
rect 156340 3454 157288 3482
rect 156340 400 156368 3454
rect 157536 400 157564 7006
rect 161112 6996 161164 7002
rect 161112 6938 161164 6944
rect 159916 5704 159968 5710
rect 159916 5646 159968 5652
rect 158720 4344 158772 4350
rect 158720 4286 158772 4292
rect 158732 400 158760 4286
rect 159928 400 159956 5646
rect 161124 400 161152 6938
rect 162320 400 162348 8570
rect 165896 8560 165948 8566
rect 165896 8502 165948 8508
rect 164700 5636 164752 5642
rect 164700 5578 164752 5584
rect 163504 4276 163556 4282
rect 163504 4218 163556 4224
rect 163516 400 163544 4218
rect 164712 400 164740 5578
rect 165908 400 165936 8502
rect 169392 8492 169444 8498
rect 169392 8434 169444 8440
rect 168196 5568 168248 5574
rect 168196 5510 168248 5516
rect 167092 4208 167144 4214
rect 167092 4150 167144 4156
rect 167104 400 167132 4150
rect 168208 400 168236 5510
rect 169404 400 169432 8434
rect 169864 4826 169892 210394
rect 169956 4894 169984 210462
rect 169944 4888 169996 4894
rect 170048 4865 170076 220102
rect 170324 210458 170352 220102
rect 170692 210526 170720 220102
rect 170680 210520 170732 210526
rect 170680 210462 170732 210468
rect 170312 210452 170364 210458
rect 170312 210394 170364 210400
rect 171140 12436 171192 12442
rect 171140 12378 171192 12384
rect 169944 4830 169996 4836
rect 170034 4856 170090 4865
rect 169852 4820 169904 4826
rect 170034 4791 170090 4800
rect 170588 4820 170640 4826
rect 169852 4762 169904 4768
rect 170588 4762 170640 4768
rect 170600 400 170628 4762
rect 171152 3369 171180 12378
rect 171244 6186 171272 220102
rect 171796 212566 171824 220116
rect 172256 217297 172284 220116
rect 172638 220102 172744 220130
rect 172242 217288 172298 217297
rect 172242 217223 172298 217232
rect 171416 212560 171468 212566
rect 171416 212502 171468 212508
rect 171784 212560 171836 212566
rect 171784 212502 171836 212508
rect 171428 205630 171456 212502
rect 171416 205624 171468 205630
rect 171416 205566 171468 205572
rect 171600 205624 171652 205630
rect 171600 205566 171652 205572
rect 171612 202858 171640 205566
rect 171520 202830 171640 202858
rect 171520 196042 171548 202830
rect 171508 196036 171560 196042
rect 171508 195978 171560 195984
rect 171508 193248 171560 193254
rect 171508 193190 171560 193196
rect 171520 176474 171548 193190
rect 171428 176446 171548 176474
rect 171428 164218 171456 176446
rect 171416 164212 171468 164218
rect 171416 164154 171468 164160
rect 171600 164212 171652 164218
rect 171600 164154 171652 164160
rect 171612 154601 171640 164154
rect 171414 154592 171470 154601
rect 171414 154527 171470 154536
rect 171598 154592 171654 154601
rect 171598 154527 171654 154536
rect 171428 144906 171456 154527
rect 171416 144900 171468 144906
rect 171416 144842 171468 144848
rect 171600 144900 171652 144906
rect 171600 144842 171652 144848
rect 171612 135289 171640 144842
rect 171414 135280 171470 135289
rect 171414 135215 171470 135224
rect 171598 135280 171654 135289
rect 171598 135215 171654 135224
rect 171428 125594 171456 135215
rect 171416 125588 171468 125594
rect 171416 125530 171468 125536
rect 171416 116000 171468 116006
rect 171416 115942 171468 115948
rect 171428 106282 171456 115942
rect 171416 106276 171468 106282
rect 171416 106218 171468 106224
rect 171416 96688 171468 96694
rect 171416 96630 171468 96636
rect 171428 86970 171456 96630
rect 171416 86964 171468 86970
rect 171416 86906 171468 86912
rect 171416 77308 171468 77314
rect 171416 77250 171468 77256
rect 171428 67590 171456 77250
rect 171416 67584 171468 67590
rect 171416 67526 171468 67532
rect 171416 57996 171468 58002
rect 171416 57938 171468 57944
rect 171428 48278 171456 57938
rect 171416 48272 171468 48278
rect 171416 48214 171468 48220
rect 171416 38684 171468 38690
rect 171416 38626 171468 38632
rect 171428 28966 171456 38626
rect 171416 28960 171468 28966
rect 171416 28902 171468 28908
rect 171324 19372 171376 19378
rect 171324 19314 171376 19320
rect 171336 12442 171364 19314
rect 171324 12436 171376 12442
rect 171324 12378 171376 12384
rect 171232 6180 171284 6186
rect 171232 6122 171284 6128
rect 171784 6180 171836 6186
rect 171784 6122 171836 6128
rect 171138 3360 171194 3369
rect 171138 3295 171194 3304
rect 171796 400 171824 6122
rect 172716 4962 172744 220102
rect 172808 220102 173098 220130
rect 173176 220102 173466 220130
rect 172808 6254 172836 220102
rect 173176 210610 173204 220102
rect 173820 212566 173848 220116
rect 174096 220102 174294 220130
rect 173992 215348 174044 215354
rect 173992 215290 174044 215296
rect 173256 212560 173308 212566
rect 173254 212528 173256 212537
rect 173808 212560 173860 212566
rect 173308 212528 173310 212537
rect 173254 212463 173310 212472
rect 173438 212528 173494 212537
rect 173808 212502 173860 212508
rect 173438 212463 173494 212472
rect 172900 210582 173204 210610
rect 172796 6248 172848 6254
rect 172796 6190 172848 6196
rect 172704 4956 172756 4962
rect 172704 4898 172756 4904
rect 172900 3466 172928 210582
rect 173360 202910 173388 202941
rect 173452 202910 173480 212463
rect 173348 202904 173400 202910
rect 173440 202904 173492 202910
rect 173400 202852 173440 202858
rect 173492 202852 173572 202858
rect 173348 202846 173572 202852
rect 173360 202830 173572 202846
rect 173544 193254 173572 202830
rect 173164 193248 173216 193254
rect 173164 193190 173216 193196
rect 173532 193248 173584 193254
rect 173532 193190 173584 193196
rect 173176 173942 173204 193190
rect 173072 173936 173124 173942
rect 173072 173878 173124 173884
rect 173164 173936 173216 173942
rect 173164 173878 173216 173884
rect 173084 164218 173112 173878
rect 173072 164212 173124 164218
rect 173072 164154 173124 164160
rect 173256 164212 173308 164218
rect 173256 164154 173308 164160
rect 173268 154601 173296 164154
rect 173070 154592 173126 154601
rect 173070 154527 173126 154536
rect 173254 154592 173310 154601
rect 173254 154527 173310 154536
rect 173084 144906 173112 154527
rect 173072 144900 173124 144906
rect 173072 144842 173124 144848
rect 173256 144900 173308 144906
rect 173256 144842 173308 144848
rect 173268 135289 173296 144842
rect 173070 135280 173126 135289
rect 173070 135215 173126 135224
rect 173254 135280 173310 135289
rect 173254 135215 173310 135224
rect 173084 125594 173112 135215
rect 173072 125588 173124 125594
rect 173072 125530 173124 125536
rect 173072 116000 173124 116006
rect 173072 115942 173124 115948
rect 173084 106282 173112 115942
rect 173072 106276 173124 106282
rect 173072 106218 173124 106224
rect 173072 96688 173124 96694
rect 173072 96630 173124 96636
rect 173084 86970 173112 96630
rect 173072 86964 173124 86970
rect 173072 86906 173124 86912
rect 173072 77308 173124 77314
rect 173072 77250 173124 77256
rect 173084 67590 173112 77250
rect 173072 67584 173124 67590
rect 173072 67526 173124 67532
rect 173072 57996 173124 58002
rect 173072 57938 173124 57944
rect 173084 28966 173112 57938
rect 173072 28960 173124 28966
rect 173072 28902 173124 28908
rect 173164 28960 173216 28966
rect 173164 28902 173216 28908
rect 172980 8424 173032 8430
rect 172980 8366 173032 8372
rect 172888 3460 172940 3466
rect 172888 3402 172940 3408
rect 172992 400 173020 8366
rect 173176 3534 173204 28902
rect 174004 8974 174032 215290
rect 173992 8968 174044 8974
rect 173992 8910 174044 8916
rect 174096 5030 174124 220102
rect 174648 215354 174676 220116
rect 175108 217394 175136 220116
rect 175476 217734 175504 220116
rect 175568 220102 175950 220130
rect 176028 220102 176318 220130
rect 175464 217728 175516 217734
rect 175464 217670 175516 217676
rect 175096 217388 175148 217394
rect 175096 217330 175148 217336
rect 174636 215348 174688 215354
rect 174636 215290 174688 215296
rect 175372 210452 175424 210458
rect 175372 210394 175424 210400
rect 175384 9042 175412 210394
rect 175372 9036 175424 9042
rect 175372 8978 175424 8984
rect 175372 6248 175424 6254
rect 175372 6190 175424 6196
rect 174084 5024 174136 5030
rect 174084 4966 174136 4972
rect 174176 4888 174228 4894
rect 174176 4830 174228 4836
rect 173164 3528 173216 3534
rect 173164 3470 173216 3476
rect 174188 400 174216 4830
rect 175384 400 175412 6190
rect 175568 5098 175596 220102
rect 176028 210458 176056 220102
rect 176016 210452 176068 210458
rect 176016 210394 176068 210400
rect 176568 8968 176620 8974
rect 176568 8910 176620 8916
rect 175556 5092 175608 5098
rect 175556 5034 175608 5040
rect 176580 400 176608 8910
rect 176672 3602 176700 220116
rect 176764 220102 177146 220130
rect 177224 220102 177514 220130
rect 176764 3670 176792 220102
rect 177224 210440 177252 220102
rect 177960 212566 177988 220116
rect 178328 217326 178356 220116
rect 178788 217462 178816 220116
rect 178776 217456 178828 217462
rect 178776 217398 178828 217404
rect 178316 217320 178368 217326
rect 178316 217262 178368 217268
rect 179156 212566 179184 220116
rect 179420 213852 179472 213858
rect 179420 213794 179472 213800
rect 177304 212560 177356 212566
rect 177304 212502 177356 212508
rect 177948 212560 178000 212566
rect 177948 212502 178000 212508
rect 178868 212560 178920 212566
rect 178868 212502 178920 212508
rect 179144 212560 179196 212566
rect 179144 212502 179196 212508
rect 176856 210412 177252 210440
rect 176856 6225 176884 210412
rect 177316 195242 177344 212502
rect 177132 195214 177344 195242
rect 177132 179382 177160 195214
rect 178880 187814 178908 212502
rect 178868 187808 178920 187814
rect 178868 187750 178920 187756
rect 178224 187740 178276 187746
rect 178224 187682 178276 187688
rect 178236 186454 178264 187682
rect 178224 186448 178276 186454
rect 178224 186390 178276 186396
rect 178132 186312 178184 186318
rect 178132 186254 178184 186260
rect 177120 179376 177172 179382
rect 177120 179318 177172 179324
rect 178144 179330 178172 186254
rect 178144 179302 178264 179330
rect 178236 176746 178264 179302
rect 178052 176718 178264 176746
rect 177120 173188 177172 173194
rect 177120 173130 177172 173136
rect 177132 168366 177160 173130
rect 177120 168360 177172 168366
rect 177120 168302 177172 168308
rect 177120 158772 177172 158778
rect 177120 158714 177172 158720
rect 177132 149054 177160 158714
rect 178052 158710 178080 176718
rect 178040 158704 178092 158710
rect 178040 158646 178092 158652
rect 178132 158704 178184 158710
rect 178132 158646 178184 158652
rect 178144 149054 178172 158646
rect 177120 149048 177172 149054
rect 177120 148990 177172 148996
rect 178132 149048 178184 149054
rect 178132 148990 178184 148996
rect 177120 139528 177172 139534
rect 177120 139470 177172 139476
rect 178132 139528 178184 139534
rect 178132 139470 178184 139476
rect 177132 139398 177160 139470
rect 178144 139398 178172 139470
rect 177120 139392 177172 139398
rect 177120 139334 177172 139340
rect 178132 139392 178184 139398
rect 178132 139334 178184 139340
rect 177120 129804 177172 129810
rect 177120 129746 177172 129752
rect 178408 129804 178460 129810
rect 178408 129746 178460 129752
rect 177132 110498 177160 129746
rect 178420 122754 178448 129746
rect 178328 122726 178448 122754
rect 178328 120086 178356 122726
rect 178316 120080 178368 120086
rect 178316 120022 178368 120028
rect 176936 110492 176988 110498
rect 176936 110434 176988 110440
rect 177120 110492 177172 110498
rect 177120 110434 177172 110440
rect 178500 110492 178552 110498
rect 178500 110434 178552 110440
rect 176948 104922 176976 110434
rect 178512 106962 178540 110434
rect 178132 106956 178184 106962
rect 178132 106898 178184 106904
rect 178500 106956 178552 106962
rect 178500 106898 178552 106904
rect 176936 104916 176988 104922
rect 176936 104858 176988 104864
rect 177028 104916 177080 104922
rect 177028 104858 177080 104864
rect 177040 102134 177068 104858
rect 177028 102128 177080 102134
rect 177028 102070 177080 102076
rect 178144 102066 178172 106898
rect 177948 102060 178000 102066
rect 177948 102002 178000 102008
rect 178132 102060 178184 102066
rect 178132 102002 178184 102008
rect 177960 95146 177988 102002
rect 177960 95130 178080 95146
rect 177960 95124 178092 95130
rect 177960 95118 178040 95124
rect 178040 95066 178092 95072
rect 177120 92540 177172 92546
rect 177120 92482 177172 92488
rect 177132 85610 177160 92482
rect 178132 91112 178184 91118
rect 178132 91054 178184 91060
rect 177028 85604 177080 85610
rect 177028 85546 177080 85552
rect 177120 85604 177172 85610
rect 177120 85546 177172 85552
rect 177040 63510 177068 85546
rect 178144 81394 178172 91054
rect 178132 81388 178184 81394
rect 178132 81330 178184 81336
rect 178316 63572 178368 63578
rect 178316 63514 178368 63520
rect 177028 63504 177080 63510
rect 178328 63481 178356 63514
rect 177028 63446 177080 63452
rect 178038 63472 178094 63481
rect 178038 63407 178094 63416
rect 178314 63472 178370 63481
rect 178314 63407 178370 63416
rect 177120 57928 177172 57934
rect 177120 57870 177172 57876
rect 177132 35986 177160 57870
rect 178052 53854 178080 63407
rect 178040 53848 178092 53854
rect 178040 53790 178092 53796
rect 178132 53848 178184 53854
rect 178132 53790 178184 53796
rect 177040 35958 177160 35986
rect 178144 35970 178172 53790
rect 178132 35964 178184 35970
rect 177040 31090 177068 35958
rect 178132 35906 178184 35912
rect 178224 35964 178276 35970
rect 178224 35906 178276 35912
rect 178236 31822 178264 35906
rect 178224 31816 178276 31822
rect 178224 31758 178276 31764
rect 178132 31748 178184 31754
rect 178132 31690 178184 31696
rect 177040 31062 177160 31090
rect 177132 16726 177160 31062
rect 178144 26246 178172 31690
rect 178132 26240 178184 26246
rect 178132 26182 178184 26188
rect 177120 16720 177172 16726
rect 177120 16662 177172 16668
rect 177028 16652 177080 16658
rect 177028 16594 177080 16600
rect 178132 16652 178184 16658
rect 178132 16594 178184 16600
rect 177040 9110 177068 16594
rect 177028 9104 177080 9110
rect 177028 9046 177080 9052
rect 177764 9036 177816 9042
rect 177764 8978 177816 8984
rect 176842 6216 176898 6225
rect 176842 6151 176898 6160
rect 176752 3664 176804 3670
rect 176752 3606 176804 3612
rect 176660 3596 176712 3602
rect 176660 3538 176712 3544
rect 177776 400 177804 8978
rect 178144 6322 178172 16594
rect 178132 6316 178184 6322
rect 178132 6258 178184 6264
rect 178960 6316 179012 6322
rect 178960 6258 179012 6264
rect 178972 400 179000 6258
rect 179432 3738 179460 213794
rect 179512 210452 179564 210458
rect 179512 210394 179564 210400
rect 179524 6390 179552 210394
rect 179616 10334 179644 220116
rect 179984 213858 180012 220116
rect 180076 220102 180366 220130
rect 180826 220102 181024 220130
rect 179972 213852 180024 213858
rect 179972 213794 180024 213800
rect 180076 210458 180104 220102
rect 180156 212560 180208 212566
rect 180156 212502 180208 212508
rect 180064 210452 180116 210458
rect 180064 210394 180116 210400
rect 180168 195226 180196 212502
rect 180892 210452 180944 210458
rect 180892 210394 180944 210400
rect 180064 195220 180116 195226
rect 180064 195162 180116 195168
rect 180156 195220 180208 195226
rect 180156 195162 180208 195168
rect 180076 189038 180104 195162
rect 180064 189032 180116 189038
rect 180064 188974 180116 188980
rect 179972 179444 180024 179450
rect 179972 179386 180024 179392
rect 179984 179330 180012 179386
rect 179984 179302 180104 179330
rect 180076 176746 180104 179302
rect 179892 176718 180104 176746
rect 179892 151842 179920 176718
rect 179880 151836 179932 151842
rect 179880 151778 179932 151784
rect 179972 151836 180024 151842
rect 179972 151778 180024 151784
rect 179984 140758 180012 151778
rect 179972 140752 180024 140758
rect 179972 140694 180024 140700
rect 180156 131164 180208 131170
rect 180156 131106 180208 131112
rect 180168 127702 180196 131106
rect 179972 127696 180024 127702
rect 179972 127638 180024 127644
rect 180156 127696 180208 127702
rect 180156 127638 180208 127644
rect 179984 102134 180012 127638
rect 179972 102128 180024 102134
rect 179972 102070 180024 102076
rect 179972 92540 180024 92546
rect 179972 92482 180024 92488
rect 179984 82822 180012 92482
rect 179972 82816 180024 82822
rect 179972 82758 180024 82764
rect 179972 73228 180024 73234
rect 179972 73170 180024 73176
rect 179984 63510 180012 73170
rect 179972 63504 180024 63510
rect 179972 63446 180024 63452
rect 179972 53848 180024 53854
rect 179972 53790 180024 53796
rect 179984 45694 180012 53790
rect 179972 45688 180024 45694
rect 179972 45630 180024 45636
rect 180064 35964 180116 35970
rect 180064 35906 180116 35912
rect 180076 31822 180104 35906
rect 180064 31816 180116 31822
rect 180064 31758 180116 31764
rect 179972 31748 180024 31754
rect 179972 31690 180024 31696
rect 179984 26246 180012 31690
rect 179972 26240 180024 26246
rect 179972 26182 180024 26188
rect 179972 16652 180024 16658
rect 179972 16594 180024 16600
rect 179604 10328 179656 10334
rect 179604 10270 179656 10276
rect 179984 8702 180012 16594
rect 180156 9104 180208 9110
rect 180156 9046 180208 9052
rect 179972 8696 180024 8702
rect 179972 8638 180024 8644
rect 179512 6384 179564 6390
rect 179512 6326 179564 6332
rect 179420 3732 179472 3738
rect 179420 3674 179472 3680
rect 180168 400 180196 9046
rect 180904 6458 180932 210394
rect 180996 11762 181024 220102
rect 181180 217598 181208 220116
rect 181272 220102 181654 220130
rect 181916 220102 182022 220130
rect 182376 220102 182482 220130
rect 182560 220102 182850 220130
rect 181168 217592 181220 217598
rect 181168 217534 181220 217540
rect 181272 210458 181300 220102
rect 181916 217598 181944 220102
rect 181352 217592 181404 217598
rect 181352 217534 181404 217540
rect 181904 217592 181956 217598
rect 181904 217534 181956 217540
rect 181260 210452 181312 210458
rect 181260 210394 181312 210400
rect 181364 210338 181392 217534
rect 181180 210310 181392 210338
rect 181180 186386 181208 210310
rect 182272 205692 182324 205698
rect 182272 205634 182324 205640
rect 182284 195922 182312 205634
rect 182192 195894 182312 195922
rect 182192 186386 182220 195894
rect 181168 186380 181220 186386
rect 181168 186322 181220 186328
rect 182180 186380 182232 186386
rect 182180 186322 182232 186328
rect 181076 186312 181128 186318
rect 181076 186254 181128 186260
rect 181088 179382 181116 186254
rect 182180 182232 182232 182238
rect 182180 182174 182232 182180
rect 182192 182034 182220 182174
rect 182180 182028 182232 182034
rect 182180 181970 182232 181976
rect 181076 179376 181128 179382
rect 181076 179318 181128 179324
rect 182272 176588 182324 176594
rect 182272 176530 182324 176536
rect 182284 171086 182312 176530
rect 182272 171080 182324 171086
rect 182272 171022 182324 171028
rect 181352 169788 181404 169794
rect 181352 169730 181404 169736
rect 181364 166138 181392 169730
rect 181088 166110 181392 166138
rect 181088 161430 181116 166110
rect 182180 161492 182232 161498
rect 182180 161434 182232 161440
rect 181076 161424 181128 161430
rect 181076 161366 181128 161372
rect 182192 161362 182220 161434
rect 182180 161356 182232 161362
rect 182180 161298 182232 161304
rect 182180 156732 182232 156738
rect 182180 156674 182232 156680
rect 181076 151836 181128 151842
rect 181076 151778 181128 151784
rect 181088 142118 181116 151778
rect 182192 142118 182220 156674
rect 181076 142112 181128 142118
rect 181076 142054 181128 142060
rect 182180 142112 182232 142118
rect 182180 142054 182232 142060
rect 181168 132592 181220 132598
rect 181168 132534 181220 132540
rect 181180 132462 181208 132534
rect 181168 132456 181220 132462
rect 181168 132398 181220 132404
rect 182180 124228 182232 124234
rect 182180 124170 182232 124176
rect 181076 122868 181128 122874
rect 181076 122810 181128 122816
rect 181088 122738 181116 122810
rect 182192 122806 182220 124170
rect 182180 122800 182232 122806
rect 182180 122742 182232 122748
rect 181076 122732 181128 122738
rect 181076 122674 181128 122680
rect 182180 118040 182232 118046
rect 182180 117982 182232 117988
rect 181076 111920 181128 111926
rect 181076 111862 181128 111868
rect 181088 111790 181116 111862
rect 181076 111784 181128 111790
rect 181076 111726 181128 111732
rect 182192 109070 182220 117982
rect 182180 109064 182232 109070
rect 182180 109006 182232 109012
rect 182180 108928 182232 108934
rect 182180 108870 182232 108876
rect 182192 104786 182220 108870
rect 182180 104780 182232 104786
rect 182180 104722 182232 104728
rect 181076 102264 181128 102270
rect 181076 102206 181128 102212
rect 181088 102134 181116 102206
rect 181076 102128 181128 102134
rect 181076 102070 181128 102076
rect 181444 102128 181496 102134
rect 181444 102070 181496 102076
rect 181456 85490 181484 102070
rect 182272 99340 182324 99346
rect 182272 99282 182324 99288
rect 182284 93838 182312 99282
rect 182272 93832 182324 93838
rect 182272 93774 182324 93780
rect 181364 85462 181484 85490
rect 181364 84130 181392 85462
rect 182180 84244 182232 84250
rect 182180 84186 182232 84192
rect 181364 84102 181484 84130
rect 181456 75936 181484 84102
rect 181272 75908 181484 75936
rect 181272 74526 181300 75908
rect 181260 74520 181312 74526
rect 181260 74462 181312 74468
rect 181076 64932 181128 64938
rect 181076 64874 181128 64880
rect 181088 58682 181116 64874
rect 181076 58676 181128 58682
rect 181076 58618 181128 58624
rect 181168 53848 181220 53854
rect 181168 53790 181220 53796
rect 181180 45694 181208 53790
rect 181168 45688 181220 45694
rect 181168 45630 181220 45636
rect 181076 45620 181128 45626
rect 181076 45562 181128 45568
rect 181088 45506 181116 45562
rect 181088 45478 181392 45506
rect 181364 44130 181392 45478
rect 181352 44124 181404 44130
rect 181352 44066 181404 44072
rect 182192 41478 182220 84186
rect 182376 77246 182404 220102
rect 182560 205698 182588 220102
rect 183204 217530 183232 220116
rect 183664 217666 183692 220116
rect 183756 220102 184046 220130
rect 183652 217660 183704 217666
rect 183652 217602 183704 217608
rect 183192 217524 183244 217530
rect 183192 217466 183244 217472
rect 182548 205692 182600 205698
rect 182548 205634 182600 205640
rect 182364 77240 182416 77246
rect 182364 77182 182416 77188
rect 182364 77104 182416 77110
rect 182364 77046 182416 77052
rect 182180 41472 182232 41478
rect 182180 41414 182232 41420
rect 182180 27668 182232 27674
rect 182180 27610 182232 27616
rect 181076 26308 181128 26314
rect 181076 26250 181128 26256
rect 181088 26194 181116 26250
rect 182192 26246 182220 27610
rect 182180 26240 182232 26246
rect 181088 26178 181208 26194
rect 182180 26182 182232 26188
rect 181088 26172 181220 26178
rect 181088 26166 181168 26172
rect 181168 26114 181220 26120
rect 181352 26172 181404 26178
rect 181352 26114 181404 26120
rect 181364 17898 181392 26114
rect 182376 18018 182404 77046
rect 182456 26240 182508 26246
rect 182456 26182 182508 26188
rect 182364 18012 182416 18018
rect 182364 17954 182416 17960
rect 181272 17870 181392 17898
rect 180984 11756 181036 11762
rect 180984 11698 181036 11704
rect 181272 8362 181300 17870
rect 182364 17808 182416 17814
rect 182364 17750 182416 17756
rect 181076 8356 181128 8362
rect 181076 8298 181128 8304
rect 181260 8356 181312 8362
rect 181260 8298 181312 8304
rect 182180 8356 182232 8362
rect 182180 8298 182232 8304
rect 180892 6452 180944 6458
rect 180892 6394 180944 6400
rect 181088 3806 181116 8298
rect 182192 8242 182220 8298
rect 182192 8214 182312 8242
rect 182284 6526 182312 8214
rect 182272 6520 182324 6526
rect 182272 6462 182324 6468
rect 182376 3874 182404 17750
rect 182468 8362 182496 26182
rect 182456 8356 182508 8362
rect 182456 8298 182508 8304
rect 183756 6594 183784 220102
rect 184492 212566 184520 220116
rect 184584 220102 184874 220130
rect 185136 220102 185334 220130
rect 184020 212560 184072 212566
rect 184020 212502 184072 212508
rect 184480 212560 184532 212566
rect 184480 212502 184532 212508
rect 183836 208412 183888 208418
rect 183836 208354 183888 208360
rect 183744 6588 183796 6594
rect 183744 6530 183796 6536
rect 182548 6384 182600 6390
rect 182548 6326 182600 6332
rect 182364 3868 182416 3874
rect 182364 3810 182416 3816
rect 181076 3800 181128 3806
rect 181076 3742 181128 3748
rect 181352 3460 181404 3466
rect 181352 3402 181404 3408
rect 181364 400 181392 3402
rect 182560 400 182588 6326
rect 183848 4010 183876 208354
rect 184032 205578 184060 212502
rect 184584 208418 184612 220102
rect 184572 208412 184624 208418
rect 184572 208354 184624 208360
rect 184032 205550 184152 205578
rect 184124 201482 184152 205550
rect 184112 201476 184164 201482
rect 184112 201418 184164 201424
rect 184296 201476 184348 201482
rect 184296 201418 184348 201424
rect 184308 191865 184336 201418
rect 184018 191856 184074 191865
rect 184018 191791 184074 191800
rect 184294 191856 184350 191865
rect 184294 191791 184350 191800
rect 184032 183666 184060 191791
rect 184020 183660 184072 183666
rect 184020 183602 184072 183608
rect 184112 183660 184164 183666
rect 184112 183602 184164 183608
rect 184124 182170 184152 183602
rect 184112 182164 184164 182170
rect 184112 182106 184164 182112
rect 184204 182164 184256 182170
rect 184204 182106 184256 182112
rect 184216 169130 184244 182106
rect 184124 169102 184244 169130
rect 184124 164218 184152 169102
rect 184020 164212 184072 164218
rect 184020 164154 184072 164160
rect 184112 164212 184164 164218
rect 184112 164154 184164 164160
rect 184032 147762 184060 164154
rect 184020 147756 184072 147762
rect 184020 147698 184072 147704
rect 184020 147620 184072 147626
rect 184020 147562 184072 147568
rect 184032 135250 184060 147562
rect 183928 135244 183980 135250
rect 183928 135186 183980 135192
rect 184020 135244 184072 135250
rect 184020 135186 184072 135192
rect 183940 128330 183968 135186
rect 183940 128302 184060 128330
rect 184032 125610 184060 128302
rect 184032 125594 184152 125610
rect 183928 125588 183980 125594
rect 184032 125588 184164 125594
rect 184032 125582 184112 125588
rect 183928 125530 183980 125536
rect 184112 125530 184164 125536
rect 183940 118674 183968 125530
rect 183940 118646 184060 118674
rect 184032 115938 184060 118646
rect 184020 115932 184072 115938
rect 184020 115874 184072 115880
rect 184112 108860 184164 108866
rect 184112 108802 184164 108808
rect 184124 99498 184152 108802
rect 184124 99470 184244 99498
rect 184216 99362 184244 99470
rect 184124 99334 184244 99362
rect 184124 75970 184152 99334
rect 184032 75942 184152 75970
rect 184032 75886 184060 75942
rect 184020 75880 184072 75886
rect 184020 75822 184072 75828
rect 184112 66292 184164 66298
rect 184112 66234 184164 66240
rect 184124 57934 184152 66234
rect 183928 57928 183980 57934
rect 183928 57870 183980 57876
rect 184112 57928 184164 57934
rect 184112 57870 184164 57876
rect 183940 55214 183968 57870
rect 183928 55208 183980 55214
rect 183928 55150 183980 55156
rect 183928 45620 183980 45626
rect 183928 45562 183980 45568
rect 183940 38706 183968 45562
rect 183940 38678 184060 38706
rect 184032 33810 184060 38678
rect 184032 33782 184244 33810
rect 184216 31634 184244 33782
rect 184124 31606 184244 31634
rect 184124 28966 184152 31606
rect 184020 28960 184072 28966
rect 184020 28902 184072 28908
rect 184112 28960 184164 28966
rect 184112 28902 184164 28908
rect 184032 9602 184060 28902
rect 183940 9574 184060 9602
rect 183836 4004 183888 4010
rect 183836 3946 183888 3952
rect 183940 3942 183968 9574
rect 185136 6662 185164 220102
rect 185688 217802 185716 220116
rect 185676 217796 185728 217802
rect 185676 217738 185728 217744
rect 186148 216782 186176 220116
rect 186136 216776 186188 216782
rect 186136 216718 186188 216724
rect 185584 216708 185636 216714
rect 185584 216650 185636 216656
rect 185124 6656 185176 6662
rect 185124 6598 185176 6604
rect 185596 4078 185624 216650
rect 186412 210452 186464 210458
rect 186412 210394 186464 210400
rect 186424 6730 186452 210394
rect 186412 6724 186464 6730
rect 186412 6666 186464 6672
rect 186044 6452 186096 6458
rect 186044 6394 186096 6400
rect 185584 4072 185636 4078
rect 185584 4014 185636 4020
rect 183928 3936 183980 3942
rect 183928 3878 183980 3884
rect 183744 3596 183796 3602
rect 183744 3538 183796 3544
rect 183756 400 183784 3538
rect 184848 3528 184900 3534
rect 184848 3470 184900 3476
rect 184860 400 184888 3470
rect 186056 400 186084 6394
rect 186516 5166 186544 220116
rect 186608 220102 186898 220130
rect 186608 210458 186636 220102
rect 187344 217870 187372 220116
rect 187726 220102 187832 220130
rect 187332 217864 187384 217870
rect 187332 217806 187384 217812
rect 186964 217524 187016 217530
rect 186964 217466 187016 217472
rect 186596 210452 186648 210458
rect 186596 210394 186648 210400
rect 186504 5160 186556 5166
rect 186504 5102 186556 5108
rect 186976 4146 187004 217466
rect 187804 5234 187832 220102
rect 187896 220102 188186 220130
rect 187896 7585 187924 220102
rect 188344 217660 188396 217666
rect 188344 217602 188396 217608
rect 187976 210452 188028 210458
rect 187976 210394 188028 210400
rect 187882 7576 187938 7585
rect 187882 7511 187938 7520
rect 187988 5302 188016 210394
rect 187976 5296 188028 5302
rect 187976 5238 188028 5244
rect 187792 5228 187844 5234
rect 187792 5170 187844 5176
rect 187240 4956 187292 4962
rect 187240 4898 187292 4904
rect 186964 4140 187016 4146
rect 186964 4082 187016 4088
rect 187252 400 187280 4898
rect 188356 3398 188384 217602
rect 188540 216714 188568 220116
rect 188632 220102 189014 220130
rect 189184 220102 189382 220130
rect 188528 216708 188580 216714
rect 188528 216650 188580 216656
rect 188632 210458 188660 220102
rect 188620 210452 188672 210458
rect 188620 210394 188672 210400
rect 189184 7614 189212 220102
rect 189736 217258 189764 220116
rect 189724 217252 189776 217258
rect 189724 217194 189776 217200
rect 190196 212566 190224 220116
rect 189356 212560 189408 212566
rect 189356 212502 189408 212508
rect 190184 212560 190236 212566
rect 190184 212502 190236 212508
rect 189368 205578 189396 212502
rect 189368 205550 189488 205578
rect 189460 186386 189488 205550
rect 189448 186380 189500 186386
rect 189448 186322 189500 186328
rect 189540 186244 189592 186250
rect 189540 186186 189592 186192
rect 189552 172582 189580 186186
rect 189448 172576 189500 172582
rect 189448 172518 189500 172524
rect 189540 172576 189592 172582
rect 189540 172518 189592 172524
rect 189460 164218 189488 172518
rect 189356 164212 189408 164218
rect 189356 164154 189408 164160
rect 189448 164212 189500 164218
rect 189448 164154 189500 164160
rect 189368 147762 189396 164154
rect 189356 147756 189408 147762
rect 189356 147698 189408 147704
rect 189356 147620 189408 147626
rect 189356 147562 189408 147568
rect 189368 128382 189396 147562
rect 189356 128376 189408 128382
rect 189356 128318 189408 128324
rect 189448 128308 189500 128314
rect 189448 128250 189500 128256
rect 189460 116113 189488 128250
rect 189446 116104 189502 116113
rect 189446 116039 189502 116048
rect 189354 115968 189410 115977
rect 189354 115903 189356 115912
rect 189408 115903 189410 115912
rect 189448 115932 189500 115938
rect 189356 115874 189408 115880
rect 189448 115874 189500 115880
rect 189460 99498 189488 115874
rect 189460 99470 189580 99498
rect 189552 99362 189580 99470
rect 189460 99334 189580 99362
rect 189460 75954 189488 99334
rect 189356 75948 189408 75954
rect 189356 75890 189408 75896
rect 189448 75948 189500 75954
rect 189448 75890 189500 75896
rect 189368 53122 189396 75890
rect 189368 53094 189488 53122
rect 189460 48278 189488 53094
rect 189448 48272 189500 48278
rect 189448 48214 189500 48220
rect 189540 48272 189592 48278
rect 189540 48214 189592 48220
rect 189552 40730 189580 48214
rect 189540 40724 189592 40730
rect 189540 40666 189592 40672
rect 189540 27668 189592 27674
rect 189540 27610 189592 27616
rect 189552 9722 189580 27610
rect 189264 9716 189316 9722
rect 189264 9658 189316 9664
rect 189540 9716 189592 9722
rect 189540 9658 189592 9664
rect 189276 9602 189304 9658
rect 189276 9574 189396 9602
rect 189172 7608 189224 7614
rect 189172 7550 189224 7556
rect 189368 5370 189396 9574
rect 190564 7682 190592 220116
rect 191024 217530 191052 220116
rect 191116 220102 191406 220130
rect 191866 220102 191972 220130
rect 191012 217524 191064 217530
rect 191012 217466 191064 217472
rect 191116 210474 191144 220102
rect 191196 217796 191248 217802
rect 191196 217738 191248 217744
rect 190656 210446 191144 210474
rect 190552 7676 190604 7682
rect 190552 7618 190604 7624
rect 190656 5438 190684 210446
rect 191208 208298 191236 217738
rect 191116 208270 191236 208298
rect 191116 196058 191144 208270
rect 191024 196030 191144 196058
rect 191024 195922 191052 196030
rect 191024 195894 191144 195922
rect 191116 167090 191144 195894
rect 191024 167062 191144 167090
rect 191024 166954 191052 167062
rect 191024 166926 191144 166954
rect 191116 154737 191144 166926
rect 191102 154728 191158 154737
rect 191102 154663 191158 154672
rect 191102 154592 191158 154601
rect 191102 154527 191158 154536
rect 191116 153202 191144 154527
rect 191104 153196 191156 153202
rect 191104 153138 191156 153144
rect 191196 153196 191248 153202
rect 191196 153138 191248 153144
rect 191208 139890 191236 153138
rect 191116 139862 191236 139890
rect 191116 128450 191144 139862
rect 191104 128444 191156 128450
rect 191104 128386 191156 128392
rect 191012 128308 191064 128314
rect 191012 128250 191064 128256
rect 191024 125594 191052 128250
rect 191012 125588 191064 125594
rect 191012 125530 191064 125536
rect 191196 125588 191248 125594
rect 191196 125530 191248 125536
rect 191208 120578 191236 125530
rect 191116 120550 191236 120578
rect 191116 106457 191144 120550
rect 191102 106448 191158 106457
rect 191102 106383 191158 106392
rect 191010 106312 191066 106321
rect 191010 106247 191066 106256
rect 191024 95266 191052 106247
rect 191012 95260 191064 95266
rect 191012 95202 191064 95208
rect 191196 95260 191248 95266
rect 191196 95202 191248 95208
rect 191208 87038 191236 95202
rect 191196 87032 191248 87038
rect 191196 86974 191248 86980
rect 191104 86964 191156 86970
rect 191104 86906 191156 86912
rect 191116 84182 191144 86906
rect 191104 84176 191156 84182
rect 191104 84118 191156 84124
rect 191288 74588 191340 74594
rect 191288 74530 191340 74536
rect 191300 74474 191328 74530
rect 191116 74446 191328 74474
rect 191116 65113 191144 74446
rect 191102 65104 191158 65113
rect 191102 65039 191158 65048
rect 191010 64968 191066 64977
rect 191066 64926 191144 64954
rect 191010 64903 191066 64912
rect 191116 54097 191144 64926
rect 191102 54088 191158 54097
rect 191102 54023 191158 54032
rect 191102 53952 191158 53961
rect 191102 53887 191158 53896
rect 191116 53825 191144 53887
rect 190918 53816 190974 53825
rect 190918 53751 190974 53760
rect 191102 53816 191158 53825
rect 191102 53751 191158 53760
rect 190932 44198 190960 53751
rect 191116 44198 191144 44229
rect 190920 44192 190972 44198
rect 190920 44134 190972 44140
rect 191104 44192 191156 44198
rect 191156 44140 191236 44146
rect 191104 44134 191236 44140
rect 191116 44118 191236 44134
rect 191208 38690 191236 44118
rect 191196 38684 191248 38690
rect 191196 38626 191248 38632
rect 191104 38616 191156 38622
rect 191104 38558 191156 38564
rect 191116 12458 191144 38558
rect 191024 12430 191144 12458
rect 190644 5432 190696 5438
rect 190644 5374 190696 5380
rect 189356 5364 189408 5370
rect 189356 5306 189408 5312
rect 190828 5024 190880 5030
rect 190828 4966 190880 4972
rect 189632 3732 189684 3738
rect 189632 3674 189684 3680
rect 188436 3664 188488 3670
rect 188436 3606 188488 3612
rect 188344 3392 188396 3398
rect 188344 3334 188396 3340
rect 188448 400 188476 3606
rect 189644 400 189672 3674
rect 190840 400 190868 4966
rect 191024 3330 191052 12430
rect 191944 7750 191972 220102
rect 192220 217326 192248 220116
rect 192208 217320 192260 217326
rect 192208 217262 192260 217268
rect 192484 217320 192536 217326
rect 192484 217262 192536 217268
rect 192392 212560 192444 212566
rect 192392 212502 192444 212508
rect 192024 210452 192076 210458
rect 192024 210394 192076 210400
rect 192036 9178 192064 210394
rect 192404 201482 192432 212502
rect 192392 201476 192444 201482
rect 192392 201418 192444 201424
rect 192116 193180 192168 193186
rect 192116 193122 192168 193128
rect 192128 183598 192156 193122
rect 192116 183592 192168 183598
rect 192116 183534 192168 183540
rect 192208 183592 192260 183598
rect 192208 183534 192260 183540
rect 192220 182170 192248 183534
rect 192208 182164 192260 182170
rect 192208 182106 192260 182112
rect 192208 176112 192260 176118
rect 192208 176054 192260 176060
rect 192220 156806 192248 176054
rect 192208 156800 192260 156806
rect 192208 156742 192260 156748
rect 192116 153264 192168 153270
rect 192168 153212 192248 153218
rect 192116 153206 192248 153212
rect 192128 153190 192248 153206
rect 192220 124166 192248 153190
rect 192208 124160 192260 124166
rect 192208 124102 192260 124108
rect 192300 124160 192352 124166
rect 192300 124102 192352 124108
rect 192312 122806 192340 124102
rect 192300 122800 192352 122806
rect 192300 122742 192352 122748
rect 192392 110424 192444 110430
rect 192392 110366 192444 110372
rect 192404 95266 192432 110366
rect 192392 95260 192444 95266
rect 192392 95202 192444 95208
rect 192392 95124 192444 95130
rect 192392 95066 192444 95072
rect 192404 90438 192432 95066
rect 192116 90432 192168 90438
rect 192116 90374 192168 90380
rect 192392 90432 192444 90438
rect 192392 90374 192444 90380
rect 192128 85626 192156 90374
rect 192128 85598 192248 85626
rect 192220 84182 192248 85598
rect 192208 84176 192260 84182
rect 192208 84118 192260 84124
rect 192208 66292 192260 66298
rect 192208 66234 192260 66240
rect 192220 51134 192248 66234
rect 192208 51128 192260 51134
rect 192208 51070 192260 51076
rect 192116 51060 192168 51066
rect 192116 51002 192168 51008
rect 192128 42106 192156 51002
rect 192128 42078 192340 42106
rect 192312 26058 192340 42078
rect 192220 26030 192340 26058
rect 192220 19310 192248 26030
rect 192208 19304 192260 19310
rect 192208 19246 192260 19252
rect 192116 9716 192168 9722
rect 192116 9658 192168 9664
rect 192024 9172 192076 9178
rect 192024 9114 192076 9120
rect 191932 7744 191984 7750
rect 191932 7686 191984 7692
rect 192128 5506 192156 9658
rect 192116 5500 192168 5506
rect 192116 5442 192168 5448
rect 192024 3868 192076 3874
rect 192024 3810 192076 3816
rect 191012 3324 191064 3330
rect 191012 3266 191064 3272
rect 192036 400 192064 3810
rect 192496 3194 192524 217262
rect 192576 217252 192628 217258
rect 192576 217194 192628 217200
rect 192588 3262 192616 217194
rect 192680 212566 192708 220116
rect 192772 220102 193062 220130
rect 192668 212560 192720 212566
rect 192668 212502 192720 212508
rect 192772 210458 192800 220102
rect 193416 217666 193444 220116
rect 193508 220102 193890 220130
rect 193968 220102 194258 220130
rect 193404 217660 193456 217666
rect 193404 217602 193456 217608
rect 192760 210452 192812 210458
rect 192760 210394 192812 210400
rect 193312 210452 193364 210458
rect 193312 210394 193364 210400
rect 193324 10402 193352 210394
rect 193312 10396 193364 10402
rect 193312 10338 193364 10344
rect 193508 4758 193536 220102
rect 193864 212900 193916 212906
rect 193864 212842 193916 212848
rect 193496 4752 193548 4758
rect 193496 4694 193548 4700
rect 193220 3800 193272 3806
rect 193220 3742 193272 3748
rect 192576 3256 192628 3262
rect 192576 3198 192628 3204
rect 192484 3188 192536 3194
rect 192484 3130 192536 3136
rect 193232 400 193260 3742
rect 193876 3126 193904 212842
rect 193968 210458 193996 220102
rect 194704 217938 194732 220116
rect 194796 220102 195086 220130
rect 194692 217932 194744 217938
rect 194692 217874 194744 217880
rect 194692 216368 194744 216374
rect 194692 216310 194744 216316
rect 194704 210934 194732 216310
rect 194692 210928 194744 210934
rect 194692 210870 194744 210876
rect 193956 210452 194008 210458
rect 193956 210394 194008 210400
rect 194796 6798 194824 220102
rect 195428 217660 195480 217666
rect 195428 217602 195480 217608
rect 195244 217592 195296 217598
rect 195244 217534 195296 217540
rect 195152 210928 195204 210934
rect 195152 210870 195204 210876
rect 195164 191842 195192 210870
rect 194980 191814 195192 191842
rect 194980 186946 195008 191814
rect 194980 186918 195100 186946
rect 195072 172582 195100 186918
rect 194968 172576 195020 172582
rect 194968 172518 195020 172524
rect 195060 172576 195112 172582
rect 195060 172518 195112 172524
rect 194980 154737 195008 172518
rect 194966 154728 195022 154737
rect 194966 154663 195022 154672
rect 194966 154592 195022 154601
rect 194966 154527 195022 154536
rect 194980 143585 195008 154527
rect 194966 143576 195022 143585
rect 194966 143511 195022 143520
rect 194966 142216 195022 142225
rect 194966 142151 195022 142160
rect 194980 140758 195008 142151
rect 194968 140752 195020 140758
rect 194968 140694 195020 140700
rect 194876 131164 194928 131170
rect 194876 131106 194928 131112
rect 194888 124234 194916 131106
rect 194876 124228 194928 124234
rect 194876 124170 194928 124176
rect 194968 124228 195020 124234
rect 194968 124170 195020 124176
rect 194980 116006 195008 124170
rect 194968 116000 195020 116006
rect 194968 115942 195020 115948
rect 194876 115932 194928 115938
rect 194876 115874 194928 115880
rect 194888 114510 194916 115874
rect 194876 114504 194928 114510
rect 194876 114446 194928 114452
rect 194968 104916 195020 104922
rect 194968 104858 195020 104864
rect 194980 95198 195008 104858
rect 194968 95192 195020 95198
rect 194968 95134 195020 95140
rect 194876 85604 194928 85610
rect 194876 85546 194928 85552
rect 194888 77246 194916 85546
rect 194876 77240 194928 77246
rect 194876 77182 194928 77188
rect 194968 66292 195020 66298
rect 194968 66234 195020 66240
rect 194980 66201 195008 66234
rect 194966 66192 195022 66201
rect 194966 66127 195022 66136
rect 194874 57896 194930 57905
rect 194874 57831 194930 57840
rect 194888 53122 194916 57831
rect 194888 53094 195008 53122
rect 194980 46918 195008 53094
rect 194968 46912 195020 46918
rect 194968 46854 195020 46860
rect 195152 46912 195204 46918
rect 195152 46854 195204 46860
rect 195164 37369 195192 46854
rect 195150 37360 195206 37369
rect 195150 37295 195206 37304
rect 194874 37224 194930 37233
rect 194874 37159 194930 37168
rect 194888 26246 194916 37159
rect 194876 26240 194928 26246
rect 194876 26182 194928 26188
rect 194968 16652 195020 16658
rect 194968 16594 195020 16600
rect 194980 12458 195008 16594
rect 194888 12430 195008 12458
rect 194888 10470 194916 12430
rect 194876 10464 194928 10470
rect 194876 10406 194928 10412
rect 194784 6792 194836 6798
rect 194784 6734 194836 6740
rect 194416 5092 194468 5098
rect 194416 5034 194468 5040
rect 193864 3120 193916 3126
rect 193864 3062 193916 3068
rect 194428 400 194456 5034
rect 195256 2990 195284 217534
rect 195336 217524 195388 217530
rect 195336 217466 195388 217472
rect 195348 3058 195376 217466
rect 195336 3052 195388 3058
rect 195336 2994 195388 3000
rect 195244 2984 195296 2990
rect 195244 2926 195296 2932
rect 195440 2922 195468 217602
rect 195532 216374 195560 220116
rect 195900 217802 195928 220116
rect 196176 220102 196282 220130
rect 196360 220102 196742 220130
rect 195888 217796 195940 217802
rect 195888 217738 195940 217744
rect 195520 216368 195572 216374
rect 195520 216310 195572 216316
rect 196072 205692 196124 205698
rect 196072 205634 196124 205640
rect 196084 196058 196112 205634
rect 195992 196030 196112 196058
rect 195992 195922 196020 196030
rect 195992 195894 196112 195922
rect 196084 167090 196112 195894
rect 195992 167062 196112 167090
rect 195992 166954 196020 167062
rect 195992 166926 196112 166954
rect 196084 147778 196112 166926
rect 195992 147750 196112 147778
rect 195992 147642 196020 147750
rect 195992 147614 196112 147642
rect 196084 128466 196112 147614
rect 195992 128438 196112 128466
rect 195992 128330 196020 128438
rect 195992 128302 196112 128330
rect 196084 109154 196112 128302
rect 195992 109126 196112 109154
rect 195992 109018 196020 109126
rect 195992 108990 196112 109018
rect 196084 89842 196112 108990
rect 195992 89814 196112 89842
rect 195992 89706 196020 89814
rect 195992 89678 196112 89706
rect 196084 70394 196112 89678
rect 195992 70366 196112 70394
rect 195992 70258 196020 70366
rect 195992 70230 196112 70258
rect 196084 51082 196112 70230
rect 195992 51054 196112 51082
rect 195992 50946 196020 51054
rect 195992 50918 196112 50946
rect 196084 31890 196112 50918
rect 196072 31884 196124 31890
rect 196072 31826 196124 31832
rect 196072 31748 196124 31754
rect 196072 31690 196124 31696
rect 196084 12458 196112 31690
rect 195992 12430 196112 12458
rect 195992 10538 196020 12430
rect 195980 10532 196032 10538
rect 195980 10474 196032 10480
rect 196176 7818 196204 220102
rect 196360 205698 196388 220102
rect 197096 218006 197124 220116
rect 197084 218000 197136 218006
rect 197084 217942 197136 217948
rect 196624 217932 196676 217938
rect 196624 217874 196676 217880
rect 196348 205692 196400 205698
rect 196348 205634 196400 205640
rect 196164 7812 196216 7818
rect 196164 7754 196216 7760
rect 195612 3936 195664 3942
rect 195612 3878 195664 3884
rect 195428 2916 195480 2922
rect 195428 2858 195480 2864
rect 195624 400 195652 3878
rect 196636 2854 196664 217874
rect 197452 205760 197504 205766
rect 197452 205702 197504 205708
rect 197464 10606 197492 205702
rect 197452 10600 197504 10606
rect 197452 10542 197504 10548
rect 197556 7886 197584 220116
rect 197648 220102 197938 220130
rect 197648 205766 197676 220102
rect 198384 217258 198412 220116
rect 198372 217252 198424 217258
rect 198372 217194 198424 217200
rect 197636 205760 197688 205766
rect 197636 205702 197688 205708
rect 198752 7954 198780 220116
rect 198936 220102 199226 220130
rect 198832 208344 198884 208350
rect 198832 208286 198884 208292
rect 198844 8022 198872 208286
rect 198936 10674 198964 220102
rect 199580 217326 199608 220116
rect 199672 220102 199962 220130
rect 200224 220102 200422 220130
rect 199568 217320 199620 217326
rect 199568 217262 199620 217268
rect 199672 208350 199700 220102
rect 199660 208344 199712 208350
rect 199660 208286 199712 208292
rect 200224 10742 200252 220102
rect 200776 217190 200804 220116
rect 200764 217184 200816 217190
rect 200764 217126 200816 217132
rect 201236 212566 201264 220116
rect 201408 217320 201460 217326
rect 201408 217262 201460 217268
rect 200856 212560 200908 212566
rect 200856 212502 200908 212508
rect 201224 212560 201276 212566
rect 201224 212502 201276 212508
rect 200868 198098 200896 212502
rect 200500 198070 200896 198098
rect 200500 176746 200528 198070
rect 200408 176718 200528 176746
rect 200408 154737 200436 176718
rect 200394 154728 200450 154737
rect 200394 154663 200450 154672
rect 200394 154592 200450 154601
rect 200394 154527 200450 154536
rect 200408 147762 200436 154527
rect 200396 147756 200448 147762
rect 200396 147698 200448 147704
rect 200396 147620 200448 147626
rect 200396 147562 200448 147568
rect 200408 135425 200436 147562
rect 200394 135416 200450 135425
rect 200394 135351 200450 135360
rect 200394 135280 200450 135289
rect 200394 135215 200450 135224
rect 200408 129010 200436 135215
rect 200316 128982 200436 129010
rect 200316 124166 200344 128982
rect 200304 124160 200356 124166
rect 200304 124102 200356 124108
rect 200580 115864 200632 115870
rect 200580 115806 200632 115812
rect 200592 96665 200620 115806
rect 200394 96656 200450 96665
rect 200394 96591 200450 96600
rect 200578 96656 200634 96665
rect 200578 96591 200634 96600
rect 200408 85678 200436 96591
rect 200396 85672 200448 85678
rect 200396 85614 200448 85620
rect 200304 85604 200356 85610
rect 200304 85546 200356 85552
rect 200316 77314 200344 85546
rect 200304 77308 200356 77314
rect 200304 77250 200356 77256
rect 200396 77308 200448 77314
rect 200396 77250 200448 77256
rect 200408 61470 200436 77250
rect 200396 61464 200448 61470
rect 200396 61406 200448 61412
rect 200488 48340 200540 48346
rect 200488 48282 200540 48288
rect 200500 37330 200528 48282
rect 200396 37324 200448 37330
rect 200396 37266 200448 37272
rect 200488 37324 200540 37330
rect 200488 37266 200540 37272
rect 200408 27674 200436 37266
rect 200396 27668 200448 27674
rect 200396 27610 200448 27616
rect 200396 26308 200448 26314
rect 200396 26250 200448 26256
rect 200408 22166 200436 26250
rect 200396 22160 200448 22166
rect 200396 22102 200448 22108
rect 200396 22024 200448 22030
rect 200396 21966 200448 21972
rect 200212 10736 200264 10742
rect 200212 10678 200264 10684
rect 198924 10668 198976 10674
rect 198924 10610 198976 10616
rect 200408 8090 200436 21966
rect 200396 8084 200448 8090
rect 200396 8026 200448 8032
rect 198832 8016 198884 8022
rect 198832 7958 198884 7964
rect 198740 7948 198792 7954
rect 198740 7890 198792 7896
rect 197544 7880 197596 7886
rect 197544 7822 197596 7828
rect 198004 5160 198056 5166
rect 198004 5102 198056 5108
rect 196808 3256 196860 3262
rect 196808 3198 196860 3204
rect 196624 2848 196676 2854
rect 196624 2790 196676 2796
rect 196820 400 196848 3198
rect 198016 400 198044 5102
rect 199200 4140 199252 4146
rect 199200 4082 199252 4088
rect 199212 400 199240 4082
rect 201420 3126 201448 217262
rect 201500 39976 201552 39982
rect 201498 39944 201500 39953
rect 201552 39944 201554 39953
rect 201498 39879 201554 39888
rect 201604 10810 201632 220116
rect 202064 212906 202092 220116
rect 202052 212900 202104 212906
rect 202052 212842 202104 212848
rect 202432 212566 202460 220116
rect 202524 220102 202814 220130
rect 201868 212560 201920 212566
rect 201868 212502 201920 212508
rect 202420 212560 202472 212566
rect 202420 212502 202472 212508
rect 201684 210452 201736 210458
rect 201684 210394 201736 210400
rect 201696 10878 201724 210394
rect 201880 205578 201908 212502
rect 202524 210458 202552 220102
rect 203260 217054 203288 220116
rect 203524 217456 203576 217462
rect 203524 217398 203576 217404
rect 203248 217048 203300 217054
rect 203248 216990 203300 216996
rect 203432 212560 203484 212566
rect 203432 212502 203484 212508
rect 202512 210452 202564 210458
rect 202512 210394 202564 210400
rect 202972 210452 203024 210458
rect 202972 210394 203024 210400
rect 201880 205550 202000 205578
rect 201972 176746 202000 205550
rect 201880 176718 202000 176746
rect 201880 154737 201908 176718
rect 201866 154728 201922 154737
rect 201866 154663 201922 154672
rect 201866 154592 201922 154601
rect 201866 154527 201922 154536
rect 201880 147762 201908 154527
rect 201868 147756 201920 147762
rect 201868 147698 201920 147704
rect 201868 147620 201920 147626
rect 201868 147562 201920 147568
rect 201880 135425 201908 147562
rect 201866 135416 201922 135425
rect 201866 135351 201922 135360
rect 201866 135280 201922 135289
rect 201866 135215 201922 135224
rect 201880 133890 201908 135215
rect 201868 133884 201920 133890
rect 201868 133826 201920 133832
rect 201776 124228 201828 124234
rect 201776 124170 201828 124176
rect 201788 116006 201816 124170
rect 201776 116000 201828 116006
rect 201776 115942 201828 115948
rect 201868 116000 201920 116006
rect 201868 115942 201920 115948
rect 201880 114510 201908 115942
rect 201868 114504 201920 114510
rect 201868 114446 201920 114452
rect 202052 104916 202104 104922
rect 202052 104858 202104 104864
rect 202064 96665 202092 104858
rect 201866 96656 201922 96665
rect 201866 96591 201922 96600
rect 202050 96656 202106 96665
rect 202050 96591 202106 96600
rect 201880 86970 201908 96591
rect 201868 86964 201920 86970
rect 201868 86906 201920 86912
rect 201868 77308 201920 77314
rect 201868 77250 201920 77256
rect 201880 61470 201908 77250
rect 201868 61464 201920 61470
rect 201868 61406 201920 61412
rect 202052 53984 202104 53990
rect 202052 53926 202104 53932
rect 202064 47002 202092 53926
rect 201972 46974 202092 47002
rect 201972 45558 202000 46974
rect 201960 45552 202012 45558
rect 201960 45494 202012 45500
rect 201866 40080 201922 40089
rect 201866 40015 201922 40024
rect 201880 39982 201908 40015
rect 201868 39976 201920 39982
rect 201868 39918 201920 39924
rect 201868 27668 201920 27674
rect 201868 27610 201920 27616
rect 201684 10872 201736 10878
rect 201684 10814 201736 10820
rect 201592 10804 201644 10810
rect 201592 10746 201644 10752
rect 201880 8158 201908 27610
rect 202984 10946 203012 210394
rect 203444 202858 203472 212502
rect 203352 202830 203472 202858
rect 203352 193254 203380 202830
rect 203248 193248 203300 193254
rect 203248 193190 203300 193196
rect 203340 193248 203392 193254
rect 203340 193190 203392 193196
rect 203260 171154 203288 193190
rect 203156 171148 203208 171154
rect 203156 171090 203208 171096
rect 203248 171148 203300 171154
rect 203248 171090 203300 171096
rect 203168 161430 203196 171090
rect 203156 161424 203208 161430
rect 203156 161366 203208 161372
rect 203156 144900 203208 144906
rect 203156 144842 203208 144848
rect 203168 143562 203196 144842
rect 203168 143534 203288 143562
rect 203260 134026 203288 143534
rect 203248 134020 203300 134026
rect 203248 133962 203300 133968
rect 203064 132524 203116 132530
rect 203064 132466 203116 132472
rect 203076 124166 203104 132466
rect 203064 124160 203116 124166
rect 203064 124102 203116 124108
rect 203248 114572 203300 114578
rect 203248 114514 203300 114520
rect 203260 96642 203288 114514
rect 203168 96614 203288 96642
rect 203168 87145 203196 96614
rect 203154 87136 203210 87145
rect 203154 87071 203210 87080
rect 203062 87000 203118 87009
rect 203062 86935 203118 86944
rect 203076 80714 203104 86935
rect 203064 80708 203116 80714
rect 203064 80650 203116 80656
rect 203064 71120 203116 71126
rect 203064 71062 203116 71068
rect 203076 66230 203104 71062
rect 203064 66224 203116 66230
rect 203064 66166 203116 66172
rect 203340 66224 203392 66230
rect 203340 66166 203392 66172
rect 203352 64870 203380 66166
rect 203340 64864 203392 64870
rect 203340 64806 203392 64812
rect 203064 55276 203116 55282
rect 203064 55218 203116 55224
rect 203076 38706 203104 55218
rect 203076 38678 203196 38706
rect 203168 28966 203196 38678
rect 203156 28960 203208 28966
rect 203156 28902 203208 28908
rect 203248 28960 203300 28966
rect 203248 28902 203300 28908
rect 203260 22012 203288 28902
rect 203168 21984 203288 22012
rect 202972 10940 203024 10946
rect 202972 10882 203024 10888
rect 203168 8226 203196 21984
rect 203156 8220 203208 8226
rect 203156 8162 203208 8168
rect 201868 8152 201920 8158
rect 201868 8094 201920 8100
rect 201500 5228 201552 5234
rect 201500 5170 201552 5176
rect 200396 3120 200448 3126
rect 200396 3062 200448 3068
rect 201408 3120 201460 3126
rect 201408 3062 201460 3068
rect 200408 400 200436 3062
rect 201512 400 201540 5170
rect 203536 4146 203564 217398
rect 203628 212566 203656 220116
rect 203720 220102 204102 220130
rect 203616 212560 203668 212566
rect 203616 212502 203668 212508
rect 203720 210458 203748 220102
rect 204456 217530 204484 220116
rect 204548 220102 204930 220130
rect 205008 220102 205298 220130
rect 204444 217524 204496 217530
rect 204444 217466 204496 217472
rect 204168 217388 204220 217394
rect 204168 217330 204220 217336
rect 203708 210452 203760 210458
rect 203708 210394 203760 210400
rect 203524 4140 203576 4146
rect 203524 4082 203576 4088
rect 202696 3120 202748 3126
rect 202696 3062 202748 3068
rect 202708 400 202736 3062
rect 204180 490 204208 217330
rect 204352 210452 204404 210458
rect 204352 210394 204404 210400
rect 204364 11014 204392 210394
rect 204352 11008 204404 11014
rect 204352 10950 204404 10956
rect 204548 8294 204576 220102
rect 204904 217524 204956 217530
rect 204904 217466 204956 217472
rect 204536 8288 204588 8294
rect 204536 8230 204588 8236
rect 204916 3262 204944 217466
rect 205008 210458 205036 220102
rect 205652 217122 205680 220116
rect 205836 220102 206126 220130
rect 206204 220102 206494 220130
rect 205640 217116 205692 217122
rect 205640 217058 205692 217064
rect 205732 214600 205784 214606
rect 205732 214542 205784 214548
rect 204996 210452 205048 210458
rect 204996 210394 205048 210400
rect 205744 10266 205772 214542
rect 205732 10260 205784 10266
rect 205732 10202 205784 10208
rect 205836 7546 205864 220102
rect 206204 214606 206232 220102
rect 206940 217598 206968 220116
rect 207216 220102 207322 220130
rect 207400 220102 207782 220130
rect 206928 217592 206980 217598
rect 206928 217534 206980 217540
rect 206192 214600 206244 214606
rect 206192 214542 206244 214548
rect 207112 209840 207164 209846
rect 207112 209782 207164 209788
rect 207124 10198 207152 209782
rect 207112 10192 207164 10198
rect 207112 10134 207164 10140
rect 205824 7540 205876 7546
rect 205824 7482 205876 7488
rect 207216 7478 207244 220102
rect 207400 209846 207428 220102
rect 208136 216986 208164 220116
rect 208308 217592 208360 217598
rect 208308 217534 208360 217540
rect 208124 216980 208176 216986
rect 208124 216922 208176 216928
rect 207388 209840 207440 209846
rect 207388 209782 207440 209788
rect 207204 7472 207256 7478
rect 207204 7414 207256 7420
rect 205088 5296 205140 5302
rect 205088 5238 205140 5244
rect 204904 3256 204956 3262
rect 204904 3198 204956 3204
rect 203904 462 204208 490
rect 203904 400 203932 462
rect 205100 400 205128 5238
rect 206284 4072 206336 4078
rect 206284 4014 206336 4020
rect 206296 400 206324 4014
rect 208320 3194 208348 217534
rect 208492 214600 208544 214606
rect 208492 214542 208544 214548
rect 208504 10130 208532 214542
rect 208492 10124 208544 10130
rect 208492 10066 208544 10072
rect 208596 7410 208624 220116
rect 208688 220102 208978 220130
rect 208688 214606 208716 220102
rect 209044 217796 209096 217802
rect 209044 217738 209096 217744
rect 208676 214600 208728 214606
rect 208676 214542 208728 214548
rect 208584 7404 208636 7410
rect 208584 7346 208636 7352
rect 208676 5364 208728 5370
rect 208676 5306 208728 5312
rect 207480 3188 207532 3194
rect 207480 3130 207532 3136
rect 208308 3188 208360 3194
rect 208308 3130 208360 3136
rect 207492 400 207520 3130
rect 208688 400 208716 5306
rect 209056 3126 209084 217738
rect 209332 217666 209360 220116
rect 209320 217660 209372 217666
rect 209320 217602 209372 217608
rect 209792 7342 209820 220116
rect 210160 217734 210188 220116
rect 210148 217728 210200 217734
rect 210148 217670 210200 217676
rect 210620 216918 210648 220116
rect 210804 220102 211002 220130
rect 211264 220102 211462 220130
rect 211540 220102 211830 220130
rect 211908 220102 212198 220130
rect 212658 220102 212764 220130
rect 210608 216912 210660 216918
rect 210608 216854 210660 216860
rect 210804 215354 210832 220102
rect 209872 215348 209924 215354
rect 209872 215290 209924 215296
rect 210792 215348 210844 215354
rect 210792 215290 210844 215296
rect 209780 7336 209832 7342
rect 209780 7278 209832 7284
rect 209884 7274 209912 215290
rect 211264 11830 211292 220102
rect 211540 216850 211568 220102
rect 211908 217682 211936 220102
rect 212356 217864 212408 217870
rect 212356 217806 212408 217812
rect 211724 217654 211936 217682
rect 212264 217660 212316 217666
rect 211528 216844 211580 216850
rect 211528 216786 211580 216792
rect 211724 214554 211752 217654
rect 212264 217602 212316 217608
rect 212276 216714 212304 217602
rect 211804 216708 211856 216714
rect 211804 216650 211856 216656
rect 212264 216708 212316 216714
rect 212264 216650 212316 216656
rect 211356 214526 211752 214554
rect 211252 11824 211304 11830
rect 211252 11766 211304 11772
rect 209872 7268 209924 7274
rect 209872 7210 209924 7216
rect 211356 7206 211384 214526
rect 211712 176724 211764 176730
rect 211712 176666 211764 176672
rect 211724 171086 211752 176666
rect 211712 171080 211764 171086
rect 211712 171022 211764 171028
rect 211344 7200 211396 7206
rect 211344 7142 211396 7148
rect 211816 4146 211844 216650
rect 212368 212673 212396 217806
rect 212354 212664 212410 212673
rect 212354 212599 212410 212608
rect 211894 212562 211950 212571
rect 212356 212560 212408 212566
rect 211894 212497 211950 212506
rect 212170 212528 212226 212537
rect 211896 212492 211948 212497
rect 212170 212463 212226 212472
rect 212354 212528 212356 212537
rect 212408 212528 212410 212537
rect 212354 212463 212410 212472
rect 211896 212434 211948 212440
rect 212184 202910 212212 212463
rect 211988 202904 212040 202910
rect 211988 202846 212040 202852
rect 212172 202904 212224 202910
rect 212172 202846 212224 202852
rect 212448 202904 212500 202910
rect 212448 202846 212500 202852
rect 212000 195786 212028 202846
rect 211908 195758 212028 195786
rect 211908 182186 211936 195758
rect 211908 182158 212028 182186
rect 212000 176730 212028 182158
rect 211988 176724 212040 176730
rect 211988 176666 212040 176672
rect 212460 164218 212488 202846
rect 212448 164212 212500 164218
rect 212448 164154 212500 164160
rect 211896 154624 211948 154630
rect 211896 154566 211948 154572
rect 212448 154624 212500 154630
rect 212448 154566 212500 154572
rect 211908 147694 211936 154566
rect 212460 149682 212488 154566
rect 212368 149654 212488 149682
rect 211896 147688 211948 147694
rect 211896 147630 211948 147636
rect 211988 147620 212040 147626
rect 211988 147562 212040 147568
rect 212000 144906 212028 147562
rect 211988 144900 212040 144906
rect 211988 144842 212040 144848
rect 212368 140758 212396 149654
rect 212356 140752 212408 140758
rect 212356 140694 212408 140700
rect 211896 135312 211948 135318
rect 211896 135254 211948 135260
rect 211908 128382 211936 135254
rect 212356 131164 212408 131170
rect 212356 131106 212408 131112
rect 211896 128376 211948 128382
rect 211896 128318 211948 128324
rect 211988 128308 212040 128314
rect 211988 128250 212040 128256
rect 212000 125594 212028 128250
rect 211988 125588 212040 125594
rect 211988 125530 212040 125536
rect 212368 121446 212396 131106
rect 212356 121440 212408 121446
rect 212356 121382 212408 121388
rect 211896 116000 211948 116006
rect 211896 115942 211948 115948
rect 211908 109070 211936 115942
rect 212356 113144 212408 113150
rect 212356 113086 212408 113092
rect 211896 109064 211948 109070
rect 211896 109006 211948 109012
rect 211988 108996 212040 109002
rect 211988 108938 212040 108944
rect 212000 106282 212028 108938
rect 212368 108338 212396 113086
rect 212276 108310 212396 108338
rect 211988 106276 212040 106282
rect 211988 106218 212040 106224
rect 211988 100088 212040 100094
rect 211988 100030 212040 100036
rect 212000 86970 212028 100030
rect 212276 90386 212304 108310
rect 212276 90358 212488 90386
rect 211896 86964 211948 86970
rect 211896 86906 211948 86912
rect 211988 86964 212040 86970
rect 211988 86906 212040 86912
rect 211908 70514 211936 86906
rect 212460 85542 212488 90358
rect 212264 85536 212316 85542
rect 212264 85478 212316 85484
rect 212448 85536 212500 85542
rect 212448 85478 212500 85484
rect 211896 70508 211948 70514
rect 211896 70450 211948 70456
rect 211896 70372 211948 70378
rect 211896 70314 211948 70320
rect 211908 58177 211936 70314
rect 212276 66230 212304 85478
rect 212264 66224 212316 66230
rect 212264 66166 212316 66172
rect 212356 66224 212408 66230
rect 212356 66166 212408 66172
rect 211894 58168 211950 58177
rect 211894 58103 211950 58112
rect 211986 57896 212042 57905
rect 211986 57831 212042 57840
rect 212000 48278 212028 57831
rect 212368 48362 212396 66166
rect 212368 48334 212488 48362
rect 212460 48278 212488 48334
rect 211896 48272 211948 48278
rect 211896 48214 211948 48220
rect 211988 48272 212040 48278
rect 211988 48214 212040 48220
rect 212448 48272 212500 48278
rect 212448 48214 212500 48220
rect 211908 38622 211936 48214
rect 212448 40112 212500 40118
rect 212446 40080 212448 40089
rect 212500 40080 212502 40089
rect 212446 40015 212502 40024
rect 211896 38616 211948 38622
rect 211896 38558 211948 38564
rect 211988 38616 212040 38622
rect 211988 38558 212040 38564
rect 212000 33674 212028 38558
rect 212356 37324 212408 37330
rect 212356 37266 212408 37272
rect 212000 33646 212120 33674
rect 212092 27606 212120 33646
rect 212368 27690 212396 37266
rect 212276 27662 212396 27690
rect 212276 27606 212304 27662
rect 212080 27600 212132 27606
rect 212080 27542 212132 27548
rect 212172 27600 212224 27606
rect 212172 27542 212224 27548
rect 212264 27600 212316 27606
rect 212264 27542 212316 27548
rect 212184 12442 212212 27542
rect 212264 19304 212316 19310
rect 212264 19246 212316 19252
rect 212276 12578 212304 19246
rect 212264 12572 212316 12578
rect 212264 12514 212316 12520
rect 211896 12436 211948 12442
rect 211896 12378 211948 12384
rect 212172 12436 212224 12442
rect 212172 12378 212224 12384
rect 211068 4140 211120 4146
rect 211068 4082 211120 4088
rect 211804 4140 211856 4146
rect 211804 4082 211856 4088
rect 209872 3256 209924 3262
rect 209872 3198 209924 3204
rect 209044 3120 209096 3126
rect 209044 3062 209096 3068
rect 209884 400 209912 3198
rect 211080 400 211108 4082
rect 211908 4078 211936 12378
rect 212736 11898 212764 220102
rect 213012 217938 213040 220116
rect 213196 220102 213486 220130
rect 213564 220102 213854 220130
rect 213932 220102 214314 220130
rect 214484 220102 214682 220130
rect 214760 220102 215142 220130
rect 215312 220102 215510 220130
rect 215588 220102 215878 220130
rect 216048 220102 216338 220130
rect 216706 220102 216812 220130
rect 213000 217932 213052 217938
rect 213000 217874 213052 217880
rect 212816 214600 212868 214606
rect 213196 214554 213224 220102
rect 213564 214606 213592 220102
rect 212816 214542 212868 214548
rect 212724 11892 212776 11898
rect 212724 11834 212776 11840
rect 212264 9716 212316 9722
rect 212264 9658 212316 9664
rect 211896 4072 211948 4078
rect 211896 4014 211948 4020
rect 212276 400 212304 9658
rect 212828 4690 212856 214542
rect 212920 214526 213224 214554
rect 213552 214600 213604 214606
rect 213552 214542 213604 214548
rect 212920 9246 212948 214526
rect 212908 9240 212960 9246
rect 212908 9182 212960 9188
rect 213932 6866 213960 220102
rect 214484 217682 214512 220102
rect 214116 217654 214512 217682
rect 214012 214600 214064 214606
rect 214012 214542 214064 214548
rect 214024 9450 214052 214542
rect 214116 22098 214144 217654
rect 214760 214606 214788 220102
rect 215208 217932 215260 217938
rect 215208 217874 215260 217880
rect 214748 214600 214800 214606
rect 214748 214542 214800 214548
rect 214104 22092 214156 22098
rect 214104 22034 214156 22040
rect 214288 22092 214340 22098
rect 214288 22034 214340 22040
rect 214300 19310 214328 22034
rect 214288 19304 214340 19310
rect 214288 19246 214340 19252
rect 214288 9716 214340 9722
rect 214288 9658 214340 9664
rect 214012 9444 214064 9450
rect 214012 9386 214064 9392
rect 214300 9314 214328 9658
rect 214288 9308 214340 9314
rect 214288 9250 214340 9256
rect 213920 6860 213972 6866
rect 213920 6802 213972 6808
rect 212816 4684 212868 4690
rect 212816 4626 212868 4632
rect 215220 4146 215248 217874
rect 215312 6118 215340 220102
rect 215392 210452 215444 210458
rect 215392 210394 215444 210400
rect 215404 9518 215432 210394
rect 215392 9512 215444 9518
rect 215392 9454 215444 9460
rect 215588 9382 215616 220102
rect 216048 210458 216076 220102
rect 216036 210452 216088 210458
rect 216036 210394 216088 210400
rect 216678 202872 216734 202881
rect 216678 202807 216734 202816
rect 216692 193254 216720 202807
rect 216680 193248 216732 193254
rect 216680 193190 216732 193196
rect 216678 183560 216734 183569
rect 216678 183495 216734 183504
rect 216692 173942 216720 183495
rect 216680 173936 216732 173942
rect 216680 173878 216732 173884
rect 215576 9376 215628 9382
rect 215576 9318 215628 9324
rect 215300 6112 215352 6118
rect 215300 6054 215352 6060
rect 216784 6050 216812 220102
rect 216864 215620 216916 215626
rect 216864 215562 216916 215568
rect 216876 9586 216904 215562
rect 217152 215354 217180 220116
rect 217520 215626 217548 220116
rect 217508 215620 217560 215626
rect 217508 215562 217560 215568
rect 217140 215348 217192 215354
rect 217140 215290 217192 215296
rect 216956 212560 217008 212566
rect 216956 212502 217008 212508
rect 216968 202881 216996 212502
rect 217980 211177 218008 220116
rect 218164 220102 218362 220130
rect 218440 220102 218730 220130
rect 218808 220102 219190 220130
rect 219452 220102 219558 220130
rect 219636 220102 220018 220130
rect 217046 211168 217102 211177
rect 217046 211103 217048 211112
rect 217100 211103 217102 211112
rect 217966 211168 218022 211177
rect 217966 211103 218022 211112
rect 217048 211074 217100 211080
rect 218060 210452 218112 210458
rect 218060 210394 218112 210400
rect 216954 202872 217010 202881
rect 216954 202807 217010 202816
rect 217140 201544 217192 201550
rect 217140 201486 217192 201492
rect 216956 193248 217008 193254
rect 216956 193190 217008 193196
rect 216968 183569 216996 193190
rect 217152 193186 217180 201486
rect 217140 193180 217192 193186
rect 217140 193122 217192 193128
rect 217232 193180 217284 193186
rect 217232 193122 217284 193128
rect 217244 186946 217272 193122
rect 217244 186918 217456 186946
rect 216954 183560 217010 183569
rect 216954 183495 217010 183504
rect 217428 182186 217456 186918
rect 217336 182158 217456 182186
rect 217336 180810 217364 182158
rect 217324 180804 217376 180810
rect 217324 180746 217376 180752
rect 216956 173936 217008 173942
rect 216956 173878 217008 173884
rect 216968 9654 216996 173878
rect 217416 171148 217468 171154
rect 217416 171090 217468 171096
rect 217428 164286 217456 171090
rect 217232 164280 217284 164286
rect 217232 164222 217284 164228
rect 217416 164280 217468 164286
rect 217416 164222 217468 164228
rect 217244 161430 217272 164222
rect 217232 161424 217284 161430
rect 217232 161366 217284 161372
rect 217140 151836 217192 151842
rect 217140 151778 217192 151784
rect 217152 147694 217180 151778
rect 217140 147688 217192 147694
rect 217140 147630 217192 147636
rect 217232 147620 217284 147626
rect 217232 147562 217284 147568
rect 217244 133958 217272 147562
rect 217140 133952 217192 133958
rect 217140 133894 217192 133900
rect 217232 133952 217284 133958
rect 217232 133894 217284 133900
rect 217152 124250 217180 133894
rect 217152 124222 217272 124250
rect 217244 111858 217272 124222
rect 217048 111852 217100 111858
rect 217048 111794 217100 111800
rect 217232 111852 217284 111858
rect 217232 111794 217284 111800
rect 217060 111722 217088 111794
rect 217048 111716 217100 111722
rect 217048 111658 217100 111664
rect 217232 102196 217284 102202
rect 217232 102138 217284 102144
rect 217244 95402 217272 102138
rect 217232 95396 217284 95402
rect 217232 95338 217284 95344
rect 217232 84244 217284 84250
rect 217232 84186 217284 84192
rect 217244 80186 217272 84186
rect 217244 80158 217364 80186
rect 217336 75954 217364 80158
rect 217140 75948 217192 75954
rect 217140 75890 217192 75896
rect 217324 75948 217376 75954
rect 217324 75890 217376 75896
rect 217152 75818 217180 75890
rect 217140 75812 217192 75818
rect 217140 75754 217192 75760
rect 217232 66292 217284 66298
rect 217232 66234 217284 66240
rect 217244 56658 217272 66234
rect 217152 56630 217272 56658
rect 217152 51762 217180 56630
rect 217152 51734 217272 51762
rect 217244 37330 217272 51734
rect 217140 37324 217192 37330
rect 217140 37266 217192 37272
rect 217232 37324 217284 37330
rect 217232 37266 217284 37272
rect 217152 22166 217180 37266
rect 217140 22160 217192 22166
rect 217140 22102 217192 22108
rect 217140 22024 217192 22030
rect 217140 21966 217192 21972
rect 216956 9648 217008 9654
rect 216956 9590 217008 9596
rect 216864 9580 216916 9586
rect 216864 9522 216916 9528
rect 216772 6044 216824 6050
rect 216772 5986 216824 5992
rect 217152 5982 217180 21966
rect 217140 5976 217192 5982
rect 217140 5918 217192 5924
rect 218072 5914 218100 210394
rect 218164 8906 218192 220102
rect 218440 217682 218468 220102
rect 218704 218000 218756 218006
rect 218704 217942 218756 217948
rect 218256 217654 218468 217682
rect 218152 8900 218204 8906
rect 218152 8842 218204 8848
rect 218256 8838 218284 217654
rect 218244 8832 218296 8838
rect 218244 8774 218296 8780
rect 218060 5908 218112 5914
rect 218060 5850 218112 5856
rect 218716 4146 218744 217942
rect 218808 210458 218836 220102
rect 219348 217252 219400 217258
rect 219348 217194 219400 217200
rect 218796 210452 218848 210458
rect 218796 210394 218848 210400
rect 214656 4140 214708 4146
rect 214656 4082 214708 4088
rect 215208 4140 215260 4146
rect 215208 4082 215260 4088
rect 217048 4140 217100 4146
rect 217048 4082 217100 4088
rect 218704 4140 218756 4146
rect 218704 4082 218756 4088
rect 213460 4004 213512 4010
rect 213460 3946 213512 3952
rect 213472 400 213500 3946
rect 214668 400 214696 4082
rect 215852 4072 215904 4078
rect 215852 4014 215904 4020
rect 215864 400 215892 4014
rect 217060 400 217088 4082
rect 218152 3188 218204 3194
rect 218152 3130 218204 3136
rect 218164 400 218192 3130
rect 219360 400 219388 217194
rect 219452 4622 219480 220102
rect 219530 93800 219586 93809
rect 219530 93735 219586 93744
rect 219544 84250 219572 93735
rect 219532 84244 219584 84250
rect 219532 84186 219584 84192
rect 219636 8770 219664 220102
rect 220372 215762 220400 220116
rect 219808 215756 219860 215762
rect 219808 215698 219860 215704
rect 220360 215756 220412 215762
rect 220360 215698 220412 215704
rect 219820 205698 219848 215698
rect 219808 205692 219860 205698
rect 219808 205634 219860 205640
rect 219808 202904 219860 202910
rect 219808 202846 219860 202852
rect 219820 196042 219848 202846
rect 219808 196036 219860 196042
rect 219808 195978 219860 195984
rect 219716 195968 219768 195974
rect 219716 195910 219768 195916
rect 219728 193225 219756 195910
rect 219714 193216 219770 193225
rect 219714 193151 219770 193160
rect 219990 193216 220046 193225
rect 219990 193151 220046 193160
rect 220004 173942 220032 193151
rect 219808 173936 219860 173942
rect 219808 173878 219860 173884
rect 219992 173936 220044 173942
rect 219992 173878 220044 173884
rect 219820 157434 219848 173878
rect 219728 157406 219848 157434
rect 219728 157298 219756 157406
rect 219728 157270 219848 157298
rect 219820 136354 219848 157270
rect 219820 136326 220032 136354
rect 220004 133929 220032 136326
rect 219806 133920 219862 133929
rect 219806 133855 219862 133864
rect 219990 133920 220046 133929
rect 219990 133855 220046 133864
rect 219820 117994 219848 133855
rect 219820 117966 219940 117994
rect 219912 113150 219940 117966
rect 219900 113144 219952 113150
rect 219900 113086 219952 113092
rect 219808 103624 219860 103630
rect 219808 103566 219860 103572
rect 219820 103494 219848 103566
rect 219808 103488 219860 103494
rect 219808 103430 219860 103436
rect 219716 93900 219768 93906
rect 219716 93842 219768 93848
rect 219728 93809 219756 93842
rect 219714 93800 219770 93809
rect 219714 93735 219770 93744
rect 219808 84244 219860 84250
rect 219808 84186 219860 84192
rect 219820 70514 219848 84186
rect 219808 70508 219860 70514
rect 219808 70450 219860 70456
rect 219716 66292 219768 66298
rect 219716 66234 219768 66240
rect 219728 56642 219756 66234
rect 219716 56636 219768 56642
rect 219716 56578 219768 56584
rect 219808 56636 219860 56642
rect 219808 56578 219860 56584
rect 219820 51354 219848 56578
rect 219728 51326 219848 51354
rect 219728 51082 219756 51326
rect 219728 51054 219848 51082
rect 219820 42498 219848 51054
rect 219808 42492 219860 42498
rect 219808 42434 219860 42440
rect 220726 40216 220782 40225
rect 220726 40151 220782 40160
rect 220740 40118 220768 40151
rect 220728 40112 220780 40118
rect 220728 40054 220780 40060
rect 219992 35964 220044 35970
rect 219992 35906 220044 35912
rect 220004 27674 220032 35906
rect 219808 27668 219860 27674
rect 219808 27610 219860 27616
rect 219992 27668 220044 27674
rect 219992 27610 220044 27616
rect 219820 27554 219848 27610
rect 219728 27526 219848 27554
rect 219728 18086 219756 27526
rect 219716 18080 219768 18086
rect 219716 18022 219768 18028
rect 219808 18012 219860 18018
rect 219808 17954 219860 17960
rect 219624 8764 219676 8770
rect 219624 8706 219676 8712
rect 219820 5846 219848 17954
rect 219808 5840 219860 5846
rect 219808 5782 219860 5788
rect 219440 4616 219492 4622
rect 219440 4558 219492 4564
rect 220832 4554 220860 220116
rect 221108 220102 221214 220130
rect 221384 220102 221674 220130
rect 221752 220102 222042 220130
rect 220912 210520 220964 210526
rect 220912 210462 220964 210468
rect 220820 4548 220872 4554
rect 220820 4490 220872 4496
rect 220924 4486 220952 210462
rect 221004 210452 221056 210458
rect 221004 210394 221056 210400
rect 221016 5778 221044 210394
rect 221108 10062 221136 220102
rect 221384 210458 221412 220102
rect 221752 210526 221780 220102
rect 221740 210520 221792 210526
rect 221740 210462 221792 210468
rect 221372 210452 221424 210458
rect 221372 210394 221424 210400
rect 222292 210452 222344 210458
rect 222292 210394 222344 210400
rect 222200 206508 222252 206514
rect 222200 206450 222252 206456
rect 221096 10056 221148 10062
rect 221096 9998 221148 10004
rect 221004 5772 221056 5778
rect 221004 5714 221056 5720
rect 220912 4480 220964 4486
rect 220912 4422 220964 4428
rect 222212 4418 222240 206450
rect 222304 7138 222332 210394
rect 222396 9994 222424 220116
rect 222488 220102 222870 220130
rect 222948 220102 223238 220130
rect 222488 210458 222516 220102
rect 222476 210452 222528 210458
rect 222476 210394 222528 210400
rect 222948 206514 222976 220102
rect 223764 218136 223816 218142
rect 223764 218078 223816 218084
rect 223580 208548 223632 208554
rect 223580 208490 223632 208496
rect 222936 206508 222988 206514
rect 222936 206450 222988 206456
rect 222384 9988 222436 9994
rect 222384 9930 222436 9936
rect 222292 7132 222344 7138
rect 222292 7074 222344 7080
rect 222200 4412 222252 4418
rect 222200 4354 222252 4360
rect 223592 4350 223620 208490
rect 223776 7070 223804 218078
rect 223868 9926 223896 220238
rect 228284 220238 228574 220266
rect 230598 220238 230796 220266
rect 223960 220102 224066 220130
rect 224144 220102 224526 220130
rect 224604 220102 224894 220130
rect 225064 220102 225262 220130
rect 225524 220102 225722 220130
rect 225800 220102 226090 220130
rect 226444 220102 226550 220130
rect 226628 220102 226918 220130
rect 227088 220102 227378 220130
rect 227746 220102 227852 220130
rect 223960 218142 223988 220102
rect 223948 218136 224000 218142
rect 223948 218078 224000 218084
rect 224040 218000 224092 218006
rect 224040 217942 224092 217948
rect 224052 196058 224080 217942
rect 224144 208554 224172 220102
rect 224604 218006 224632 220102
rect 224592 218000 224644 218006
rect 224592 217942 224644 217948
rect 224960 210452 225012 210458
rect 224960 210394 225012 210400
rect 224132 208548 224184 208554
rect 224132 208490 224184 208496
rect 223960 196030 224080 196058
rect 223960 186386 223988 196030
rect 223948 186380 224000 186386
rect 223948 186322 224000 186328
rect 224040 186244 224092 186250
rect 224040 186186 224092 186192
rect 224052 182170 224080 186186
rect 224040 182164 224092 182170
rect 224040 182106 224092 182112
rect 224040 172576 224092 172582
rect 224040 172518 224092 172524
rect 224052 157978 224080 172518
rect 224052 157950 224264 157978
rect 224236 154442 224264 157950
rect 224144 154414 224264 154442
rect 224144 144974 224172 154414
rect 224040 144968 224092 144974
rect 224040 144910 224092 144916
rect 224132 144968 224184 144974
rect 224132 144910 224184 144916
rect 224052 138394 224080 144910
rect 224052 138366 224264 138394
rect 224236 133929 224264 138366
rect 224038 133920 224094 133929
rect 224038 133855 224094 133864
rect 224222 133920 224278 133929
rect 224222 133855 224278 133864
rect 224052 118810 224080 133855
rect 224052 118782 224172 118810
rect 224144 117994 224172 118782
rect 224052 117966 224172 117994
rect 224052 99550 224080 117966
rect 224040 99544 224092 99550
rect 224040 99486 224092 99492
rect 224132 95260 224184 95266
rect 224132 95202 224184 95208
rect 224144 85610 224172 95202
rect 224040 85604 224092 85610
rect 224040 85546 224092 85552
rect 224132 85604 224184 85610
rect 224132 85546 224184 85552
rect 224052 77382 224080 85546
rect 224040 77376 224092 77382
rect 224040 77318 224092 77324
rect 223948 77240 224000 77246
rect 223948 77182 224000 77188
rect 223960 67590 223988 77182
rect 223948 67584 224000 67590
rect 223948 67526 224000 67532
rect 224040 67516 224092 67522
rect 224040 67458 224092 67464
rect 224052 51134 224080 67458
rect 224040 51128 224092 51134
rect 224040 51070 224092 51076
rect 224040 50992 224092 50998
rect 224040 50934 224092 50940
rect 224052 28914 224080 50934
rect 223960 28886 224080 28914
rect 223960 19378 223988 28886
rect 223948 19372 224000 19378
rect 223948 19314 224000 19320
rect 224040 19372 224092 19378
rect 224040 19314 224092 19320
rect 223856 9920 223908 9926
rect 223856 9862 223908 9868
rect 223764 7064 223816 7070
rect 223764 7006 223816 7012
rect 224052 5710 224080 19314
rect 224040 5704 224092 5710
rect 224040 5646 224092 5652
rect 223580 4344 223632 4350
rect 223580 4286 223632 4292
rect 224972 4282 225000 210394
rect 225064 7002 225092 220102
rect 225524 211154 225552 220102
rect 225432 211126 225552 211154
rect 225432 209778 225460 211126
rect 225800 210458 225828 220102
rect 226248 217184 226300 217190
rect 226248 217126 226300 217132
rect 225788 210452 225840 210458
rect 225788 210394 225840 210400
rect 225144 209772 225196 209778
rect 225144 209714 225196 209720
rect 225420 209772 225472 209778
rect 225420 209714 225472 209720
rect 225156 200161 225184 209714
rect 225142 200152 225198 200161
rect 225142 200087 225198 200096
rect 225326 200152 225382 200161
rect 225326 200087 225382 200096
rect 225340 190482 225368 200087
rect 225340 190466 225460 190482
rect 225236 190460 225288 190466
rect 225340 190460 225472 190466
rect 225340 190454 225420 190460
rect 225236 190402 225288 190408
rect 225420 190402 225472 190408
rect 225248 180849 225276 190402
rect 225432 190371 225460 190402
rect 225234 180840 225290 180849
rect 225234 180775 225290 180784
rect 225510 180840 225566 180849
rect 225510 180775 225566 180784
rect 225524 176882 225552 180775
rect 225432 176854 225552 176882
rect 225432 172514 225460 176854
rect 225420 172508 225472 172514
rect 225420 172450 225472 172456
rect 225420 162716 225472 162722
rect 225420 162658 225472 162664
rect 225432 160070 225460 162658
rect 225420 160064 225472 160070
rect 225420 160006 225472 160012
rect 225604 160064 225656 160070
rect 225604 160006 225656 160012
rect 225616 158710 225644 160006
rect 225604 158704 225656 158710
rect 225604 158646 225656 158652
rect 225604 150340 225656 150346
rect 225604 150282 225656 150288
rect 225616 140826 225644 150282
rect 225236 140820 225288 140826
rect 225236 140762 225288 140768
rect 225604 140820 225656 140826
rect 225604 140762 225656 140768
rect 225248 140706 225276 140762
rect 225326 140720 225382 140729
rect 225248 140678 225326 140706
rect 225326 140655 225382 140664
rect 225510 140720 225566 140729
rect 225510 140655 225566 140664
rect 225524 133822 225552 140655
rect 225328 133816 225380 133822
rect 225328 133758 225380 133764
rect 225512 133816 225564 133822
rect 225512 133758 225564 133764
rect 225340 122806 225368 133758
rect 225236 122800 225288 122806
rect 225236 122742 225288 122748
rect 225328 122800 225380 122806
rect 225328 122742 225380 122748
rect 225248 117858 225276 122742
rect 225248 117830 225368 117858
rect 225340 99686 225368 117830
rect 225328 99680 225380 99686
rect 225328 99622 225380 99628
rect 225328 95260 225380 95266
rect 225328 95202 225380 95208
rect 225340 86970 225368 95202
rect 225236 86964 225288 86970
rect 225236 86906 225288 86912
rect 225328 86964 225380 86970
rect 225328 86906 225380 86912
rect 225248 80730 225276 86906
rect 225248 80702 225460 80730
rect 225432 77194 225460 80702
rect 225340 77166 225460 77194
rect 225340 67658 225368 77166
rect 225236 67652 225288 67658
rect 225236 67594 225288 67600
rect 225328 67652 225380 67658
rect 225328 67594 225380 67600
rect 225248 56574 225276 67594
rect 225236 56568 225288 56574
rect 225236 56510 225288 56516
rect 225512 56568 225564 56574
rect 225512 56510 225564 56516
rect 225524 37330 225552 56510
rect 225236 37324 225288 37330
rect 225236 37266 225288 37272
rect 225512 37324 225564 37330
rect 225512 37266 225564 37272
rect 225248 8634 225276 37266
rect 225236 8628 225288 8634
rect 225236 8570 225288 8576
rect 225052 6996 225104 7002
rect 225052 6938 225104 6944
rect 224960 4276 225012 4282
rect 224960 4218 225012 4224
rect 221740 4140 221792 4146
rect 221740 4082 221792 4088
rect 220544 2916 220596 2922
rect 220544 2858 220596 2864
rect 220556 400 220584 2858
rect 221752 400 221780 4082
rect 226260 3942 226288 217126
rect 226340 210452 226392 210458
rect 226340 210394 226392 210400
rect 226352 4214 226380 210394
rect 226444 5642 226472 220102
rect 226628 8566 226656 220102
rect 227088 210458 227116 220102
rect 227628 217116 227680 217122
rect 227628 217058 227680 217064
rect 227076 210452 227128 210458
rect 227076 210394 227128 210400
rect 226616 8560 226668 8566
rect 226616 8502 226668 8508
rect 226432 5636 226484 5642
rect 226432 5578 226484 5584
rect 226340 4208 226392 4214
rect 226340 4150 226392 4156
rect 225328 3936 225380 3942
rect 225328 3878 225380 3884
rect 226248 3936 226300 3942
rect 226248 3878 226300 3884
rect 224132 3120 224184 3126
rect 224132 3062 224184 3068
rect 222936 3052 222988 3058
rect 222936 2994 222988 3000
rect 222948 400 222976 2994
rect 224144 400 224172 3062
rect 225340 400 225368 3878
rect 227640 3466 227668 217058
rect 227824 5574 227852 220102
rect 228008 220102 228206 220130
rect 227904 210452 227956 210458
rect 227904 210394 227956 210400
rect 227916 6186 227944 210394
rect 228008 8498 228036 220102
rect 228284 182170 228312 220238
rect 228652 220102 228942 220130
rect 228652 210458 228680 220102
rect 229388 212537 229416 220116
rect 229480 220102 229770 220130
rect 229848 220102 230230 220130
rect 229374 212528 229430 212537
rect 229374 212463 229430 212472
rect 229480 210458 229508 220102
rect 229744 216980 229796 216986
rect 229744 216922 229796 216928
rect 229558 212528 229614 212537
rect 229558 212463 229614 212472
rect 228640 210452 228692 210458
rect 228640 210394 228692 210400
rect 229100 210452 229152 210458
rect 229100 210394 229152 210400
rect 229468 210452 229520 210458
rect 229468 210394 229520 210400
rect 228272 182164 228324 182170
rect 228272 182106 228324 182112
rect 228364 182164 228416 182170
rect 228364 182106 228416 182112
rect 228376 158710 228404 182106
rect 228364 158704 228416 158710
rect 228364 158646 228416 158652
rect 228548 158704 228600 158710
rect 228548 158646 228600 158652
rect 228560 157350 228588 158646
rect 228548 157344 228600 157350
rect 228548 157286 228600 157292
rect 228180 139460 228232 139466
rect 228180 139402 228232 139408
rect 228192 139346 228220 139402
rect 228270 139360 228326 139369
rect 228192 139318 228270 139346
rect 228270 139295 228326 139304
rect 228454 139360 228510 139369
rect 228454 139295 228510 139304
rect 228468 133822 228496 139295
rect 228272 133816 228324 133822
rect 228272 133758 228324 133764
rect 228456 133816 228508 133822
rect 228456 133758 228508 133764
rect 228284 122754 228312 133758
rect 228284 122726 228404 122754
rect 228376 110922 228404 122726
rect 228284 110894 228404 110922
rect 228284 99634 228312 110894
rect 228284 99606 228404 99634
rect 228376 99362 228404 99606
rect 228284 99334 228404 99362
rect 228284 86970 228312 99334
rect 228180 86964 228232 86970
rect 228180 86906 228232 86912
rect 228272 86964 228324 86970
rect 228272 86906 228324 86912
rect 228192 85542 228220 86906
rect 228180 85536 228232 85542
rect 228180 85478 228232 85484
rect 228272 85536 228324 85542
rect 228272 85478 228324 85484
rect 228284 75970 228312 85478
rect 228192 75942 228312 75970
rect 228192 55214 228220 75942
rect 228180 55208 228232 55214
rect 228180 55150 228232 55156
rect 228272 46912 228324 46918
rect 228272 46854 228324 46860
rect 228284 45558 228312 46854
rect 228180 45552 228232 45558
rect 228180 45494 228232 45500
rect 228272 45552 228324 45558
rect 228272 45494 228324 45500
rect 228192 17898 228220 45494
rect 228192 17870 228312 17898
rect 228284 8514 228312 17870
rect 227996 8492 228048 8498
rect 227996 8434 228048 8440
rect 228192 8486 228312 8514
rect 227904 6180 227956 6186
rect 227904 6122 227956 6128
rect 227812 5568 227864 5574
rect 227812 5510 227864 5516
rect 228192 4826 228220 8486
rect 229112 4894 229140 210394
rect 229572 210338 229600 212463
rect 229480 210310 229600 210338
rect 229192 207052 229244 207058
rect 229192 206994 229244 207000
rect 229204 6254 229232 206994
rect 229480 200122 229508 210310
rect 229468 200116 229520 200122
rect 229468 200058 229520 200064
rect 229560 200116 229612 200122
rect 229560 200058 229612 200064
rect 229572 182209 229600 200058
rect 229282 182200 229338 182209
rect 229558 182200 229614 182209
rect 229282 182135 229284 182144
rect 229336 182135 229338 182144
rect 229468 182164 229520 182170
rect 229284 182106 229336 182112
rect 229558 182135 229614 182144
rect 229468 182106 229520 182112
rect 229480 176474 229508 182106
rect 229388 176446 229508 176474
rect 229388 172514 229416 176446
rect 229376 172508 229428 172514
rect 229376 172450 229428 172456
rect 229376 164212 229428 164218
rect 229376 164154 229428 164160
rect 229388 162874 229416 164154
rect 229388 162858 229508 162874
rect 229388 162852 229520 162858
rect 229388 162846 229468 162852
rect 229468 162794 229520 162800
rect 229284 153264 229336 153270
rect 229284 153206 229336 153212
rect 229296 142118 229324 153206
rect 229284 142112 229336 142118
rect 229284 142054 229336 142060
rect 229376 142112 229428 142118
rect 229376 142054 229428 142060
rect 229388 125769 229416 142054
rect 229374 125760 229430 125769
rect 229374 125695 229430 125704
rect 229282 125624 229338 125633
rect 229282 125559 229338 125568
rect 229296 122806 229324 125559
rect 229284 122800 229336 122806
rect 229284 122742 229336 122748
rect 229284 118040 229336 118046
rect 229284 117982 229336 117988
rect 229296 100042 229324 117982
rect 229296 100014 229508 100042
rect 229480 99226 229508 100014
rect 229388 99198 229508 99226
rect 229388 91882 229416 99198
rect 229388 91854 229508 91882
rect 229480 87009 229508 91854
rect 229282 87000 229338 87009
rect 229282 86935 229284 86944
rect 229336 86935 229338 86944
rect 229466 87000 229522 87009
rect 229466 86935 229522 86944
rect 229284 86906 229336 86912
rect 229376 86896 229428 86902
rect 229376 86838 229428 86844
rect 229388 77518 229416 86838
rect 229376 77512 229428 77518
rect 229376 77454 229428 77460
rect 229376 77376 229428 77382
rect 229376 77318 229428 77324
rect 229388 77194 229416 77318
rect 229296 77166 229416 77194
rect 229296 67590 229324 77166
rect 229284 67584 229336 67590
rect 229284 67526 229336 67532
rect 229376 67516 229428 67522
rect 229376 67458 229428 67464
rect 229388 51134 229416 67458
rect 229376 51128 229428 51134
rect 229376 51070 229428 51076
rect 229376 50992 229428 50998
rect 229376 50934 229428 50940
rect 229388 38622 229416 50934
rect 229284 38616 229336 38622
rect 229284 38558 229336 38564
rect 229376 38616 229428 38622
rect 229376 38558 229428 38564
rect 229296 19378 229324 38558
rect 229284 19372 229336 19378
rect 229284 19314 229336 19320
rect 229376 19372 229428 19378
rect 229376 19314 229428 19320
rect 229388 8430 229416 19314
rect 229376 8424 229428 8430
rect 229376 8366 229428 8372
rect 229192 6248 229244 6254
rect 229192 6190 229244 6196
rect 229100 4888 229152 4894
rect 229100 4830 229152 4836
rect 228180 4820 228232 4826
rect 228180 4762 228232 4768
rect 226524 3460 226576 3466
rect 226524 3402 226576 3408
rect 227628 3460 227680 3466
rect 227628 3402 227680 3408
rect 226536 400 226564 3402
rect 228916 3188 228968 3194
rect 228916 3130 228968 3136
rect 227720 2848 227772 2854
rect 227720 2790 227772 2796
rect 227732 400 227760 2790
rect 228928 400 228956 3130
rect 229756 3058 229784 216922
rect 229848 207058 229876 220102
rect 230388 217048 230440 217054
rect 230388 216990 230440 216996
rect 229836 207052 229888 207058
rect 229836 206994 229888 207000
rect 229744 3052 229796 3058
rect 229744 2994 229796 3000
rect 230400 490 230428 216990
rect 230480 210452 230532 210458
rect 230480 210394 230532 210400
rect 230492 6322 230520 210394
rect 230664 205896 230716 205902
rect 230664 205838 230716 205844
rect 230572 191140 230624 191146
rect 230572 191082 230624 191088
rect 230584 181490 230612 191082
rect 230572 181484 230624 181490
rect 230572 181426 230624 181432
rect 230572 152108 230624 152114
rect 230572 152050 230624 152056
rect 230584 142866 230612 152050
rect 230572 142860 230624 142866
rect 230572 142802 230624 142808
rect 230572 16788 230624 16794
rect 230572 16730 230624 16736
rect 230584 8974 230612 16730
rect 230676 9042 230704 205838
rect 230768 191146 230796 220238
rect 235552 220238 235934 220266
rect 276690 220238 277072 220266
rect 230860 220102 231058 220130
rect 231136 220102 231426 220130
rect 231688 220102 231794 220130
rect 231964 220102 232254 220130
rect 232332 220102 232622 220130
rect 232792 220102 233082 220130
rect 233252 220102 233450 220130
rect 233528 220102 233910 220130
rect 233988 220102 234278 220130
rect 234738 220102 234844 220130
rect 230860 205902 230888 220102
rect 231136 210458 231164 220102
rect 231688 215234 231716 220102
rect 231412 215206 231716 215234
rect 231124 210452 231176 210458
rect 231124 210394 231176 210400
rect 230848 205896 230900 205902
rect 230848 205838 230900 205844
rect 231412 200122 231440 215206
rect 231860 210452 231912 210458
rect 231860 210394 231912 210400
rect 230848 200116 230900 200122
rect 230848 200058 230900 200064
rect 231400 200116 231452 200122
rect 231400 200058 231452 200064
rect 230756 191140 230808 191146
rect 230756 191082 230808 191088
rect 230860 190505 230888 200058
rect 230846 190496 230902 190505
rect 230846 190431 230902 190440
rect 231030 190496 231086 190505
rect 231030 190431 231086 190440
rect 231044 186454 231072 190431
rect 231032 186448 231084 186454
rect 231032 186390 231084 186396
rect 230940 186312 230992 186318
rect 230940 186254 230992 186260
rect 230952 182170 230980 186254
rect 230940 182164 230992 182170
rect 230940 182106 230992 182112
rect 231032 182164 231084 182170
rect 231032 182106 231084 182112
rect 230756 181484 230808 181490
rect 230756 181426 230808 181432
rect 230768 171850 230796 181426
rect 230768 171822 230980 171850
rect 230952 162330 230980 171822
rect 231044 169130 231072 182106
rect 231044 169102 231256 169130
rect 230768 162302 230980 162330
rect 230768 152114 230796 162302
rect 231228 154601 231256 169102
rect 230938 154592 230994 154601
rect 230938 154527 230994 154536
rect 231214 154592 231270 154601
rect 231214 154527 231270 154536
rect 230952 153202 230980 154527
rect 230940 153196 230992 153202
rect 230940 153138 230992 153144
rect 231768 153196 231820 153202
rect 231768 153138 231820 153144
rect 230756 152108 230808 152114
rect 230756 152050 230808 152056
rect 230940 144900 230992 144906
rect 230940 144842 230992 144848
rect 230952 143562 230980 144842
rect 231780 143585 231808 153138
rect 231766 143576 231822 143585
rect 230952 143534 231072 143562
rect 230756 142860 230808 142866
rect 230756 142802 230808 142808
rect 230768 133226 230796 142802
rect 231044 135250 231072 143534
rect 231766 143511 231822 143520
rect 231032 135244 231084 135250
rect 231032 135186 231084 135192
rect 231216 135244 231268 135250
rect 231216 135186 231268 135192
rect 230768 133198 230980 133226
rect 230952 123570 230980 133198
rect 231228 129010 231256 135186
rect 231136 128982 231256 129010
rect 231136 124166 231164 128982
rect 231124 124160 231176 124166
rect 231124 124102 231176 124108
rect 230768 123542 230980 123570
rect 230768 113898 230796 123542
rect 231032 114572 231084 114578
rect 231032 114514 231084 114520
rect 230756 113892 230808 113898
rect 230756 113834 230808 113840
rect 230940 113892 230992 113898
rect 230940 113834 230992 113840
rect 230756 111104 230808 111110
rect 230756 111046 230808 111052
rect 230768 104394 230796 111046
rect 230768 104366 230888 104394
rect 230756 104236 230808 104242
rect 230756 104178 230808 104184
rect 230768 94586 230796 104178
rect 230756 94580 230808 94586
rect 230756 94522 230808 94528
rect 230860 94466 230888 104366
rect 230952 104242 230980 113834
rect 231044 111110 231072 114514
rect 231032 111104 231084 111110
rect 231032 111046 231084 111052
rect 230940 104236 230992 104242
rect 230940 104178 230992 104184
rect 230940 94580 230992 94586
rect 230940 94522 230992 94528
rect 230768 94438 230888 94466
rect 230768 85082 230796 94438
rect 230768 85054 230888 85082
rect 230756 84924 230808 84930
rect 230756 84866 230808 84872
rect 230768 75274 230796 84866
rect 230756 75268 230808 75274
rect 230756 75210 230808 75216
rect 230860 75154 230888 85054
rect 230952 84930 230980 94522
rect 230940 84924 230992 84930
rect 230940 84866 230992 84872
rect 230940 75268 230992 75274
rect 230940 75210 230992 75216
rect 230768 75126 230888 75154
rect 230768 65958 230796 75126
rect 230756 65952 230808 65958
rect 230756 65894 230808 65900
rect 230952 61010 230980 75210
rect 230768 60982 230980 61010
rect 230768 55842 230796 60982
rect 231032 56636 231084 56642
rect 231032 56578 231084 56584
rect 231044 56506 231072 56578
rect 231032 56500 231084 56506
rect 231032 56442 231084 56448
rect 231400 56500 231452 56506
rect 231400 56442 231452 56448
rect 230768 55814 230980 55842
rect 230952 38690 230980 55814
rect 231412 47002 231440 56442
rect 231228 46974 231440 47002
rect 231228 45558 231256 46974
rect 231216 45552 231268 45558
rect 231216 45494 231268 45500
rect 231308 45552 231360 45558
rect 231308 45494 231360 45500
rect 230756 38684 230808 38690
rect 230756 38626 230808 38632
rect 230940 38684 230992 38690
rect 230940 38626 230992 38632
rect 230768 36530 230796 38626
rect 230768 36502 230980 36530
rect 230952 26874 230980 36502
rect 231320 29102 231348 45494
rect 231308 29096 231360 29102
rect 231308 29038 231360 29044
rect 231124 28960 231176 28966
rect 231124 28902 231176 28908
rect 230768 26846 230980 26874
rect 230768 16794 230796 26846
rect 231136 26654 231164 28902
rect 230940 26648 230992 26654
rect 230940 26590 230992 26596
rect 231124 26648 231176 26654
rect 231124 26590 231176 26596
rect 230756 16788 230808 16794
rect 230756 16730 230808 16736
rect 230952 9110 230980 26590
rect 230940 9104 230992 9110
rect 230940 9046 230992 9052
rect 230664 9036 230716 9042
rect 230664 8978 230716 8984
rect 230572 8968 230624 8974
rect 230572 8910 230624 8916
rect 230480 6316 230532 6322
rect 230480 6258 230532 6264
rect 231872 3602 231900 210394
rect 231860 3596 231912 3602
rect 231860 3538 231912 3544
rect 231964 3398 231992 220102
rect 232332 216322 232360 220102
rect 232504 216844 232556 216850
rect 232504 216786 232556 216792
rect 232056 216294 232360 216322
rect 232056 212537 232084 216294
rect 232042 212528 232098 212537
rect 232042 212463 232098 212472
rect 232318 212528 232374 212537
rect 232318 212463 232374 212472
rect 232332 202910 232360 212463
rect 232136 202904 232188 202910
rect 232136 202846 232188 202852
rect 232320 202904 232372 202910
rect 232320 202846 232372 202852
rect 232148 198150 232176 202846
rect 232136 198144 232188 198150
rect 232136 198086 232188 198092
rect 232044 198076 232096 198082
rect 232044 198018 232096 198024
rect 232056 193225 232084 198018
rect 232042 193216 232098 193225
rect 232042 193151 232098 193160
rect 232226 193216 232282 193225
rect 232226 193151 232282 193160
rect 232148 183598 232176 183629
rect 232240 183598 232268 193151
rect 232136 183592 232188 183598
rect 232228 183592 232280 183598
rect 232188 183540 232228 183546
rect 232136 183534 232280 183540
rect 232148 183518 232268 183534
rect 232240 174010 232268 183518
rect 232136 174004 232188 174010
rect 232136 173946 232188 173952
rect 232228 174004 232280 174010
rect 232228 173946 232280 173952
rect 232148 167142 232176 173946
rect 232136 167136 232188 167142
rect 232136 167078 232188 167084
rect 232136 167000 232188 167006
rect 232136 166942 232188 166948
rect 232148 157282 232176 166942
rect 232136 157276 232188 157282
rect 232136 157218 232188 157224
rect 232044 157140 232096 157146
rect 232044 157082 232096 157088
rect 232056 153202 232084 157082
rect 232044 153196 232096 153202
rect 232044 153138 232096 153144
rect 232042 143576 232098 143585
rect 232042 143511 232098 143520
rect 232056 139262 232084 143511
rect 232044 139256 232096 139262
rect 232044 139198 232096 139204
rect 232320 139256 232372 139262
rect 232320 139198 232372 139204
rect 232332 124234 232360 139198
rect 232228 124228 232280 124234
rect 232228 124170 232280 124176
rect 232320 124228 232372 124234
rect 232320 124170 232372 124176
rect 232240 124114 232268 124170
rect 232240 124086 232360 124114
rect 232332 122806 232360 124086
rect 232320 122800 232372 122806
rect 232320 122742 232372 122748
rect 232228 113212 232280 113218
rect 232228 113154 232280 113160
rect 232240 99226 232268 113154
rect 232056 99198 232268 99226
rect 232056 96626 232084 99198
rect 232044 96620 232096 96626
rect 232044 96562 232096 96568
rect 232228 96620 232280 96626
rect 232228 96562 232280 96568
rect 232240 77314 232268 96562
rect 232228 77308 232280 77314
rect 232228 77250 232280 77256
rect 232228 75948 232280 75954
rect 232228 75890 232280 75896
rect 232240 67658 232268 75890
rect 232044 67652 232096 67658
rect 232044 67594 232096 67600
rect 232228 67652 232280 67658
rect 232228 67594 232280 67600
rect 232056 61418 232084 67594
rect 232056 61390 232268 61418
rect 232240 60704 232268 61390
rect 232148 60676 232268 60704
rect 232148 51134 232176 60676
rect 232136 51128 232188 51134
rect 232136 51070 232188 51076
rect 232044 51060 232096 51066
rect 232044 51002 232096 51008
rect 232056 46918 232084 51002
rect 232044 46912 232096 46918
rect 232044 46854 232096 46860
rect 232044 37324 232096 37330
rect 232044 37266 232096 37272
rect 232056 29034 232084 37266
rect 232044 29028 232096 29034
rect 232044 28970 232096 28976
rect 232136 29028 232188 29034
rect 232136 28970 232188 28976
rect 232148 6390 232176 28970
rect 232136 6384 232188 6390
rect 232136 6326 232188 6332
rect 232516 3618 232544 216786
rect 232792 210458 232820 220102
rect 232780 210452 232832 210458
rect 232780 210394 232832 210400
rect 233252 3942 233280 220102
rect 233332 210452 233384 210458
rect 233332 210394 233384 210400
rect 233344 4962 233372 210394
rect 233528 6458 233556 220102
rect 233988 210458 234016 220102
rect 233976 210452 234028 210458
rect 233976 210394 234028 210400
rect 234620 210384 234672 210390
rect 234620 210326 234672 210332
rect 233516 6452 233568 6458
rect 233516 6394 233568 6400
rect 233332 4956 233384 4962
rect 233332 4898 233384 4904
rect 233240 3936 233292 3942
rect 233240 3878 233292 3884
rect 233700 3936 233752 3942
rect 233700 3878 233752 3884
rect 232424 3590 232544 3618
rect 232424 3466 232452 3590
rect 232412 3460 232464 3466
rect 232412 3402 232464 3408
rect 232504 3460 232556 3466
rect 232504 3402 232556 3408
rect 231952 3392 232004 3398
rect 231952 3334 232004 3340
rect 231308 3052 231360 3058
rect 231308 2994 231360 3000
rect 230124 462 230428 490
rect 230124 400 230152 462
rect 231320 400 231348 2994
rect 232516 400 232544 3402
rect 233712 400 233740 3878
rect 234632 3738 234660 210326
rect 234816 205766 234844 220102
rect 234908 220102 235106 220130
rect 235276 220102 235474 220130
rect 234908 210390 234936 220102
rect 235276 217682 235304 220102
rect 235092 217654 235304 217682
rect 234896 210384 234948 210390
rect 234896 210326 234948 210332
rect 235092 210202 235120 217654
rect 235552 212514 235580 220238
rect 236104 220102 236302 220130
rect 235552 212486 235672 212514
rect 234908 210174 235120 210202
rect 234804 205760 234856 205766
rect 234804 205702 234856 205708
rect 234804 205624 234856 205630
rect 234804 205566 234856 205572
rect 234816 198014 234844 205566
rect 234804 198008 234856 198014
rect 234804 197950 234856 197956
rect 234804 41472 234856 41478
rect 234804 41414 234856 41420
rect 234816 31822 234844 41414
rect 234804 31816 234856 31822
rect 234804 31758 234856 31764
rect 234712 31748 234764 31754
rect 234712 31690 234764 31696
rect 234724 25158 234752 31690
rect 234712 25152 234764 25158
rect 234712 25094 234764 25100
rect 234712 12504 234764 12510
rect 234712 12446 234764 12452
rect 234620 3732 234672 3738
rect 234620 3674 234672 3680
rect 234724 3670 234752 12446
rect 234908 5030 234936 210174
rect 235644 198082 235672 212486
rect 236000 210452 236052 210458
rect 236000 210394 236052 210400
rect 234988 198076 235040 198082
rect 234988 198018 235040 198024
rect 235632 198076 235684 198082
rect 235632 198018 235684 198024
rect 235000 183598 235028 198018
rect 235172 198008 235224 198014
rect 235172 197950 235224 197956
rect 234988 183592 235040 183598
rect 235080 183592 235132 183598
rect 234988 183534 235040 183540
rect 235078 183560 235080 183569
rect 235132 183560 235134 183569
rect 235078 183495 235134 183504
rect 235184 164393 235212 197950
rect 235354 183560 235410 183569
rect 235354 183495 235410 183504
rect 235170 164384 235226 164393
rect 235170 164319 235226 164328
rect 235368 164286 235396 183495
rect 235264 164280 235316 164286
rect 235078 164248 235134 164257
rect 235264 164222 235316 164228
rect 235356 164280 235408 164286
rect 235356 164222 235408 164228
rect 235078 164183 235080 164192
rect 235132 164183 235134 164192
rect 235080 164154 235132 164160
rect 235172 164144 235224 164150
rect 235172 164086 235224 164092
rect 235184 154562 235212 164086
rect 234988 154556 235040 154562
rect 234988 154498 235040 154504
rect 235172 154556 235224 154562
rect 235172 154498 235224 154504
rect 235000 145058 235028 154498
rect 235000 145030 235120 145058
rect 234988 142860 235040 142866
rect 234988 142802 235040 142808
rect 235000 138009 235028 142802
rect 235092 142118 235120 145030
rect 235276 142866 235304 164222
rect 235264 142860 235316 142866
rect 235264 142802 235316 142808
rect 235080 142112 235132 142118
rect 235080 142054 235132 142060
rect 235172 142044 235224 142050
rect 235172 141986 235224 141992
rect 234986 138000 235042 138009
rect 234986 137935 235042 137944
rect 235184 125769 235212 141986
rect 235262 138000 235318 138009
rect 235262 137935 235318 137944
rect 235170 125760 235226 125769
rect 235170 125695 235226 125704
rect 235078 125624 235134 125633
rect 235078 125559 235080 125568
rect 235132 125559 235134 125568
rect 235080 125530 235132 125536
rect 235172 125520 235224 125526
rect 235172 125462 235224 125468
rect 235184 106457 235212 125462
rect 235276 118726 235304 137935
rect 235264 118720 235316 118726
rect 235264 118662 235316 118668
rect 235264 116000 235316 116006
rect 235264 115942 235316 115948
rect 235170 106448 235226 106457
rect 235170 106383 235226 106392
rect 235078 106312 235134 106321
rect 235078 106247 235080 106256
rect 235132 106247 235134 106256
rect 235080 106218 235132 106224
rect 235172 106208 235224 106214
rect 235172 106150 235224 106156
rect 235184 96626 235212 106150
rect 235276 99414 235304 115942
rect 235264 99408 235316 99414
rect 235264 99350 235316 99356
rect 235264 96688 235316 96694
rect 235264 96630 235316 96636
rect 235172 96620 235224 96626
rect 235172 96562 235224 96568
rect 235078 87000 235134 87009
rect 235078 86935 235080 86944
rect 235132 86935 235134 86944
rect 235080 86906 235132 86912
rect 235172 86896 235224 86902
rect 235172 86838 235224 86844
rect 235184 67726 235212 86838
rect 235276 80102 235304 96630
rect 235356 96620 235408 96626
rect 235356 96562 235408 96568
rect 235368 87009 235396 96562
rect 235354 87000 235410 87009
rect 235354 86935 235410 86944
rect 235264 80096 235316 80102
rect 235264 80038 235316 80044
rect 235264 77308 235316 77314
rect 235264 77250 235316 77256
rect 235172 67720 235224 67726
rect 235172 67662 235224 67668
rect 235080 67652 235132 67658
rect 235080 67594 235132 67600
rect 235092 66230 235120 67594
rect 235080 66224 235132 66230
rect 235080 66166 235132 66172
rect 235172 66156 235224 66162
rect 235172 66098 235224 66104
rect 234988 65544 235040 65550
rect 234988 65486 235040 65492
rect 235000 60654 235028 65486
rect 234988 60648 235040 60654
rect 234988 60590 235040 60596
rect 235184 48414 235212 66098
rect 235276 65550 235304 77250
rect 235264 65544 235316 65550
rect 235264 65486 235316 65492
rect 235264 60648 235316 60654
rect 235264 60590 235316 60596
rect 235276 51134 235304 60590
rect 235264 51128 235316 51134
rect 235264 51070 235316 51076
rect 235356 51060 235408 51066
rect 235356 51002 235408 51008
rect 235172 48408 235224 48414
rect 235172 48350 235224 48356
rect 235080 48340 235132 48346
rect 235080 48282 235132 48288
rect 235092 41478 235120 48282
rect 235080 41472 235132 41478
rect 234986 41440 235042 41449
rect 235368 41449 235396 51002
rect 235080 41414 235132 41420
rect 235354 41440 235410 41449
rect 234986 41375 235042 41384
rect 235354 41375 235410 41384
rect 235000 41290 235028 41375
rect 235000 41262 235120 41290
rect 235092 38622 235120 41262
rect 235080 38616 235132 38622
rect 235080 38558 235132 38564
rect 235264 38616 235316 38622
rect 235264 38558 235316 38564
rect 235172 25152 235224 25158
rect 235172 25094 235224 25100
rect 235184 12510 235212 25094
rect 235172 12504 235224 12510
rect 235172 12446 235224 12452
rect 234896 5024 234948 5030
rect 234896 4966 234948 4972
rect 234804 4004 234856 4010
rect 234804 3946 234856 3952
rect 234712 3664 234764 3670
rect 234712 3606 234764 3612
rect 234816 400 234844 3946
rect 235276 3874 235304 38558
rect 235264 3868 235316 3874
rect 235264 3810 235316 3816
rect 236012 3806 236040 210394
rect 236000 3800 236052 3806
rect 236000 3742 236052 3748
rect 236104 3602 236132 220102
rect 236748 212566 236776 220116
rect 236840 220102 237130 220130
rect 236276 212560 236328 212566
rect 236276 212502 236328 212508
rect 236736 212560 236788 212566
rect 236736 212502 236788 212508
rect 236288 205630 236316 212502
rect 236840 210458 236868 220102
rect 237576 217530 237604 220116
rect 237668 220102 237958 220130
rect 237564 217524 237616 217530
rect 237564 217466 237616 217472
rect 237288 216912 237340 216918
rect 237288 216854 237340 216860
rect 236828 210452 236880 210458
rect 236828 210394 236880 210400
rect 236276 205624 236328 205630
rect 236276 205566 236328 205572
rect 236460 205624 236512 205630
rect 236460 205566 236512 205572
rect 236472 197826 236500 205566
rect 236380 197798 236500 197826
rect 236380 186266 236408 197798
rect 236288 186238 236408 186266
rect 236288 182170 236316 186238
rect 236276 182164 236328 182170
rect 236276 182106 236328 182112
rect 236460 182164 236512 182170
rect 236460 182106 236512 182112
rect 236472 172530 236500 182106
rect 236380 172502 236500 172530
rect 236380 171086 236408 172502
rect 236368 171080 236420 171086
rect 236368 171022 236420 171028
rect 236276 160132 236328 160138
rect 236276 160074 236328 160080
rect 236288 142254 236316 160074
rect 236184 142248 236236 142254
rect 236184 142190 236236 142196
rect 236276 142248 236328 142254
rect 236276 142190 236328 142196
rect 236196 142118 236224 142190
rect 236184 142112 236236 142118
rect 236184 142054 236236 142060
rect 236276 120692 236328 120698
rect 236276 120634 236328 120640
rect 236288 115954 236316 120634
rect 236288 115926 236408 115954
rect 236380 109138 236408 115926
rect 236368 109132 236420 109138
rect 236368 109074 236420 109080
rect 236276 108996 236328 109002
rect 236276 108938 236328 108944
rect 236288 106282 236316 108938
rect 236276 106276 236328 106282
rect 236276 106218 236328 106224
rect 236368 96688 236420 96694
rect 236368 96630 236420 96636
rect 236380 89826 236408 96630
rect 236368 89820 236420 89826
rect 236368 89762 236420 89768
rect 236368 89684 236420 89690
rect 236368 89626 236420 89632
rect 236380 86986 236408 89626
rect 236288 86970 236408 86986
rect 236276 86964 236408 86970
rect 236328 86958 236408 86964
rect 236276 86906 236328 86912
rect 236460 75948 236512 75954
rect 236460 75890 236512 75896
rect 236472 67658 236500 75890
rect 236276 67652 236328 67658
rect 236276 67594 236328 67600
rect 236460 67652 236512 67658
rect 236460 67594 236512 67600
rect 236288 61554 236316 67594
rect 236288 61526 236500 61554
rect 236472 60704 236500 61526
rect 236380 60676 236500 60704
rect 236380 48521 236408 60676
rect 236366 48512 236422 48521
rect 236366 48447 236422 48456
rect 236274 48376 236330 48385
rect 236274 48311 236330 48320
rect 236288 41478 236316 48311
rect 236276 41472 236328 41478
rect 236276 41414 236328 41420
rect 236276 41336 236328 41342
rect 236276 41278 236328 41284
rect 236288 31634 236316 41278
rect 236288 31606 236408 31634
rect 236380 28966 236408 31606
rect 236368 28960 236420 28966
rect 236368 28902 236420 28908
rect 236368 19372 236420 19378
rect 236368 19314 236420 19320
rect 236380 5098 236408 19314
rect 236368 5092 236420 5098
rect 236368 5034 236420 5040
rect 236092 3596 236144 3602
rect 236092 3538 236144 3544
rect 236000 3528 236052 3534
rect 236000 3470 236052 3476
rect 236012 400 236040 3470
rect 237300 490 237328 216854
rect 237668 5166 237696 220102
rect 238024 217524 238076 217530
rect 238024 217466 238076 217472
rect 237656 5160 237708 5166
rect 237656 5102 237708 5108
rect 238036 3126 238064 217466
rect 238312 217462 238340 220116
rect 238300 217456 238352 217462
rect 238300 217398 238352 217404
rect 238668 217456 238720 217462
rect 238668 217398 238720 217404
rect 238024 3120 238076 3126
rect 238024 3062 238076 3068
rect 238680 490 238708 217398
rect 238772 217326 238800 220116
rect 238956 220102 239154 220130
rect 238760 217320 238812 217326
rect 238760 217262 238812 217268
rect 238956 5234 238984 220102
rect 239600 217802 239628 220116
rect 239588 217796 239640 217802
rect 239588 217738 239640 217744
rect 239968 217394 239996 220116
rect 240336 220102 240442 220130
rect 239956 217388 240008 217394
rect 239956 217330 240008 217336
rect 239404 216708 239456 216714
rect 239404 216650 239456 216656
rect 238944 5228 238996 5234
rect 238944 5170 238996 5176
rect 239416 3330 239444 216650
rect 240336 5302 240364 220102
rect 240796 217870 240824 220116
rect 240784 217864 240836 217870
rect 240784 217806 240836 217812
rect 241164 217598 241192 220116
rect 241638 220102 241744 220130
rect 241152 217592 241204 217598
rect 241152 217534 241204 217540
rect 240784 217388 240836 217394
rect 240784 217330 240836 217336
rect 240324 5296 240376 5302
rect 240324 5238 240376 5244
rect 240796 4162 240824 217330
rect 241428 217320 241480 217326
rect 241428 217262 241480 217268
rect 240704 4134 240824 4162
rect 240704 3942 240732 4134
rect 241440 4078 241468 217262
rect 241716 5370 241744 220102
rect 241992 216850 242020 220116
rect 242452 217666 242480 220116
rect 242820 217734 242848 220116
rect 243096 220102 243294 220130
rect 242808 217728 242860 217734
rect 242808 217670 242860 217676
rect 242440 217660 242492 217666
rect 242440 217602 242492 217608
rect 241980 216844 242032 216850
rect 241980 216786 242032 216792
rect 242992 210452 243044 210458
rect 242992 210394 243044 210400
rect 241704 5364 241756 5370
rect 241704 5306 241756 5312
rect 240784 4072 240836 4078
rect 240784 4014 240836 4020
rect 241428 4072 241480 4078
rect 241428 4014 241480 4020
rect 240692 3936 240744 3942
rect 240692 3878 240744 3884
rect 239588 3664 239640 3670
rect 239588 3606 239640 3612
rect 239404 3324 239456 3330
rect 239404 3266 239456 3272
rect 237208 462 237328 490
rect 238404 462 238708 490
rect 237208 400 237236 462
rect 238404 400 238432 462
rect 239600 400 239628 3606
rect 240796 400 240824 4014
rect 241980 3936 242032 3942
rect 241980 3878 242032 3884
rect 241992 400 242020 3878
rect 243004 3874 243032 210394
rect 242992 3868 243044 3874
rect 242992 3810 243044 3816
rect 243096 3738 243124 220102
rect 243648 217938 243676 220116
rect 243832 220102 244122 220130
rect 243636 217932 243688 217938
rect 243636 217874 243688 217880
rect 243544 216844 243596 216850
rect 243544 216786 243596 216792
rect 243084 3732 243136 3738
rect 243084 3674 243136 3680
rect 243176 3732 243228 3738
rect 243176 3674 243228 3680
rect 243188 400 243216 3674
rect 243556 3262 243584 216786
rect 243832 210458 243860 220102
rect 244476 218006 244504 220116
rect 244464 218000 244516 218006
rect 244464 217942 244516 217948
rect 244844 216714 244872 220116
rect 245304 217258 245332 220116
rect 245568 217592 245620 217598
rect 245568 217534 245620 217540
rect 245292 217252 245344 217258
rect 245292 217194 245344 217200
rect 244924 216776 244976 216782
rect 244924 216718 244976 216724
rect 244832 216708 244884 216714
rect 244832 216650 244884 216656
rect 243820 210452 243872 210458
rect 243820 210394 243872 210400
rect 244372 3596 244424 3602
rect 244372 3538 244424 3544
rect 243544 3256 243596 3262
rect 243544 3198 243596 3204
rect 244384 400 244412 3538
rect 244936 2990 244964 216718
rect 245016 216708 245068 216714
rect 245016 216650 245068 216656
rect 245028 4146 245056 216650
rect 245016 4140 245068 4146
rect 245016 4082 245068 4088
rect 245580 3602 245608 217534
rect 245672 217530 245700 220116
rect 245660 217524 245712 217530
rect 245660 217466 245712 217472
rect 246132 216714 246160 220116
rect 246500 216986 246528 220116
rect 246488 216980 246540 216986
rect 246488 216922 246540 216928
rect 246960 216850 246988 220116
rect 247328 217190 247356 220116
rect 247316 217184 247368 217190
rect 247316 217126 247368 217132
rect 247696 217122 247724 220116
rect 247776 217660 247828 217666
rect 247776 217602 247828 217608
rect 247684 217116 247736 217122
rect 247684 217058 247736 217064
rect 246948 216844 247000 216850
rect 246948 216786 247000 216792
rect 246120 216708 246172 216714
rect 246120 216650 246172 216656
rect 247684 216708 247736 216714
rect 247684 216650 247736 216656
rect 246764 3800 246816 3806
rect 246764 3742 246816 3748
rect 245568 3596 245620 3602
rect 245568 3538 245620 3544
rect 245568 3392 245620 3398
rect 245568 3334 245620 3340
rect 244924 2984 244976 2990
rect 244924 2926 244976 2932
rect 245580 400 245608 3334
rect 246776 400 246804 3742
rect 247696 3194 247724 216650
rect 247788 4010 247816 217602
rect 248156 216782 248184 220116
rect 248328 217524 248380 217530
rect 248328 217466 248380 217472
rect 248144 216776 248196 216782
rect 248144 216718 248196 216724
rect 247776 4004 247828 4010
rect 247776 3946 247828 3952
rect 247684 3188 247736 3194
rect 247684 3130 247736 3136
rect 248340 490 248368 217466
rect 248524 216714 248552 220116
rect 248984 217054 249012 220116
rect 249076 220102 249366 220130
rect 248972 217048 249024 217054
rect 248972 216990 249024 216996
rect 248512 216708 248564 216714
rect 248512 216650 248564 216656
rect 249076 214554 249104 220102
rect 249340 217048 249392 217054
rect 249340 216990 249392 216996
rect 249156 216708 249208 216714
rect 249156 216650 249208 216656
rect 248616 214526 249104 214554
rect 248616 3058 248644 214526
rect 249168 214418 249196 216650
rect 249076 214390 249196 214418
rect 249076 3466 249104 214390
rect 249352 214282 249380 216990
rect 249812 216714 249840 220116
rect 249904 220102 250194 220130
rect 249904 217394 249932 220102
rect 250640 217666 250668 220116
rect 250732 220102 251022 220130
rect 250628 217660 250680 217666
rect 250628 217602 250680 217608
rect 249892 217388 249944 217394
rect 249892 217330 249944 217336
rect 249800 216708 249852 216714
rect 249800 216650 249852 216656
rect 250732 214554 250760 220102
rect 251376 216918 251404 220116
rect 251836 217462 251864 220116
rect 251824 217456 251876 217462
rect 251824 217398 251876 217404
rect 251364 216912 251416 216918
rect 251364 216854 251416 216860
rect 251916 216912 251968 216918
rect 251916 216854 251968 216860
rect 250904 216844 250956 216850
rect 250904 216786 250956 216792
rect 250812 216776 250864 216782
rect 250812 216718 250864 216724
rect 249168 214254 249380 214282
rect 249996 214526 250760 214554
rect 249168 3942 249196 214254
rect 249156 3936 249208 3942
rect 249156 3878 249208 3884
rect 249996 3534 250024 214526
rect 250824 214418 250852 216718
rect 250456 214390 250852 214418
rect 250456 3670 250484 214390
rect 250916 214282 250944 216786
rect 251824 216708 251876 216714
rect 251824 216650 251876 216656
rect 250548 214254 250944 214282
rect 250444 3664 250496 3670
rect 250444 3606 250496 3612
rect 249984 3528 250036 3534
rect 249984 3470 250036 3476
rect 249064 3460 249116 3466
rect 249064 3402 249116 3408
rect 249156 3460 249208 3466
rect 249156 3402 249208 3408
rect 248604 3052 248656 3058
rect 248604 2994 248656 3000
rect 247972 462 248368 490
rect 247972 400 248000 462
rect 249168 400 249196 3402
rect 250548 3398 250576 214254
rect 251836 3738 251864 216650
rect 251824 3732 251876 3738
rect 251824 3674 251876 3680
rect 251456 3528 251508 3534
rect 251456 3470 251508 3476
rect 250536 3392 250588 3398
rect 250536 3334 250588 3340
rect 250352 3324 250404 3330
rect 250352 3266 250404 3272
rect 250364 400 250392 3266
rect 251468 400 251496 3470
rect 251928 3466 251956 216854
rect 252204 216782 252232 220116
rect 252664 217326 252692 220116
rect 252652 217320 252704 217326
rect 252652 217262 252704 217268
rect 253032 217054 253060 220116
rect 253020 217048 253072 217054
rect 253020 216990 253072 216996
rect 252468 216980 252520 216986
rect 252468 216922 252520 216928
rect 252192 216776 252244 216782
rect 252192 216718 252244 216724
rect 252480 3534 252508 216922
rect 253492 216714 253520 220116
rect 253860 217598 253888 220116
rect 253848 217592 253900 217598
rect 253848 217534 253900 217540
rect 254228 216850 254256 220116
rect 254412 220102 254702 220130
rect 254216 216844 254268 216850
rect 254216 216786 254268 216792
rect 253480 216708 253532 216714
rect 253480 216650 253532 216656
rect 254412 215234 254440 220102
rect 255056 217530 255084 220116
rect 255228 217660 255280 217666
rect 255228 217602 255280 217608
rect 255044 217524 255096 217530
rect 255044 217466 255096 217472
rect 254584 216844 254636 216850
rect 254584 216786 254636 216792
rect 254228 215206 254440 215234
rect 254228 205714 254256 215206
rect 254136 205686 254256 205714
rect 254136 3806 254164 205686
rect 254124 3800 254176 3806
rect 254124 3742 254176 3748
rect 252468 3528 252520 3534
rect 252468 3470 252520 3476
rect 251916 3460 251968 3466
rect 251916 3402 251968 3408
rect 253848 3256 253900 3262
rect 253848 3198 253900 3204
rect 252652 3052 252704 3058
rect 252652 2994 252704 3000
rect 252664 400 252692 2994
rect 253860 400 253888 3198
rect 254596 3058 254624 216786
rect 254584 3052 254636 3058
rect 254584 2994 254636 3000
rect 255240 490 255268 217602
rect 255516 216918 255544 220116
rect 255608 220102 255898 220130
rect 255504 216912 255556 216918
rect 255504 216854 255556 216860
rect 255608 3330 255636 220102
rect 256344 216986 256372 220116
rect 256608 217728 256660 217734
rect 256608 217670 256660 217676
rect 256332 216980 256384 216986
rect 256332 216922 256384 216928
rect 255596 3324 255648 3330
rect 255596 3266 255648 3272
rect 256620 490 256648 217670
rect 256712 216850 256740 220116
rect 256896 220102 257186 220130
rect 256700 216844 256752 216850
rect 256700 216786 256752 216792
rect 256896 3262 256924 220102
rect 257540 217666 257568 220116
rect 257908 217734 257936 220116
rect 258092 220102 258382 220130
rect 258644 220102 258750 220130
rect 259210 220102 259408 220130
rect 257896 217728 257948 217734
rect 258092 217682 258120 220102
rect 258644 217682 258672 220102
rect 257896 217670 257948 217676
rect 257528 217660 257580 217666
rect 257528 217602 257580 217608
rect 258000 217654 258120 217682
rect 258276 217654 258672 217682
rect 258000 4146 258028 217654
rect 258276 207738 258304 217654
rect 258264 207732 258316 207738
rect 258264 207674 258316 207680
rect 258356 202904 258408 202910
rect 258356 202846 258408 202852
rect 258368 167074 258396 202846
rect 258172 167068 258224 167074
rect 258172 167010 258224 167016
rect 258356 167068 258408 167074
rect 258356 167010 258408 167016
rect 258184 166954 258212 167010
rect 258184 166926 258304 166954
rect 258276 164218 258304 166926
rect 258264 164212 258316 164218
rect 258264 164154 258316 164160
rect 258264 157344 258316 157350
rect 258264 157286 258316 157292
rect 258276 154578 258304 157286
rect 258276 154550 258396 154578
rect 258368 147694 258396 154550
rect 258172 147688 258224 147694
rect 258356 147688 258408 147694
rect 258224 147636 258304 147642
rect 258172 147630 258304 147636
rect 258356 147630 258408 147636
rect 258184 147614 258304 147630
rect 258276 144906 258304 147614
rect 258264 144900 258316 144906
rect 258264 144842 258316 144848
rect 258264 137964 258316 137970
rect 258264 137906 258316 137912
rect 258276 135266 258304 137906
rect 258276 135238 258396 135266
rect 258368 128382 258396 135238
rect 258172 128376 258224 128382
rect 258356 128376 258408 128382
rect 258224 128324 258304 128330
rect 258172 128318 258304 128324
rect 258356 128318 258408 128324
rect 258184 128302 258304 128318
rect 258276 125594 258304 128302
rect 258264 125588 258316 125594
rect 258264 125530 258316 125536
rect 258264 118652 258316 118658
rect 258264 118594 258316 118600
rect 258276 115954 258304 118594
rect 258276 115926 258396 115954
rect 258368 109070 258396 115926
rect 258172 109064 258224 109070
rect 258356 109064 258408 109070
rect 258224 109012 258304 109018
rect 258172 109006 258304 109012
rect 258356 109006 258408 109012
rect 258184 108990 258304 109006
rect 258276 106282 258304 108990
rect 258264 106276 258316 106282
rect 258264 106218 258316 106224
rect 258264 99340 258316 99346
rect 258264 99282 258316 99288
rect 258276 96642 258304 99282
rect 258276 96614 258396 96642
rect 258368 89758 258396 96614
rect 258172 89752 258224 89758
rect 258356 89752 258408 89758
rect 258224 89700 258304 89706
rect 258172 89694 258304 89700
rect 258356 89694 258408 89700
rect 258184 89678 258304 89694
rect 258276 86970 258304 89678
rect 258264 86964 258316 86970
rect 258264 86906 258316 86912
rect 258356 77308 258408 77314
rect 258356 77250 258408 77256
rect 258368 77217 258396 77250
rect 258170 77208 258226 77217
rect 258170 77143 258226 77152
rect 258354 77208 258410 77217
rect 258354 77143 258410 77152
rect 258184 70446 258212 77143
rect 258172 70440 258224 70446
rect 258172 70382 258224 70388
rect 258264 70372 258316 70378
rect 258264 70314 258316 70320
rect 258276 60738 258304 70314
rect 258276 60710 258396 60738
rect 258368 48346 258396 60710
rect 258264 48340 258316 48346
rect 258264 48282 258316 48288
rect 258356 48340 258408 48346
rect 258356 48282 258408 48288
rect 258276 41426 258304 48282
rect 258276 41398 258396 41426
rect 258368 38622 258396 41398
rect 258356 38616 258408 38622
rect 258356 38558 258408 38564
rect 258264 31748 258316 31754
rect 258264 31690 258316 31696
rect 258276 22114 258304 31690
rect 258276 22086 258396 22114
rect 258368 12458 258396 22086
rect 258184 12430 258396 12458
rect 258184 4146 258212 12430
rect 259380 4146 259408 220102
rect 259564 211206 259592 220116
rect 260024 217462 260052 220116
rect 260012 217456 260064 217462
rect 260012 217398 260064 217404
rect 260392 211274 260420 220116
rect 260760 217666 260788 220116
rect 260748 217660 260800 217666
rect 260748 217602 260800 217608
rect 261220 217122 261248 220116
rect 261602 220102 261984 220130
rect 262062 220102 262168 220130
rect 261576 217660 261628 217666
rect 261576 217602 261628 217608
rect 261484 217456 261536 217462
rect 261484 217398 261536 217404
rect 261208 217116 261260 217122
rect 261208 217058 261260 217064
rect 260380 211268 260432 211274
rect 260380 211210 260432 211216
rect 259552 211200 259604 211206
rect 259552 211142 259604 211148
rect 261116 211200 261168 211206
rect 261116 211142 261168 211148
rect 261128 182170 261156 211142
rect 261116 182164 261168 182170
rect 261116 182106 261168 182112
rect 261300 182164 261352 182170
rect 261300 182106 261352 182112
rect 261312 172553 261340 182106
rect 261114 172544 261170 172553
rect 261114 172479 261170 172488
rect 261298 172544 261354 172553
rect 261298 172479 261354 172488
rect 261128 162858 261156 172479
rect 261116 162852 261168 162858
rect 261116 162794 261168 162800
rect 261116 153264 261168 153270
rect 261116 153206 261168 153212
rect 261128 143546 261156 153206
rect 261116 143540 261168 143546
rect 261116 143482 261168 143488
rect 261116 133952 261168 133958
rect 261116 133894 261168 133900
rect 261128 124166 261156 133894
rect 261116 124160 261168 124166
rect 261116 124102 261168 124108
rect 261116 114572 261168 114578
rect 261116 114514 261168 114520
rect 261128 104854 261156 114514
rect 261116 104848 261168 104854
rect 261116 104790 261168 104796
rect 261116 95260 261168 95266
rect 261116 95202 261168 95208
rect 261128 85542 261156 95202
rect 261116 85536 261168 85542
rect 261116 85478 261168 85484
rect 260932 75948 260984 75954
rect 260932 75890 260984 75896
rect 260944 67697 260972 75890
rect 260930 67688 260986 67697
rect 260930 67623 260986 67632
rect 261114 67688 261170 67697
rect 261114 67623 261170 67632
rect 261128 57934 261156 67623
rect 261024 57928 261076 57934
rect 261024 57870 261076 57876
rect 261116 57928 261168 57934
rect 261116 57870 261168 57876
rect 261036 56574 261064 57870
rect 261024 56568 261076 56574
rect 261024 56510 261076 56516
rect 261208 56500 261260 56506
rect 261208 56442 261260 56448
rect 261220 46918 261248 56442
rect 261208 46912 261260 46918
rect 261208 46854 261260 46860
rect 261300 46912 261352 46918
rect 261300 46854 261352 46860
rect 261312 38570 261340 46854
rect 261220 38542 261340 38570
rect 261220 29034 261248 38542
rect 261116 29028 261168 29034
rect 261116 28970 261168 28976
rect 261208 29028 261260 29034
rect 261208 28970 261260 28976
rect 261128 27606 261156 28970
rect 261116 27600 261168 27606
rect 261116 27542 261168 27548
rect 261116 18012 261168 18018
rect 261116 17954 261168 17960
rect 261128 12594 261156 17954
rect 261128 12566 261248 12594
rect 261220 12322 261248 12566
rect 261036 12294 261248 12322
rect 257436 4140 257488 4146
rect 257436 4082 257488 4088
rect 257988 4140 258040 4146
rect 257988 4082 258040 4088
rect 258172 4140 258224 4146
rect 258172 4082 258224 4088
rect 258632 4140 258684 4146
rect 258632 4082 258684 4088
rect 259368 4140 259420 4146
rect 259368 4082 259420 4088
rect 259828 4140 259880 4146
rect 259828 4082 259880 4088
rect 256884 3256 256936 3262
rect 256884 3198 256936 3204
rect 255056 462 255268 490
rect 256252 462 256648 490
rect 255056 400 255084 462
rect 256252 400 256280 462
rect 257448 400 257476 4082
rect 258644 400 258672 4082
rect 259840 400 259868 4082
rect 261036 400 261064 12294
rect 261496 4146 261524 217398
rect 261484 4140 261536 4146
rect 261484 4082 261536 4088
rect 261588 4078 261616 217602
rect 261956 211954 261984 220102
rect 261944 211948 261996 211954
rect 261944 211890 261996 211896
rect 261576 4072 261628 4078
rect 261576 4014 261628 4020
rect 262140 3738 262168 220102
rect 262416 217054 262444 220116
rect 262876 217734 262904 220116
rect 263258 220102 263364 220130
rect 262864 217728 262916 217734
rect 262864 217670 262916 217676
rect 262404 217048 262456 217054
rect 262404 216990 262456 216996
rect 262588 211268 262640 211274
rect 262588 211210 262640 211216
rect 262600 211138 262628 211210
rect 262588 211132 262640 211138
rect 262588 211074 262640 211080
rect 262588 205624 262640 205630
rect 262588 205566 262640 205572
rect 262600 201498 262628 205566
rect 262600 201470 262720 201498
rect 262692 196654 262720 201470
rect 262404 196648 262456 196654
rect 262404 196590 262456 196596
rect 262680 196648 262732 196654
rect 262680 196590 262732 196596
rect 262416 191842 262444 196590
rect 262416 191826 262536 191842
rect 262416 191820 262548 191826
rect 262416 191814 262496 191820
rect 262496 191762 262548 191768
rect 262508 191731 262536 191762
rect 262496 186312 262548 186318
rect 262496 186254 262548 186260
rect 262508 182186 262536 186254
rect 262508 182158 262628 182186
rect 262600 182102 262628 182158
rect 262588 182096 262640 182102
rect 262588 182038 262640 182044
rect 262588 172576 262640 172582
rect 262588 172518 262640 172524
rect 262600 166954 262628 172518
rect 262508 166926 262628 166954
rect 262508 164218 262536 166926
rect 262312 164212 262364 164218
rect 262312 164154 262364 164160
rect 262496 164212 262548 164218
rect 262496 164154 262548 164160
rect 262324 154601 262352 164154
rect 262310 154592 262366 154601
rect 262310 154527 262366 154536
rect 262586 154592 262642 154601
rect 262586 154527 262642 154536
rect 262600 147642 262628 154527
rect 262508 147614 262628 147642
rect 262508 140026 262536 147614
rect 262324 139998 262536 140026
rect 262324 135289 262352 139998
rect 262310 135280 262366 135289
rect 262310 135215 262366 135224
rect 262586 135280 262642 135289
rect 262586 135215 262642 135224
rect 262600 128330 262628 135215
rect 262508 128302 262628 128330
rect 262508 120714 262536 128302
rect 262324 120686 262536 120714
rect 262324 115977 262352 120686
rect 262310 115968 262366 115977
rect 262310 115903 262366 115912
rect 262586 115968 262642 115977
rect 262586 115903 262642 115912
rect 262600 109018 262628 115903
rect 262508 108990 262628 109018
rect 262508 101402 262536 108990
rect 262324 101374 262536 101402
rect 262324 96665 262352 101374
rect 262310 96656 262366 96665
rect 262310 96591 262366 96600
rect 262586 96656 262642 96665
rect 262586 96591 262642 96600
rect 262600 89706 262628 96591
rect 262416 89678 262628 89706
rect 262416 86970 262444 89678
rect 262404 86964 262456 86970
rect 262404 86906 262456 86912
rect 262312 77308 262364 77314
rect 262312 77250 262364 77256
rect 262324 70258 262352 77250
rect 262324 70230 262444 70258
rect 262416 60722 262444 70230
rect 262404 60716 262456 60722
rect 262404 60658 262456 60664
rect 262588 60716 262640 60722
rect 262588 60658 262640 60664
rect 262600 57934 262628 60658
rect 262588 57928 262640 57934
rect 262588 57870 262640 57876
rect 262496 48340 262548 48346
rect 262496 48282 262548 48288
rect 262508 41426 262536 48282
rect 262416 41410 262536 41426
rect 262404 41404 262536 41410
rect 262456 41398 262536 41404
rect 262588 41404 262640 41410
rect 262404 41346 262456 41352
rect 262588 41346 262640 41352
rect 262600 31770 262628 41346
rect 262508 31742 262628 31770
rect 262508 22114 262536 31742
rect 262416 22098 262536 22114
rect 262404 22092 262536 22098
rect 262456 22086 262536 22092
rect 262588 22092 262640 22098
rect 262404 22034 262456 22040
rect 262588 22034 262640 22040
rect 262220 4140 262272 4146
rect 262220 4082 262272 4088
rect 262128 3732 262180 3738
rect 262128 3674 262180 3680
rect 262232 400 262260 4082
rect 262600 3346 262628 22034
rect 263336 3466 263364 220102
rect 263508 217728 263560 217734
rect 263508 217670 263560 217676
rect 263416 217048 263468 217054
rect 263416 216990 263468 216996
rect 263428 3602 263456 216990
rect 263520 4078 263548 217670
rect 263704 216918 263732 220116
rect 264072 217394 264100 220116
rect 264440 217666 264468 220116
rect 264900 217734 264928 220116
rect 264888 217728 264940 217734
rect 264888 217670 264940 217676
rect 264428 217660 264480 217666
rect 264428 217602 264480 217608
rect 264060 217388 264112 217394
rect 264060 217330 264112 217336
rect 265268 217326 265296 220116
rect 265742 220102 265940 220130
rect 266110 220102 266308 220130
rect 265624 217728 265676 217734
rect 265624 217670 265676 217676
rect 265912 217682 265940 220102
rect 265256 217320 265308 217326
rect 265256 217262 265308 217268
rect 265256 217048 265308 217054
rect 265256 216990 265308 216996
rect 263692 216912 263744 216918
rect 263692 216854 263744 216860
rect 265268 12442 265296 216990
rect 265256 12436 265308 12442
rect 265256 12378 265308 12384
rect 264612 4140 264664 4146
rect 264612 4082 264664 4088
rect 263508 4072 263560 4078
rect 263508 4014 263560 4020
rect 263416 3596 263468 3602
rect 263416 3538 263468 3544
rect 263324 3460 263376 3466
rect 263324 3402 263376 3408
rect 262600 3318 263456 3346
rect 263428 400 263456 3318
rect 264624 400 264652 4082
rect 265636 3874 265664 217670
rect 265912 217654 266124 217682
rect 266096 215234 266124 217654
rect 266096 215206 266216 215234
rect 265808 12436 265860 12442
rect 265808 12378 265860 12384
rect 265624 3868 265676 3874
rect 265624 3810 265676 3816
rect 265820 400 265848 12378
rect 266188 3670 266216 215206
rect 266176 3664 266228 3670
rect 266176 3606 266228 3612
rect 266280 3534 266308 220102
rect 266556 217054 266584 220116
rect 266924 218006 266952 220116
rect 267306 220102 267596 220130
rect 266912 218000 266964 218006
rect 266912 217942 266964 217948
rect 267004 217388 267056 217394
rect 267004 217330 267056 217336
rect 266544 217048 266596 217054
rect 266544 216990 266596 216996
rect 266544 211948 266596 211954
rect 266544 211890 266596 211896
rect 266556 211138 266584 211890
rect 266544 211132 266596 211138
rect 266544 211074 266596 211080
rect 266728 211132 266780 211138
rect 266728 211074 266780 211080
rect 266740 191865 266768 211074
rect 266542 191856 266598 191865
rect 266542 191791 266598 191800
rect 266726 191856 266782 191865
rect 266726 191791 266782 191800
rect 266556 167090 266584 191791
rect 266464 167062 266584 167090
rect 266464 166954 266492 167062
rect 266464 166926 266584 166954
rect 266556 147778 266584 166926
rect 266464 147750 266584 147778
rect 266464 147642 266492 147750
rect 266464 147614 266584 147642
rect 266556 128466 266584 147614
rect 266464 128438 266584 128466
rect 266464 128330 266492 128438
rect 266464 128302 266584 128330
rect 266556 109154 266584 128302
rect 266464 109126 266584 109154
rect 266464 109018 266492 109126
rect 266464 108990 266584 109018
rect 266556 89842 266584 108990
rect 266464 89814 266584 89842
rect 266464 89706 266492 89814
rect 266464 89678 266584 89706
rect 266556 70394 266584 89678
rect 266464 70366 266584 70394
rect 266464 70258 266492 70366
rect 266464 70230 266584 70258
rect 266556 51082 266584 70230
rect 266464 51054 266584 51082
rect 266464 50946 266492 51054
rect 266464 50918 266584 50946
rect 266556 31890 266584 50918
rect 266544 31884 266596 31890
rect 266544 31826 266596 31832
rect 266544 31748 266596 31754
rect 266544 31690 266596 31696
rect 266556 23662 266584 31690
rect 266544 23656 266596 23662
rect 266544 23598 266596 23604
rect 266820 23656 266872 23662
rect 266820 23598 266872 23604
rect 266832 19258 266860 23598
rect 266832 19230 266952 19258
rect 266268 3528 266320 3534
rect 266268 3470 266320 3476
rect 266924 3210 266952 19230
rect 267016 3398 267044 217330
rect 267568 4010 267596 220102
rect 267752 217734 267780 220116
rect 268134 220102 268516 220130
rect 268594 220102 268884 220130
rect 268962 220102 269068 220130
rect 267740 217728 267792 217734
rect 267740 217670 267792 217676
rect 267648 217048 267700 217054
rect 267648 216990 267700 216996
rect 267556 4004 267608 4010
rect 267556 3946 267608 3952
rect 267660 3806 267688 216990
rect 268488 215234 268516 220102
rect 268488 215206 268700 215234
rect 268672 195922 268700 215206
rect 268672 195894 268792 195922
rect 268764 167090 268792 195894
rect 268672 167062 268792 167090
rect 268672 166954 268700 167062
rect 268672 166926 268792 166954
rect 268764 147778 268792 166926
rect 268672 147750 268792 147778
rect 268672 147642 268700 147750
rect 268672 147614 268792 147642
rect 268764 128466 268792 147614
rect 268672 128438 268792 128466
rect 268672 128330 268700 128438
rect 268672 128302 268792 128330
rect 268764 109154 268792 128302
rect 268672 109126 268792 109154
rect 268672 109018 268700 109126
rect 268672 108990 268792 109018
rect 268764 89842 268792 108990
rect 268672 89814 268792 89842
rect 268672 89706 268700 89814
rect 268672 89678 268792 89706
rect 268764 70394 268792 89678
rect 268672 70366 268792 70394
rect 268672 70258 268700 70366
rect 268672 70230 268792 70258
rect 268764 51082 268792 70230
rect 268672 51054 268792 51082
rect 268672 50946 268700 51054
rect 268672 50918 268792 50946
rect 268764 29209 268792 50918
rect 268750 29200 268806 29209
rect 268750 29135 268806 29144
rect 268750 29064 268806 29073
rect 268750 28999 268806 29008
rect 268764 27606 268792 28999
rect 268752 27600 268804 27606
rect 268752 27542 268804 27548
rect 268752 18012 268804 18018
rect 268752 17954 268804 17960
rect 268764 3942 268792 17954
rect 268752 3936 268804 3942
rect 268752 3878 268804 3884
rect 267648 3800 267700 3806
rect 267648 3742 267700 3748
rect 268108 3732 268160 3738
rect 268108 3674 268160 3680
rect 267004 3392 267056 3398
rect 267004 3334 267056 3340
rect 266924 3182 267044 3210
rect 267016 400 267044 3182
rect 268120 400 268148 3674
rect 268856 3330 268884 220102
rect 268936 217728 268988 217734
rect 268936 217670 268988 217676
rect 268844 3324 268896 3330
rect 268844 3266 268896 3272
rect 268948 2854 268976 217670
rect 269040 2922 269068 220102
rect 269408 217462 269436 220116
rect 269790 220102 270172 220130
rect 270250 220102 270448 220130
rect 269396 217456 269448 217462
rect 269396 217398 269448 217404
rect 269764 216912 269816 216918
rect 269764 216854 269816 216860
rect 269776 4146 269804 216854
rect 270144 210458 270172 220102
rect 270224 217456 270276 217462
rect 270224 217398 270276 217404
rect 270132 210452 270184 210458
rect 270132 210394 270184 210400
rect 270132 189916 270184 189922
rect 270132 189858 270184 189864
rect 270144 181490 270172 189858
rect 270132 181484 270184 181490
rect 270132 181426 270184 181432
rect 270132 170604 270184 170610
rect 270132 170546 270184 170552
rect 270144 162178 270172 170546
rect 270132 162172 270184 162178
rect 270132 162114 270184 162120
rect 270132 152516 270184 152522
rect 270132 152458 270184 152464
rect 270144 142866 270172 152458
rect 270132 142860 270184 142866
rect 270132 142802 270184 142808
rect 270132 131980 270184 131986
rect 270132 131922 270184 131928
rect 270144 123554 270172 131922
rect 270132 123548 270184 123554
rect 270132 123490 270184 123496
rect 270132 113892 270184 113898
rect 270132 113834 270184 113840
rect 270144 105466 270172 113834
rect 270132 105460 270184 105466
rect 270132 105402 270184 105408
rect 270132 94580 270184 94586
rect 270132 94522 270184 94528
rect 270144 86154 270172 94522
rect 270132 86148 270184 86154
rect 270132 86090 270184 86096
rect 270132 75268 270184 75274
rect 270132 75210 270184 75216
rect 270144 65550 270172 75210
rect 270132 65544 270184 65550
rect 270132 65486 270184 65492
rect 270132 54664 270184 54670
rect 270132 54606 270184 54612
rect 270144 47462 270172 54606
rect 270132 47456 270184 47462
rect 270132 47398 270184 47404
rect 270132 35352 270184 35358
rect 270132 35294 270184 35300
rect 270144 26926 270172 35294
rect 270132 26920 270184 26926
rect 270132 26862 270184 26868
rect 270132 17264 270184 17270
rect 270132 17206 270184 17212
rect 269764 4140 269816 4146
rect 269764 4082 269816 4088
rect 270144 3602 270172 17206
rect 269304 3596 269356 3602
rect 269304 3538 269356 3544
rect 270132 3596 270184 3602
rect 270132 3538 270184 3544
rect 269028 2916 269080 2922
rect 269028 2858 269080 2864
rect 268936 2848 268988 2854
rect 268936 2790 268988 2796
rect 269316 400 269344 3538
rect 270236 2990 270264 217398
rect 270316 210452 270368 210458
rect 270316 210394 270368 210400
rect 270328 189922 270356 210394
rect 270316 189916 270368 189922
rect 270316 189858 270368 189864
rect 270316 181484 270368 181490
rect 270316 181426 270368 181432
rect 270328 170610 270356 181426
rect 270316 170604 270368 170610
rect 270316 170546 270368 170552
rect 270316 162172 270368 162178
rect 270316 162114 270368 162120
rect 270328 152522 270356 162114
rect 270316 152516 270368 152522
rect 270316 152458 270368 152464
rect 270316 142860 270368 142866
rect 270316 142802 270368 142808
rect 270328 131986 270356 142802
rect 270316 131980 270368 131986
rect 270316 131922 270368 131928
rect 270316 123548 270368 123554
rect 270316 123490 270368 123496
rect 270328 113898 270356 123490
rect 270316 113892 270368 113898
rect 270316 113834 270368 113840
rect 270316 105460 270368 105466
rect 270316 105402 270368 105408
rect 270328 94586 270356 105402
rect 270316 94580 270368 94586
rect 270316 94522 270368 94528
rect 270316 86148 270368 86154
rect 270316 86090 270368 86096
rect 270328 75274 270356 86090
rect 270316 75268 270368 75274
rect 270316 75210 270368 75216
rect 270316 65544 270368 65550
rect 270316 65486 270368 65492
rect 270328 54670 270356 65486
rect 270316 54664 270368 54670
rect 270316 54606 270368 54612
rect 270316 47456 270368 47462
rect 270316 47398 270368 47404
rect 270328 35358 270356 47398
rect 270316 35352 270368 35358
rect 270316 35294 270368 35300
rect 270316 26920 270368 26926
rect 270316 26862 270368 26868
rect 270328 17270 270356 26862
rect 270316 17264 270368 17270
rect 270316 17206 270368 17212
rect 270420 3738 270448 220102
rect 270604 217734 270632 220116
rect 270592 217728 270644 217734
rect 270592 217670 270644 217676
rect 270972 216986 271000 220116
rect 270960 216980 271012 216986
rect 270960 216922 271012 216928
rect 271432 216850 271460 220116
rect 271800 217938 271828 220116
rect 271788 217932 271840 217938
rect 271788 217874 271840 217880
rect 271788 217728 271840 217734
rect 271788 217670 271840 217676
rect 271420 216844 271472 216850
rect 271420 216786 271472 216792
rect 270500 40248 270552 40254
rect 270498 40216 270500 40225
rect 270552 40216 270554 40225
rect 270498 40151 270554 40160
rect 270500 4072 270552 4078
rect 270500 4014 270552 4020
rect 270408 3732 270460 3738
rect 270408 3674 270460 3680
rect 270224 2984 270276 2990
rect 270224 2926 270276 2932
rect 270512 400 270540 4014
rect 271696 3460 271748 3466
rect 271696 3402 271748 3408
rect 271708 400 271736 3402
rect 271800 3194 271828 217670
rect 272260 217054 272288 220116
rect 272642 220102 273024 220130
rect 273102 220102 273208 220130
rect 272524 217660 272576 217666
rect 272524 217602 272576 217608
rect 272248 217048 272300 217054
rect 272248 216990 272300 216996
rect 272536 3534 272564 217602
rect 272996 205714 273024 220102
rect 272904 205686 273024 205714
rect 272904 205578 272932 205686
rect 272904 205550 273024 205578
rect 272996 196058 273024 205550
rect 272996 196030 273116 196058
rect 273088 193202 273116 196030
rect 272996 193174 273116 193202
rect 272996 172689 273024 193174
rect 272982 172680 273038 172689
rect 272982 172615 273038 172624
rect 273074 172544 273130 172553
rect 273074 172479 273130 172488
rect 273088 167142 273116 172479
rect 273076 167136 273128 167142
rect 273076 167078 273128 167084
rect 272984 166932 273036 166938
rect 272984 166874 273036 166880
rect 272996 158030 273024 166874
rect 272984 158024 273036 158030
rect 272984 157966 273036 157972
rect 273180 154698 273208 220102
rect 273456 216918 273484 220116
rect 273824 217462 273852 220116
rect 274298 220102 274588 220130
rect 273812 217456 273864 217462
rect 273812 217398 273864 217404
rect 273444 216912 273496 216918
rect 273444 216854 273496 216860
rect 273904 216844 273956 216850
rect 273904 216786 273956 216792
rect 273260 158024 273312 158030
rect 273260 157966 273312 157972
rect 273168 154692 273220 154698
rect 273168 154634 273220 154640
rect 273168 154556 273220 154562
rect 273168 154498 273220 154504
rect 273076 147756 273128 147762
rect 273076 147698 273128 147704
rect 273088 135250 273116 147698
rect 272984 135244 273036 135250
rect 272984 135186 273036 135192
rect 273076 135244 273128 135250
rect 273076 135186 273128 135192
rect 272996 128364 273024 135186
rect 272996 128336 273116 128364
rect 273088 115938 273116 128336
rect 273076 115932 273128 115938
rect 273076 115874 273128 115880
rect 273076 106344 273128 106350
rect 273076 106286 273128 106292
rect 273088 51134 273116 106286
rect 273076 51128 273128 51134
rect 273076 51070 273128 51076
rect 272984 51060 273036 51066
rect 272984 51002 273036 51008
rect 272996 45558 273024 51002
rect 272984 45552 273036 45558
rect 272984 45494 273036 45500
rect 272984 37188 273036 37194
rect 272984 37130 273036 37136
rect 272996 27742 273024 37130
rect 272984 27736 273036 27742
rect 272984 27678 273036 27684
rect 273076 27668 273128 27674
rect 273076 27610 273128 27616
rect 273088 22250 273116 27610
rect 272904 22222 273116 22250
rect 272904 18018 272932 22222
rect 272800 18012 272852 18018
rect 272800 17954 272852 17960
rect 272892 18012 272944 18018
rect 272892 17954 272944 17960
rect 272812 4010 272840 17954
rect 272892 4140 272944 4146
rect 272892 4082 272944 4088
rect 272800 4004 272852 4010
rect 272800 3946 272852 3952
rect 272524 3528 272576 3534
rect 272524 3470 272576 3476
rect 271788 3188 271840 3194
rect 271788 3130 271840 3136
rect 272904 400 272932 4082
rect 273180 3126 273208 154498
rect 273272 147762 273300 157966
rect 273260 147756 273312 147762
rect 273260 147698 273312 147704
rect 273916 7698 273944 216786
rect 273916 7670 274220 7698
rect 274192 3398 274220 7670
rect 274088 3392 274140 3398
rect 274088 3334 274140 3340
rect 274180 3392 274232 3398
rect 274180 3334 274232 3340
rect 273168 3120 273220 3126
rect 273168 3062 273220 3068
rect 274100 400 274128 3334
rect 274560 3058 274588 220102
rect 274652 217122 274680 220116
rect 275112 217190 275140 220116
rect 275480 219609 275508 220116
rect 275466 219600 275522 219609
rect 275466 219535 275522 219544
rect 275834 219464 275890 219473
rect 275834 219399 275890 219408
rect 275100 217184 275152 217190
rect 275100 217126 275152 217132
rect 274640 217116 274692 217122
rect 274640 217058 274692 217064
rect 275848 209778 275876 219399
rect 275940 217977 275968 220116
rect 275926 217968 275982 217977
rect 275926 217903 275982 217912
rect 275928 217796 275980 217802
rect 275928 217738 275980 217744
rect 275940 217705 275968 217738
rect 275926 217696 275982 217705
rect 275926 217631 275982 217640
rect 276308 217394 276336 220116
rect 276296 217388 276348 217394
rect 276296 217330 276348 217336
rect 276664 217320 276716 217326
rect 276664 217262 276716 217268
rect 275836 209772 275888 209778
rect 275836 209714 275888 209720
rect 276112 209772 276164 209778
rect 276112 209714 276164 209720
rect 276124 195294 276152 209714
rect 275836 195288 275888 195294
rect 275836 195230 275888 195236
rect 276112 195288 276164 195294
rect 276112 195230 276164 195236
rect 275848 183666 275876 195230
rect 275836 183660 275888 183666
rect 275836 183602 275888 183608
rect 275836 183524 275888 183530
rect 275836 183466 275888 183472
rect 275848 180810 275876 183466
rect 275836 180804 275888 180810
rect 275836 180746 275888 180752
rect 275928 171148 275980 171154
rect 275928 171090 275980 171096
rect 275940 162858 275968 171090
rect 275836 162852 275888 162858
rect 275836 162794 275888 162800
rect 275928 162852 275980 162858
rect 275928 162794 275980 162800
rect 275848 144922 275876 162794
rect 275848 144894 275968 144922
rect 275940 143546 275968 144894
rect 275928 143540 275980 143546
rect 275928 143482 275980 143488
rect 275836 133952 275888 133958
rect 275836 133894 275888 133900
rect 275848 130370 275876 133894
rect 275848 130342 275968 130370
rect 275940 124166 275968 130342
rect 275928 124160 275980 124166
rect 275928 124102 275980 124108
rect 276020 124160 276072 124166
rect 276020 124102 276072 124108
rect 276032 110922 276060 124102
rect 275940 110894 276060 110922
rect 275940 104854 275968 110894
rect 275928 104848 275980 104854
rect 275928 104790 275980 104796
rect 275836 95260 275888 95266
rect 275836 95202 275888 95208
rect 275848 89672 275876 95202
rect 275848 89644 275968 89672
rect 275940 84182 275968 89644
rect 275744 84176 275796 84182
rect 275744 84118 275796 84124
rect 275928 84176 275980 84182
rect 275928 84118 275980 84124
rect 275756 74610 275784 84118
rect 275756 74582 275876 74610
rect 275848 66230 275876 74582
rect 275836 66224 275888 66230
rect 275836 66166 275888 66172
rect 276020 66156 276072 66162
rect 276020 66098 276072 66104
rect 276032 64954 276060 66098
rect 275940 64926 276060 64954
rect 275940 63510 275968 64926
rect 275928 63504 275980 63510
rect 275928 63446 275980 63452
rect 275744 53848 275796 53854
rect 275744 53790 275796 53796
rect 275756 53174 275784 53790
rect 275744 53168 275796 53174
rect 275744 53110 275796 53116
rect 275928 53168 275980 53174
rect 275928 53110 275980 53116
rect 275940 48278 275968 53110
rect 275836 48272 275888 48278
rect 275836 48214 275888 48220
rect 275928 48272 275980 48278
rect 275928 48214 275980 48220
rect 275744 40248 275796 40254
rect 275742 40216 275744 40225
rect 275796 40216 275798 40225
rect 275742 40151 275798 40160
rect 275848 38622 275876 48214
rect 275836 38616 275888 38622
rect 275836 38558 275888 38564
rect 275928 33244 275980 33250
rect 275928 33186 275980 33192
rect 275940 27606 275968 33186
rect 275928 27600 275980 27606
rect 275928 27542 275980 27548
rect 275928 18012 275980 18018
rect 275928 17954 275980 17960
rect 275284 3528 275336 3534
rect 275284 3470 275336 3476
rect 274548 3052 274600 3058
rect 274548 2994 274600 3000
rect 275296 400 275324 3470
rect 275940 3262 275968 17954
rect 276676 4146 276704 217262
rect 277044 212514 277072 220238
rect 277136 217598 277164 220116
rect 277124 217592 277176 217598
rect 277124 217534 277176 217540
rect 277504 217394 277532 220116
rect 277964 217734 277992 220116
rect 278332 217802 278360 220116
rect 278320 217796 278372 217802
rect 278320 217738 278372 217744
rect 277952 217728 278004 217734
rect 277952 217670 278004 217676
rect 278688 217728 278740 217734
rect 278688 217670 278740 217676
rect 277308 217388 277360 217394
rect 277308 217330 277360 217336
rect 277492 217388 277544 217394
rect 277492 217330 277544 217336
rect 276952 212486 277072 212514
rect 276952 201521 276980 212486
rect 276938 201512 276994 201521
rect 276938 201447 276994 201456
rect 277214 201512 277270 201521
rect 277214 201447 277270 201456
rect 277228 200122 277256 201447
rect 277216 200116 277268 200122
rect 277216 200058 277268 200064
rect 277216 183592 277268 183598
rect 277216 183534 277268 183540
rect 277228 182170 277256 183534
rect 277216 182164 277268 182170
rect 277216 182106 277268 182112
rect 277124 172576 277176 172582
rect 277124 172518 277176 172524
rect 277136 167634 277164 172518
rect 277044 167606 277164 167634
rect 277044 162897 277072 167606
rect 277030 162888 277086 162897
rect 277030 162823 277086 162832
rect 277122 153232 277178 153241
rect 277032 153196 277084 153202
rect 277122 153167 277124 153176
rect 277032 153138 277084 153144
rect 277176 153167 277178 153176
rect 277124 153138 277176 153144
rect 277044 143585 277072 153138
rect 277030 143576 277086 143585
rect 277030 143511 277086 143520
rect 277214 143576 277270 143585
rect 277214 143511 277270 143520
rect 277228 133890 277256 143511
rect 277216 133884 277268 133890
rect 277216 133826 277268 133832
rect 277216 124228 277268 124234
rect 277216 124170 277268 124176
rect 277228 118794 277256 124170
rect 277216 118788 277268 118794
rect 277216 118730 277268 118736
rect 277216 104984 277268 104990
rect 277216 104926 277268 104932
rect 277228 104854 277256 104926
rect 277216 104848 277268 104854
rect 277216 104790 277268 104796
rect 277124 95260 277176 95266
rect 277124 95202 277176 95208
rect 277136 89706 277164 95202
rect 277136 89678 277256 89706
rect 277228 74662 277256 89678
rect 277124 74656 277176 74662
rect 277124 74598 277176 74604
rect 277216 74656 277268 74662
rect 277216 74598 277268 74604
rect 277136 69714 277164 74598
rect 277136 69686 277256 69714
rect 277228 63510 277256 69686
rect 277216 63504 277268 63510
rect 277216 63446 277268 63452
rect 277216 48340 277268 48346
rect 277216 48282 277268 48288
rect 277228 38706 277256 48282
rect 277136 38678 277256 38706
rect 277136 31498 277164 38678
rect 277136 31470 277256 31498
rect 277228 27606 277256 31470
rect 277216 27600 277268 27606
rect 277216 27542 277268 27548
rect 277216 9716 277268 9722
rect 277216 9658 277268 9664
rect 277228 4214 277256 9658
rect 277216 4208 277268 4214
rect 277216 4150 277268 4156
rect 276664 4140 276716 4146
rect 276664 4082 276716 4088
rect 276480 4072 276532 4078
rect 276480 4014 276532 4020
rect 275928 3256 275980 3262
rect 275928 3198 275980 3204
rect 276492 400 276520 4014
rect 277320 3330 277348 217330
rect 277676 4140 277728 4146
rect 277676 4082 277728 4088
rect 277216 3324 277268 3330
rect 277216 3266 277268 3272
rect 277308 3324 277360 3330
rect 277308 3266 277360 3272
rect 277228 3097 277256 3266
rect 277214 3088 277270 3097
rect 277214 3023 277270 3032
rect 277688 400 277716 4082
rect 278700 3738 278728 217670
rect 278792 217258 278820 220116
rect 279160 217734 279188 220116
rect 279424 218000 279476 218006
rect 279424 217942 279476 217948
rect 279148 217728 279200 217734
rect 279148 217670 279200 217676
rect 278780 217252 278832 217258
rect 278780 217194 278832 217200
rect 279436 4146 279464 217942
rect 279620 217666 279648 220116
rect 279608 217660 279660 217666
rect 279608 217602 279660 217608
rect 279988 4214 280016 220116
rect 280356 217734 280384 220116
rect 280068 217728 280120 217734
rect 280068 217670 280120 217676
rect 280344 217728 280396 217734
rect 280344 217670 280396 217676
rect 279976 4208 280028 4214
rect 279976 4150 280028 4156
rect 279424 4140 279476 4146
rect 279424 4082 279476 4088
rect 280080 3806 280108 217670
rect 280816 217326 280844 220116
rect 281198 220102 281396 220130
rect 280804 217320 280856 217326
rect 280804 217262 280856 217268
rect 281368 4282 281396 220102
rect 281448 217728 281500 217734
rect 281448 217670 281500 217676
rect 281356 4276 281408 4282
rect 281356 4218 281408 4224
rect 278872 3800 278924 3806
rect 278872 3742 278924 3748
rect 280068 3800 280120 3806
rect 280068 3742 280120 3748
rect 278688 3732 278740 3738
rect 278688 3674 278740 3680
rect 278884 400 278912 3742
rect 281460 3670 281488 217670
rect 281644 217530 281672 220116
rect 282012 218006 282040 220116
rect 282000 218000 282052 218006
rect 282000 217942 282052 217948
rect 281632 217524 281684 217530
rect 281632 217466 281684 217472
rect 282472 211177 282500 220116
rect 282840 216918 282868 220116
rect 283208 217938 283236 220116
rect 283682 220102 283788 220130
rect 284050 220102 284248 220130
rect 283196 217932 283248 217938
rect 283196 217874 283248 217880
rect 283656 217252 283708 217258
rect 283656 217194 283708 217200
rect 283564 216980 283616 216986
rect 283564 216922 283616 216928
rect 282828 216912 282880 216918
rect 282828 216854 282880 216860
rect 282458 211168 282514 211177
rect 282458 211103 282514 211112
rect 282642 211168 282698 211177
rect 282642 211103 282698 211112
rect 282656 205562 282684 211103
rect 282644 205556 282696 205562
rect 282644 205498 282696 205504
rect 282828 205556 282880 205562
rect 282828 205498 282880 205504
rect 282840 201482 282868 205498
rect 282828 201476 282880 201482
rect 282828 201418 282880 201424
rect 282828 193180 282880 193186
rect 282828 193122 282880 193128
rect 282840 191842 282868 193122
rect 282840 191814 282960 191842
rect 282932 183598 282960 191814
rect 282736 183592 282788 183598
rect 282734 183560 282736 183569
rect 282920 183592 282972 183598
rect 282788 183560 282790 183569
rect 282734 183495 282790 183504
rect 282918 183560 282920 183569
rect 282972 183560 282974 183569
rect 282918 183495 282974 183504
rect 282932 182170 282960 183495
rect 282828 182164 282880 182170
rect 282828 182106 282880 182112
rect 282920 182164 282972 182170
rect 282920 182106 282972 182112
rect 282840 164257 282868 182106
rect 282642 164248 282698 164257
rect 282642 164183 282698 164192
rect 282826 164248 282882 164257
rect 282826 164183 282882 164192
rect 282656 162858 282684 164183
rect 282644 162852 282696 162858
rect 282644 162794 282696 162800
rect 282828 162852 282880 162858
rect 282828 162794 282880 162800
rect 282840 128364 282868 162794
rect 282748 128336 282868 128364
rect 282748 125610 282776 128336
rect 282748 125582 282868 125610
rect 282840 116006 282868 125582
rect 282828 116000 282880 116006
rect 282828 115942 282880 115948
rect 282736 114572 282788 114578
rect 282736 114514 282788 114520
rect 282748 104854 282776 114514
rect 282736 104848 282788 104854
rect 282736 104790 282788 104796
rect 282736 95260 282788 95266
rect 282736 95202 282788 95208
rect 282748 89026 282776 95202
rect 282748 88998 282868 89026
rect 282840 77382 282868 88998
rect 282828 77376 282880 77382
rect 282828 77318 282880 77324
rect 282736 75948 282788 75954
rect 282736 75890 282788 75896
rect 282748 67658 282776 75890
rect 282736 67652 282788 67658
rect 282736 67594 282788 67600
rect 282828 67652 282880 67658
rect 282828 67594 282880 67600
rect 282840 53122 282868 67594
rect 282748 53094 282868 53122
rect 282748 48278 282776 53094
rect 282736 48272 282788 48278
rect 282736 48214 282788 48220
rect 282828 48272 282880 48278
rect 282828 48214 282880 48220
rect 282840 37330 282868 48214
rect 282736 37324 282788 37330
rect 282736 37266 282788 37272
rect 282828 37324 282880 37330
rect 282828 37266 282880 37272
rect 282748 26330 282776 37266
rect 282748 26302 282868 26330
rect 282840 12458 282868 26302
rect 282840 12430 282960 12458
rect 282932 12322 282960 12430
rect 282748 12294 282960 12322
rect 282748 4350 282776 12294
rect 282736 4344 282788 4350
rect 282736 4286 282788 4292
rect 282460 4140 282512 4146
rect 282460 4082 282512 4088
rect 281264 3664 281316 3670
rect 281264 3606 281316 3612
rect 281448 3664 281500 3670
rect 281448 3606 281500 3612
rect 280068 3392 280120 3398
rect 280068 3334 280120 3340
rect 280080 400 280108 3334
rect 280434 3088 280490 3097
rect 280434 3023 280436 3032
rect 280488 3023 280490 3032
rect 280436 2994 280488 3000
rect 281276 400 281304 3606
rect 282472 400 282500 4082
rect 283576 2786 283604 216922
rect 283668 4146 283696 217194
rect 283760 212566 283788 220102
rect 284116 217932 284168 217938
rect 284116 217874 284168 217880
rect 283748 212560 283800 212566
rect 283748 212502 283800 212508
rect 284024 212560 284076 212566
rect 284024 212502 284076 212508
rect 284036 211138 284064 212502
rect 283840 211132 283892 211138
rect 283840 211074 283892 211080
rect 284024 211132 284076 211138
rect 284024 211074 284076 211080
rect 283852 201521 283880 211074
rect 283838 201512 283894 201521
rect 283838 201447 283894 201456
rect 284022 201512 284078 201521
rect 284022 201447 284078 201456
rect 284036 191826 284064 201447
rect 283840 191820 283892 191826
rect 283840 191762 283892 191768
rect 284024 191820 284076 191826
rect 284024 191762 284076 191768
rect 283852 182209 283880 191762
rect 283838 182200 283894 182209
rect 283838 182135 283894 182144
rect 284022 182200 284078 182209
rect 284022 182135 284078 182144
rect 284036 172514 284064 182135
rect 283840 172508 283892 172514
rect 283840 172450 283892 172456
rect 284024 172508 284076 172514
rect 284024 172450 284076 172456
rect 283852 162897 283880 172450
rect 283838 162888 283894 162897
rect 283838 162823 283894 162832
rect 284022 162888 284078 162897
rect 284022 162823 284078 162832
rect 284036 154714 284064 162823
rect 283944 154686 284064 154714
rect 283944 153270 283972 154686
rect 283840 153264 283892 153270
rect 283840 153206 283892 153212
rect 283932 153264 283984 153270
rect 283932 153206 283984 153212
rect 283852 147744 283880 153206
rect 283852 147716 283972 147744
rect 283944 138666 283972 147716
rect 283852 138638 283972 138666
rect 283852 137986 283880 138638
rect 283852 137958 283972 137986
rect 283944 133906 283972 137958
rect 283944 133890 284064 133906
rect 283944 133884 284076 133890
rect 283944 133878 284024 133884
rect 284024 133826 284076 133832
rect 284036 133795 284064 133826
rect 284022 106312 284078 106321
rect 284022 106247 284078 106256
rect 284036 104854 284064 106247
rect 284024 104848 284076 104854
rect 284024 104790 284076 104796
rect 283932 95260 283984 95266
rect 283932 95202 283984 95208
rect 283944 85542 283972 95202
rect 283932 85536 283984 85542
rect 283932 85478 283984 85484
rect 284024 75948 284076 75954
rect 284024 75890 284076 75896
rect 284036 66230 284064 75890
rect 284024 66224 284076 66230
rect 284024 66166 284076 66172
rect 283932 56704 283984 56710
rect 283932 56646 283984 56652
rect 283944 56574 283972 56646
rect 283932 56568 283984 56574
rect 283932 56510 283984 56516
rect 284024 46980 284076 46986
rect 284024 46922 284076 46928
rect 284036 46866 284064 46922
rect 283944 46838 284064 46866
rect 283944 38554 283972 46838
rect 284128 38758 284156 217874
rect 284220 38758 284248 220102
rect 284496 217938 284524 220116
rect 284484 217932 284536 217938
rect 284484 217874 284536 217880
rect 284864 212566 284892 220116
rect 285338 220102 285628 220130
rect 285496 217932 285548 217938
rect 285496 217874 285548 217880
rect 284852 212560 284904 212566
rect 285312 212560 285364 212566
rect 284852 212502 284904 212508
rect 285232 212508 285312 212514
rect 285232 212502 285364 212508
rect 285232 212486 285352 212502
rect 285232 192001 285260 212486
rect 285218 191992 285274 192001
rect 285218 191927 285274 191936
rect 285310 191856 285366 191865
rect 285310 191791 285366 191800
rect 285324 183546 285352 191791
rect 285232 183518 285352 183546
rect 285232 182170 285260 183518
rect 285220 182164 285272 182170
rect 285220 182106 285272 182112
rect 285312 166932 285364 166938
rect 285312 166874 285364 166880
rect 285324 159338 285352 166874
rect 285324 159310 285444 159338
rect 285416 144922 285444 159310
rect 285324 144894 285444 144922
rect 285324 143546 285352 144894
rect 285312 143540 285364 143546
rect 285312 143482 285364 143488
rect 285312 137964 285364 137970
rect 285312 137906 285364 137912
rect 285324 133906 285352 137906
rect 284300 133884 284352 133890
rect 285324 133878 285444 133906
rect 284300 133826 284352 133832
rect 284312 124273 284340 133826
rect 285416 125662 285444 133878
rect 285312 125656 285364 125662
rect 285312 125598 285364 125604
rect 285404 125656 285456 125662
rect 285404 125598 285456 125604
rect 284298 124264 284354 124273
rect 284298 124199 284354 124208
rect 285324 120714 285352 125598
rect 285324 120686 285444 120714
rect 285416 109138 285444 120686
rect 285404 109132 285456 109138
rect 285404 109074 285456 109080
rect 285312 108996 285364 109002
rect 285312 108938 285364 108944
rect 285324 101402 285352 108938
rect 285324 101374 285444 101402
rect 285416 89808 285444 101374
rect 285324 89780 285444 89808
rect 285324 80730 285352 89780
rect 285232 80702 285352 80730
rect 285232 67658 285260 80702
rect 285220 67652 285272 67658
rect 285220 67594 285272 67600
rect 285312 67652 285364 67658
rect 285312 67594 285364 67600
rect 285324 66230 285352 67594
rect 285312 66224 285364 66230
rect 285312 66166 285364 66172
rect 285404 56636 285456 56642
rect 285404 56578 285456 56584
rect 285416 48346 285444 56578
rect 285312 48340 285364 48346
rect 285312 48282 285364 48288
rect 285404 48340 285456 48346
rect 285404 48282 285456 48288
rect 285324 43466 285352 48282
rect 285324 43438 285444 43466
rect 284116 38752 284168 38758
rect 284116 38694 284168 38700
rect 284208 38752 284260 38758
rect 284208 38694 284260 38700
rect 284116 38616 284168 38622
rect 284116 38558 284168 38564
rect 284208 38616 284260 38622
rect 284208 38558 284260 38564
rect 283932 38548 283984 38554
rect 283932 38490 283984 38496
rect 284128 33862 284156 38558
rect 284116 33856 284168 33862
rect 284116 33798 284168 33804
rect 284116 33720 284168 33726
rect 284116 33662 284168 33668
rect 284024 29028 284076 29034
rect 284024 28970 284076 28976
rect 284036 9790 284064 28970
rect 284024 9784 284076 9790
rect 284024 9726 284076 9732
rect 283932 8356 283984 8362
rect 283932 8298 283984 8304
rect 283944 4554 283972 8298
rect 283932 4548 283984 4554
rect 283932 4490 283984 4496
rect 284128 4418 284156 33662
rect 284116 4412 284168 4418
rect 284116 4354 284168 4360
rect 283656 4140 283708 4146
rect 283656 4082 283708 4088
rect 283656 3936 283708 3942
rect 283656 3878 283708 3884
rect 283564 2780 283616 2786
rect 283564 2722 283616 2728
rect 283668 400 283696 3878
rect 284220 3369 284248 38558
rect 284300 38548 284352 38554
rect 284300 38490 284352 38496
rect 284312 29034 284340 38490
rect 285416 31822 285444 43438
rect 285404 31816 285456 31822
rect 285404 31758 285456 31764
rect 285312 31748 285364 31754
rect 285312 31690 285364 31696
rect 284300 29028 284352 29034
rect 284300 28970 284352 28976
rect 285324 26330 285352 31690
rect 285324 26302 285444 26330
rect 285416 12510 285444 26302
rect 285404 12504 285456 12510
rect 285404 12446 285456 12452
rect 285312 12436 285364 12442
rect 285312 12378 285364 12384
rect 285324 4622 285352 12378
rect 285312 4616 285364 4622
rect 285312 4558 285364 4564
rect 285508 4486 285536 217874
rect 285496 4480 285548 4486
rect 285496 4422 285548 4428
rect 285600 3942 285628 220102
rect 285692 217258 285720 220116
rect 285680 217252 285732 217258
rect 285680 217194 285732 217200
rect 286152 212566 286180 220116
rect 286520 217938 286548 220116
rect 286796 220102 286902 220130
rect 286508 217932 286560 217938
rect 286508 217874 286560 217880
rect 286140 212560 286192 212566
rect 286140 212502 286192 212508
rect 286600 212560 286652 212566
rect 286600 212502 286652 212508
rect 286612 205698 286640 212502
rect 286600 205692 286652 205698
rect 286600 205634 286652 205640
rect 286692 205556 286744 205562
rect 286692 205498 286744 205504
rect 286704 202881 286732 205498
rect 286506 202872 286562 202881
rect 286506 202807 286562 202816
rect 286690 202872 286746 202881
rect 286690 202807 286746 202816
rect 286520 193254 286548 202807
rect 286508 193248 286560 193254
rect 286508 193190 286560 193196
rect 286692 193248 286744 193254
rect 286692 193190 286744 193196
rect 286704 183666 286732 193190
rect 286692 183660 286744 183666
rect 286692 183602 286744 183608
rect 286600 183592 286652 183598
rect 286598 183560 286600 183569
rect 286652 183560 286654 183569
rect 286598 183495 286654 183504
rect 286506 183424 286562 183433
rect 286506 183359 286562 183368
rect 286520 173942 286548 183359
rect 286508 173936 286560 173942
rect 286508 173878 286560 173884
rect 286600 173800 286652 173806
rect 286600 173742 286652 173748
rect 286612 164218 286640 173742
rect 286600 164212 286652 164218
rect 286600 164154 286652 164160
rect 286692 164212 286744 164218
rect 286692 164154 286744 164160
rect 286704 162858 286732 164154
rect 286692 162852 286744 162858
rect 286692 162794 286744 162800
rect 286692 153264 286744 153270
rect 286692 153206 286744 153212
rect 286704 144922 286732 153206
rect 286612 144894 286732 144922
rect 286612 143546 286640 144894
rect 286600 143540 286652 143546
rect 286600 143482 286652 143488
rect 286600 137964 286652 137970
rect 286600 137906 286652 137912
rect 286612 133906 286640 137906
rect 286612 133878 286732 133906
rect 286704 125662 286732 133878
rect 286600 125656 286652 125662
rect 286600 125598 286652 125604
rect 286692 125656 286744 125662
rect 286692 125598 286744 125604
rect 286612 120714 286640 125598
rect 286612 120686 286732 120714
rect 286704 115938 286732 120686
rect 286416 115932 286468 115938
rect 286416 115874 286468 115880
rect 286692 115932 286744 115938
rect 286692 115874 286744 115880
rect 286428 106321 286456 115874
rect 286414 106312 286470 106321
rect 286414 106247 286470 106256
rect 286598 106312 286654 106321
rect 286598 106247 286654 106256
rect 286612 101402 286640 106247
rect 286612 101374 286732 101402
rect 286704 89808 286732 101374
rect 286612 89780 286732 89808
rect 286612 80730 286640 89780
rect 286520 80702 286640 80730
rect 286520 67658 286548 80702
rect 286508 67652 286560 67658
rect 286508 67594 286560 67600
rect 286600 67652 286652 67658
rect 286600 67594 286652 67600
rect 286612 66230 286640 67594
rect 286600 66224 286652 66230
rect 286600 66166 286652 66172
rect 286692 56636 286744 56642
rect 286692 56578 286744 56584
rect 286704 48346 286732 56578
rect 286600 48340 286652 48346
rect 286600 48282 286652 48288
rect 286692 48340 286744 48346
rect 286692 48282 286744 48288
rect 286612 43466 286640 48282
rect 286612 43438 286732 43466
rect 286704 31822 286732 43438
rect 286692 31816 286744 31822
rect 286692 31758 286744 31764
rect 286600 31748 286652 31754
rect 286600 31690 286652 31696
rect 286612 26330 286640 31690
rect 286612 26302 286732 26330
rect 286704 12510 286732 26302
rect 286692 12504 286744 12510
rect 286692 12446 286744 12452
rect 286600 12436 286652 12442
rect 286600 12378 286652 12384
rect 286612 4758 286640 12378
rect 286796 5438 286824 220102
rect 286968 217932 287020 217938
rect 286968 217874 287020 217880
rect 286876 217252 286928 217258
rect 286876 217194 286928 217200
rect 286784 5432 286836 5438
rect 286784 5374 286836 5380
rect 286600 4752 286652 4758
rect 286600 4694 286652 4700
rect 286888 4690 286916 217194
rect 286876 4684 286928 4690
rect 286876 4626 286928 4632
rect 286980 4146 287008 217874
rect 287348 217054 287376 220116
rect 287716 217938 287744 220116
rect 287704 217932 287756 217938
rect 287704 217874 287756 217880
rect 287336 217048 287388 217054
rect 287336 216990 287388 216996
rect 288176 5302 288204 220116
rect 288348 217932 288400 217938
rect 288348 217874 288400 217880
rect 288256 217048 288308 217054
rect 288256 216990 288308 216996
rect 288268 5506 288296 216990
rect 288256 5500 288308 5506
rect 288256 5442 288308 5448
rect 288164 5296 288216 5302
rect 288164 5238 288216 5244
rect 286968 4140 287020 4146
rect 286968 4082 287020 4088
rect 285956 4004 286008 4010
rect 285956 3946 286008 3952
rect 285588 3936 285640 3942
rect 285588 3878 285640 3884
rect 284206 3360 284262 3369
rect 284206 3295 284262 3304
rect 284760 2848 284812 2854
rect 284760 2790 284812 2796
rect 284772 400 284800 2790
rect 285968 400 285996 3946
rect 287612 3936 287664 3942
rect 287664 3884 288020 3890
rect 287612 3878 288020 3884
rect 287152 3868 287204 3874
rect 287624 3862 288020 3878
rect 287152 3810 287204 3816
rect 287164 400 287192 3810
rect 287992 3806 288020 3862
rect 287980 3800 288032 3806
rect 287980 3742 288032 3748
rect 288360 3670 288388 217874
rect 288544 217326 288572 220116
rect 288532 217320 288584 217326
rect 288532 217262 288584 217268
rect 289004 212566 289032 220116
rect 289372 217938 289400 220116
rect 289556 220102 289754 220130
rect 289360 217932 289412 217938
rect 289360 217874 289412 217880
rect 288992 212560 289044 212566
rect 289360 212560 289412 212566
rect 288992 212502 289044 212508
rect 289174 212528 289230 212537
rect 289174 212463 289230 212472
rect 289358 212528 289360 212537
rect 289412 212528 289414 212537
rect 289358 212463 289414 212472
rect 289188 202910 289216 212463
rect 289176 202904 289228 202910
rect 289452 202904 289504 202910
rect 289176 202846 289228 202852
rect 289266 202872 289322 202881
rect 289266 202807 289322 202816
rect 289450 202872 289452 202881
rect 289504 202872 289506 202881
rect 289450 202807 289506 202816
rect 289280 193254 289308 202807
rect 289268 193248 289320 193254
rect 289266 193216 289268 193225
rect 289452 193248 289504 193254
rect 289320 193216 289322 193225
rect 289266 193151 289322 193160
rect 289450 193216 289452 193225
rect 289504 193216 289506 193225
rect 289450 193151 289506 193160
rect 289280 183598 289308 193151
rect 289268 183592 289320 183598
rect 289266 183560 289268 183569
rect 289452 183592 289504 183598
rect 289320 183560 289322 183569
rect 289266 183495 289322 183504
rect 289450 183560 289452 183569
rect 289504 183560 289506 183569
rect 289450 183495 289506 183504
rect 289280 173942 289308 183495
rect 289268 173936 289320 173942
rect 289268 173878 289320 173884
rect 289452 173936 289504 173942
rect 289452 173878 289504 173884
rect 289464 166818 289492 173878
rect 289372 166790 289492 166818
rect 289372 164218 289400 166790
rect 289360 164212 289412 164218
rect 289360 164154 289412 164160
rect 289452 164212 289504 164218
rect 289452 164154 289504 164160
rect 289464 162858 289492 164154
rect 289268 162852 289320 162858
rect 289268 162794 289320 162800
rect 289452 162852 289504 162858
rect 289452 162794 289504 162800
rect 289280 153241 289308 162794
rect 289266 153232 289322 153241
rect 289266 153167 289322 153176
rect 289450 153232 289506 153241
rect 289450 153167 289506 153176
rect 289464 144922 289492 153167
rect 289372 144894 289492 144922
rect 289372 143546 289400 144894
rect 289360 143540 289412 143546
rect 289360 143482 289412 143488
rect 289360 137964 289412 137970
rect 289360 137906 289412 137912
rect 289372 133906 289400 137906
rect 289372 133878 289492 133906
rect 289464 125662 289492 133878
rect 289360 125656 289412 125662
rect 289360 125598 289412 125604
rect 289452 125656 289504 125662
rect 289452 125598 289504 125604
rect 289372 120714 289400 125598
rect 289372 120686 289492 120714
rect 289464 115938 289492 120686
rect 289176 115932 289228 115938
rect 289176 115874 289228 115880
rect 289452 115932 289504 115938
rect 289452 115874 289504 115880
rect 289188 106321 289216 115874
rect 289174 106312 289230 106321
rect 289174 106247 289230 106256
rect 289358 106312 289414 106321
rect 289358 106247 289414 106256
rect 289372 101402 289400 106247
rect 289372 101374 289492 101402
rect 289464 86986 289492 101374
rect 289372 86958 289492 86986
rect 289372 85542 289400 86958
rect 289360 85536 289412 85542
rect 289360 85478 289412 85484
rect 289268 75948 289320 75954
rect 289268 75890 289320 75896
rect 289280 67658 289308 75890
rect 289268 67652 289320 67658
rect 289268 67594 289320 67600
rect 289360 67652 289412 67658
rect 289360 67594 289412 67600
rect 289372 66230 289400 67594
rect 289360 66224 289412 66230
rect 289360 66166 289412 66172
rect 289452 56636 289504 56642
rect 289452 56578 289504 56584
rect 289464 48346 289492 56578
rect 289360 48340 289412 48346
rect 289360 48282 289412 48288
rect 289452 48340 289504 48346
rect 289452 48282 289504 48288
rect 289372 43466 289400 48282
rect 289372 43438 289492 43466
rect 289464 29034 289492 43438
rect 289268 29028 289320 29034
rect 289268 28970 289320 28976
rect 289452 29028 289504 29034
rect 289452 28970 289504 28976
rect 289280 18057 289308 28970
rect 289266 18048 289322 18057
rect 289266 17983 289322 17992
rect 289266 17912 289322 17921
rect 289266 17847 289322 17856
rect 289280 13122 289308 17847
rect 289268 13116 289320 13122
rect 289268 13058 289320 13064
rect 289556 8022 289584 220102
rect 289728 217932 289780 217938
rect 289728 217874 289780 217880
rect 289636 217320 289688 217326
rect 289636 217262 289688 217268
rect 289544 8016 289596 8022
rect 289544 7958 289596 7964
rect 289648 5370 289676 217262
rect 289636 5364 289688 5370
rect 289636 5306 289688 5312
rect 289740 5234 289768 217874
rect 290200 217326 290228 220116
rect 290568 217938 290596 220116
rect 290936 220102 291042 220130
rect 290556 217932 290608 217938
rect 290556 217874 290608 217880
rect 290188 217320 290240 217326
rect 290188 217262 290240 217268
rect 290464 216980 290516 216986
rect 290464 216922 290516 216928
rect 289910 40352 289966 40361
rect 289910 40287 289966 40296
rect 289818 40216 289874 40225
rect 289924 40202 289952 40287
rect 289874 40174 289952 40202
rect 289818 40151 289874 40160
rect 289728 5228 289780 5234
rect 289728 5170 289780 5176
rect 288348 3664 288400 3670
rect 288348 3606 288400 3612
rect 289544 2984 289596 2990
rect 289544 2926 289596 2932
rect 288348 2916 288400 2922
rect 288348 2858 288400 2864
rect 288360 400 288388 2858
rect 289556 400 289584 2926
rect 290476 2922 290504 216922
rect 290936 7954 290964 220102
rect 291396 217938 291424 220116
rect 291016 217932 291068 217938
rect 291016 217874 291068 217880
rect 291384 217932 291436 217938
rect 291384 217874 291436 217880
rect 290924 7948 290976 7954
rect 290924 7890 290976 7896
rect 291028 5166 291056 217874
rect 291108 217320 291160 217326
rect 291108 217262 291160 217268
rect 291016 5160 291068 5166
rect 291016 5102 291068 5108
rect 291120 3602 291148 217262
rect 291856 216782 291884 220116
rect 292238 220102 292344 220130
rect 291844 216776 291896 216782
rect 291844 216718 291896 216724
rect 291936 215212 291988 215218
rect 291936 215154 291988 215160
rect 291948 196058 291976 215154
rect 291856 196030 291976 196058
rect 291856 193225 291884 196030
rect 291658 193216 291714 193225
rect 291658 193151 291714 193160
rect 291842 193216 291898 193225
rect 291842 193151 291898 193160
rect 291672 183598 291700 193151
rect 291660 183592 291712 183598
rect 291660 183534 291712 183540
rect 291936 183592 291988 183598
rect 291936 183534 291988 183540
rect 291948 176798 291976 183534
rect 291936 176792 291988 176798
rect 291936 176734 291988 176740
rect 291936 176588 291988 176594
rect 291936 176530 291988 176536
rect 291948 157350 291976 176530
rect 291936 157344 291988 157350
rect 291936 157286 291988 157292
rect 291936 157208 291988 157214
rect 291936 157150 291988 157156
rect 291948 154562 291976 157150
rect 291936 154556 291988 154562
rect 291936 154498 291988 154504
rect 291936 145036 291988 145042
rect 291936 144978 291988 144984
rect 291948 143546 291976 144978
rect 291844 143540 291896 143546
rect 291844 143482 291896 143488
rect 291936 143540 291988 143546
rect 291936 143482 291988 143488
rect 291856 134065 291884 143482
rect 291842 134056 291898 134065
rect 291842 133991 291898 134000
rect 291934 133920 291990 133929
rect 291752 133884 291804 133890
rect 291934 133855 291936 133864
rect 291752 133826 291804 133832
rect 291988 133855 291990 133864
rect 291936 133826 291988 133832
rect 291764 124273 291792 133826
rect 291750 124264 291806 124273
rect 291750 124199 291806 124208
rect 291934 124264 291990 124273
rect 291934 124199 291990 124208
rect 291948 124166 291976 124199
rect 291936 124160 291988 124166
rect 291936 124102 291988 124108
rect 291936 114572 291988 114578
rect 291936 114514 291988 114520
rect 291948 99362 291976 114514
rect 291948 99334 292068 99362
rect 292040 96694 292068 99334
rect 291936 96688 291988 96694
rect 291936 96630 291988 96636
rect 292028 96688 292080 96694
rect 292028 96630 292080 96636
rect 291948 80102 291976 96630
rect 291936 80096 291988 80102
rect 291936 80038 291988 80044
rect 291844 80028 291896 80034
rect 291844 79970 291896 79976
rect 291856 77330 291884 79970
rect 291856 77302 291976 77330
rect 291948 66230 291976 77302
rect 291936 66224 291988 66230
rect 291936 66166 291988 66172
rect 292028 66156 292080 66162
rect 292028 66098 292080 66104
rect 292040 51066 292068 66098
rect 291844 51060 291896 51066
rect 291844 51002 291896 51008
rect 292028 51060 292080 51066
rect 292028 51002 292080 51008
rect 291856 48210 291884 51002
rect 291752 48204 291804 48210
rect 291752 48146 291804 48152
rect 291844 48204 291896 48210
rect 291844 48146 291896 48152
rect 291764 43330 291792 48146
rect 291764 43302 291884 43330
rect 291856 31822 291884 43302
rect 291844 31816 291896 31822
rect 291844 31758 291896 31764
rect 291936 31748 291988 31754
rect 291936 31690 291988 31696
rect 291948 22166 291976 31690
rect 291936 22160 291988 22166
rect 291936 22102 291988 22108
rect 291936 22024 291988 22030
rect 291936 21966 291988 21972
rect 291948 19310 291976 21966
rect 291936 19304 291988 19310
rect 291936 19246 291988 19252
rect 291844 9716 291896 9722
rect 291844 9658 291896 9664
rect 290740 3596 290792 3602
rect 290740 3538 290792 3544
rect 291108 3596 291160 3602
rect 291108 3538 291160 3544
rect 290464 2916 290516 2922
rect 290464 2858 290516 2864
rect 290752 400 290780 3538
rect 291856 950 291884 9658
rect 292316 7886 292344 220102
rect 292488 217932 292540 217938
rect 292488 217874 292540 217880
rect 292396 216776 292448 216782
rect 292396 216718 292448 216724
rect 292304 7880 292356 7886
rect 292304 7822 292356 7828
rect 292408 5098 292436 216718
rect 292396 5092 292448 5098
rect 292396 5034 292448 5040
rect 292500 3534 292528 217874
rect 292684 217734 292712 220116
rect 292672 217728 292724 217734
rect 292672 217670 292724 217676
rect 293052 217122 293080 220116
rect 293434 220102 293724 220130
rect 293040 217116 293092 217122
rect 293040 217058 293092 217064
rect 293696 7818 293724 220102
rect 293880 217938 293908 220116
rect 293868 217932 293920 217938
rect 293868 217874 293920 217880
rect 293868 217728 293920 217734
rect 293868 217670 293920 217676
rect 293776 217116 293828 217122
rect 293776 217058 293828 217064
rect 293684 7812 293736 7818
rect 293684 7754 293736 7760
rect 293788 5030 293816 217058
rect 293776 5024 293828 5030
rect 293776 4966 293828 4972
rect 291936 3528 291988 3534
rect 291936 3470 291988 3476
rect 292488 3528 292540 3534
rect 292488 3470 292540 3476
rect 291844 944 291896 950
rect 291844 886 291896 892
rect 291948 400 291976 3470
rect 293880 3466 293908 217670
rect 294248 217054 294276 220116
rect 294236 217048 294288 217054
rect 294236 216990 294288 216996
rect 294708 212566 294736 220116
rect 295090 220102 295196 220130
rect 294696 212560 294748 212566
rect 294696 212502 294748 212508
rect 295064 212560 295116 212566
rect 295064 212502 295116 212508
rect 295076 196058 295104 212502
rect 294984 196030 295104 196058
rect 294984 195922 295012 196030
rect 294984 195894 295104 195922
rect 295076 167090 295104 195894
rect 294984 167062 295104 167090
rect 294984 166954 295012 167062
rect 294984 166926 295104 166954
rect 295076 147778 295104 166926
rect 294984 147750 295104 147778
rect 294984 147642 295012 147750
rect 294984 147614 295104 147642
rect 295076 128466 295104 147614
rect 294984 128438 295104 128466
rect 294984 128330 295012 128438
rect 294984 128302 295104 128330
rect 295076 109154 295104 128302
rect 294984 109126 295104 109154
rect 294984 109018 295012 109126
rect 294984 108990 295104 109018
rect 295076 89842 295104 108990
rect 294984 89814 295104 89842
rect 294984 89706 295012 89814
rect 294984 89678 295104 89706
rect 295076 70394 295104 89678
rect 294984 70366 295104 70394
rect 294984 70258 295012 70366
rect 294984 70230 295104 70258
rect 295076 51082 295104 70230
rect 294984 51054 295104 51082
rect 294984 50946 295012 51054
rect 294984 50918 295104 50946
rect 295076 31770 295104 50918
rect 294984 31742 295104 31770
rect 294984 31634 295012 31742
rect 294984 31606 295104 31634
rect 295076 12458 295104 31606
rect 294984 12430 295104 12458
rect 294984 7750 295012 12430
rect 294972 7744 295024 7750
rect 294972 7686 295024 7692
rect 295168 7614 295196 220102
rect 295536 217666 295564 220116
rect 295904 217734 295932 220116
rect 296286 220102 296484 220130
rect 295892 217728 295944 217734
rect 295892 217670 295944 217676
rect 295524 217660 295576 217666
rect 295524 217602 295576 217608
rect 295248 217048 295300 217054
rect 295248 216990 295300 216996
rect 295156 7608 295208 7614
rect 295156 7550 295208 7556
rect 295260 4962 295288 216990
rect 296456 14754 296484 220102
rect 296732 217734 296760 220116
rect 296536 217728 296588 217734
rect 296536 217670 296588 217676
rect 296720 217728 296772 217734
rect 296720 217670 296772 217676
rect 296444 14748 296496 14754
rect 296444 14690 296496 14696
rect 296548 7682 296576 217670
rect 296628 217660 296680 217666
rect 296628 217602 296680 217608
rect 296536 7676 296588 7682
rect 296536 7618 296588 7624
rect 295248 4956 295300 4962
rect 295248 4898 295300 4904
rect 296640 4894 296668 217602
rect 297100 217190 297128 220116
rect 297574 220102 297772 220130
rect 297088 217184 297140 217190
rect 297088 217126 297140 217132
rect 297364 216980 297416 216986
rect 297364 216922 297416 216928
rect 296628 4888 296680 4894
rect 296628 4830 296680 4836
rect 297376 3466 297404 216922
rect 297744 14686 297772 220102
rect 297824 217184 297876 217190
rect 297824 217126 297876 217132
rect 297732 14680 297784 14686
rect 297732 14622 297784 14628
rect 297836 11286 297864 217126
rect 297824 11280 297876 11286
rect 297824 11222 297876 11228
rect 297928 4865 297956 220116
rect 298008 217728 298060 217734
rect 298008 217670 298060 217676
rect 297914 4856 297970 4865
rect 298020 4826 298048 217670
rect 298388 217122 298416 220116
rect 298770 220102 299060 220130
rect 299230 220102 299428 220130
rect 298744 217864 298796 217870
rect 298744 217806 298796 217812
rect 298376 217116 298428 217122
rect 298376 217058 298428 217064
rect 297914 4791 297970 4800
rect 298008 4820 298060 4826
rect 298008 4762 298060 4768
rect 293132 3460 293184 3466
rect 293132 3402 293184 3408
rect 293868 3460 293920 3466
rect 293868 3402 293920 3408
rect 297364 3460 297416 3466
rect 297364 3402 297416 3408
rect 293144 400 293172 3402
rect 298756 3058 298784 217806
rect 299032 217682 299060 220102
rect 299032 217654 299244 217682
rect 299216 196058 299244 217654
rect 299296 217116 299348 217122
rect 299296 217058 299348 217064
rect 299032 196030 299244 196058
rect 299032 195922 299060 196030
rect 299032 195894 299152 195922
rect 299124 180826 299152 195894
rect 299124 180798 299244 180826
rect 299216 167090 299244 180798
rect 299032 167062 299244 167090
rect 299032 166954 299060 167062
rect 299032 166926 299152 166954
rect 299124 166818 299152 166926
rect 299124 166790 299244 166818
rect 299216 147830 299244 166790
rect 299204 147824 299256 147830
rect 299204 147766 299256 147772
rect 299204 144968 299256 144974
rect 299204 144910 299256 144916
rect 299216 128518 299244 144910
rect 299204 128512 299256 128518
rect 299204 128454 299256 128460
rect 299204 124228 299256 124234
rect 299204 124170 299256 124176
rect 299216 103562 299244 124170
rect 299204 103556 299256 103562
rect 299204 103498 299256 103504
rect 299204 102264 299256 102270
rect 299204 102206 299256 102212
rect 299216 102134 299244 102206
rect 298928 102128 298980 102134
rect 298928 102070 298980 102076
rect 299204 102128 299256 102134
rect 299204 102070 299256 102076
rect 298940 87009 298968 102070
rect 298926 87000 298982 87009
rect 298926 86935 298982 86944
rect 299202 87000 299258 87009
rect 299202 86935 299258 86944
rect 299216 31770 299244 86935
rect 299124 31742 299244 31770
rect 299124 14618 299152 31742
rect 299112 14612 299164 14618
rect 299112 14554 299164 14560
rect 299308 11354 299336 217058
rect 299296 11348 299348 11354
rect 299296 11290 299348 11296
rect 299400 9926 299428 220102
rect 299584 217666 299612 220116
rect 299572 217660 299624 217666
rect 299572 217602 299624 217608
rect 299952 212566 299980 220116
rect 300412 217734 300440 220116
rect 300688 220102 300794 220130
rect 300400 217728 300452 217734
rect 300400 217670 300452 217676
rect 300584 217660 300636 217666
rect 300584 217602 300636 217608
rect 300124 217184 300176 217190
rect 300124 217126 300176 217132
rect 299940 212560 299992 212566
rect 299940 212502 299992 212508
rect 299388 9920 299440 9926
rect 299388 9862 299440 9868
rect 300136 3126 300164 217126
rect 300492 212560 300544 212566
rect 300492 212502 300544 212508
rect 300504 196058 300532 212502
rect 300320 196030 300532 196058
rect 300320 195922 300348 196030
rect 300320 195894 300440 195922
rect 300412 180826 300440 195894
rect 300412 180798 300532 180826
rect 300504 167090 300532 180798
rect 300320 167062 300532 167090
rect 300320 166954 300348 167062
rect 300320 166926 300440 166954
rect 300412 166818 300440 166926
rect 300412 166790 300532 166818
rect 300504 147830 300532 166790
rect 300492 147824 300544 147830
rect 300492 147766 300544 147772
rect 300492 144968 300544 144974
rect 300492 144910 300544 144916
rect 300504 128518 300532 144910
rect 300492 128512 300544 128518
rect 300492 128454 300544 128460
rect 300492 124228 300544 124234
rect 300492 124170 300544 124176
rect 300504 109206 300532 124170
rect 300492 109200 300544 109206
rect 300492 109142 300544 109148
rect 300492 103556 300544 103562
rect 300492 103498 300544 103504
rect 300504 31770 300532 103498
rect 300412 31742 300532 31770
rect 300412 14550 300440 31742
rect 300400 14544 300452 14550
rect 300400 14486 300452 14492
rect 300596 11422 300624 217602
rect 300688 11490 300716 220102
rect 301240 217870 301268 220116
rect 301228 217864 301280 217870
rect 301228 217806 301280 217812
rect 301608 217734 301636 220116
rect 300768 217728 300820 217734
rect 300768 217670 300820 217676
rect 301596 217728 301648 217734
rect 301596 217670 301648 217676
rect 300676 11484 300728 11490
rect 300676 11426 300728 11432
rect 300584 11416 300636 11422
rect 300584 11358 300636 11364
rect 300780 9994 300808 217670
rect 301504 217456 301556 217462
rect 301504 217398 301556 217404
rect 300768 9988 300820 9994
rect 300768 9930 300820 9936
rect 301412 3460 301464 3466
rect 301412 3402 301464 3408
rect 300308 3188 300360 3194
rect 300308 3130 300360 3136
rect 299112 3120 299164 3126
rect 299112 3062 299164 3068
rect 300124 3120 300176 3126
rect 300124 3062 300176 3068
rect 295524 3052 295576 3058
rect 295524 2994 295576 3000
rect 298744 3052 298796 3058
rect 298744 2994 298796 3000
rect 294328 2848 294380 2854
rect 294328 2790 294380 2796
rect 294340 400 294368 2790
rect 295536 400 295564 2994
rect 297916 2916 297968 2922
rect 297916 2858 297968 2864
rect 296720 944 296772 950
rect 296720 886 296772 892
rect 296732 400 296760 886
rect 297928 400 297956 2858
rect 299124 400 299152 3062
rect 300320 400 300348 3130
rect 301424 400 301452 3402
rect 301516 3194 301544 217398
rect 302068 11558 302096 220116
rect 302148 217728 302200 217734
rect 302148 217670 302200 217676
rect 302056 11552 302108 11558
rect 302056 11494 302108 11500
rect 302160 10062 302188 217670
rect 302436 217054 302464 220116
rect 302424 217048 302476 217054
rect 302424 216990 302476 216996
rect 302804 216782 302832 220116
rect 303278 220102 303476 220130
rect 302884 217660 302936 217666
rect 302884 217602 302936 217608
rect 302792 216776 302844 216782
rect 302792 216718 302844 216724
rect 302148 10056 302200 10062
rect 302148 9998 302200 10004
rect 301504 3188 301556 3194
rect 301504 3130 301556 3136
rect 302608 3052 302660 3058
rect 302608 2994 302660 3000
rect 302620 400 302648 2994
rect 302896 2854 302924 217602
rect 302976 217388 303028 217394
rect 302976 217330 303028 217336
rect 302988 3262 303016 217330
rect 303448 11626 303476 220102
rect 303632 217734 303660 220116
rect 303620 217728 303672 217734
rect 303620 217670 303672 217676
rect 304092 216782 304120 220116
rect 304474 220102 304856 220130
rect 304264 217796 304316 217802
rect 304264 217738 304316 217744
rect 303528 216776 303580 216782
rect 303528 216718 303580 216724
rect 304080 216776 304132 216782
rect 304080 216718 304132 216724
rect 303436 11620 303488 11626
rect 303436 11562 303488 11568
rect 303540 10130 303568 216718
rect 303528 10124 303580 10130
rect 303528 10066 303580 10072
rect 302976 3256 303028 3262
rect 302976 3198 303028 3204
rect 303804 2984 303856 2990
rect 303804 2926 303856 2932
rect 302884 2848 302936 2854
rect 302884 2790 302936 2796
rect 303816 400 303844 2926
rect 304276 2922 304304 217738
rect 304828 11694 304856 220102
rect 304920 216918 304948 220116
rect 304908 216912 304960 216918
rect 304908 216854 304960 216860
rect 305288 216782 305316 220116
rect 305670 220102 306052 220130
rect 305736 217252 305788 217258
rect 305736 217194 305788 217200
rect 305644 216980 305696 216986
rect 305644 216922 305696 216928
rect 304908 216776 304960 216782
rect 304908 216718 304960 216724
rect 305276 216776 305328 216782
rect 305276 216718 305328 216724
rect 304816 11688 304868 11694
rect 304816 11630 304868 11636
rect 304920 10198 304948 216718
rect 304908 10192 304960 10198
rect 304908 10134 304960 10140
rect 305656 3126 305684 216922
rect 305000 3120 305052 3126
rect 305000 3062 305052 3068
rect 305644 3120 305696 3126
rect 305644 3062 305696 3068
rect 304264 2916 304316 2922
rect 304264 2858 304316 2864
rect 305012 400 305040 3062
rect 305748 2990 305776 217194
rect 306024 216866 306052 220102
rect 306116 217462 306144 220116
rect 306104 217456 306156 217462
rect 306104 217398 306156 217404
rect 306024 216838 306328 216866
rect 306196 216776 306248 216782
rect 306196 216718 306248 216724
rect 306208 10266 306236 216718
rect 306196 10260 306248 10266
rect 306196 10202 306248 10208
rect 306300 8362 306328 216838
rect 306484 216782 306512 220116
rect 306472 216776 306524 216782
rect 306472 216718 306524 216724
rect 306944 216714 306972 220116
rect 307312 217054 307340 220116
rect 307300 217048 307352 217054
rect 307300 216990 307352 216996
rect 307772 216782 307800 220116
rect 307576 216776 307628 216782
rect 307576 216718 307628 216724
rect 307760 216776 307812 216782
rect 307760 216718 307812 216724
rect 306932 216708 306984 216714
rect 306932 216650 306984 216656
rect 307588 11014 307616 216718
rect 308140 216714 308168 220116
rect 308404 218000 308456 218006
rect 308404 217942 308456 217948
rect 307668 216708 307720 216714
rect 307668 216650 307720 216656
rect 308128 216708 308180 216714
rect 308128 216650 308180 216656
rect 307576 11008 307628 11014
rect 307576 10950 307628 10956
rect 307680 8430 307708 216650
rect 307668 8424 307720 8430
rect 307668 8366 307720 8372
rect 306288 8356 306340 8362
rect 306288 8298 306340 8304
rect 306378 4176 306434 4185
rect 306378 4111 306380 4120
rect 306432 4111 306434 4120
rect 306380 4082 306432 4088
rect 307392 3324 307444 3330
rect 307392 3266 307444 3272
rect 306196 3256 306248 3262
rect 306196 3198 306248 3204
rect 305736 2984 305788 2990
rect 305736 2926 305788 2932
rect 306208 400 306236 3198
rect 307404 400 307432 3266
rect 308416 3126 308444 217942
rect 308600 216986 308628 220116
rect 308982 220102 309088 220130
rect 308588 216980 308640 216986
rect 308588 216922 308640 216928
rect 308864 216776 308916 216782
rect 308864 216718 308916 216724
rect 308876 10946 308904 216718
rect 308956 216708 309008 216714
rect 308956 216650 309008 216656
rect 308864 10940 308916 10946
rect 308864 10882 308916 10888
rect 308968 8498 308996 216650
rect 308956 8492 309008 8498
rect 308956 8434 309008 8440
rect 309060 5574 309088 220102
rect 309336 216714 309364 220116
rect 309810 220102 310100 220130
rect 310178 220102 310468 220130
rect 309784 217524 309836 217530
rect 309784 217466 309836 217472
rect 309324 216708 309376 216714
rect 309324 216650 309376 216656
rect 309796 6882 309824 217466
rect 310072 217190 310100 220102
rect 310060 217184 310112 217190
rect 310060 217126 310112 217132
rect 310336 216708 310388 216714
rect 310336 216650 310388 216656
rect 310348 8566 310376 216650
rect 310336 8560 310388 8566
rect 310336 8502 310388 8508
rect 309704 6854 309824 6882
rect 309048 5568 309100 5574
rect 309048 5510 309100 5516
rect 309704 3330 309732 6854
rect 310440 5642 310468 220102
rect 310624 216714 310652 220116
rect 310992 217394 311020 220116
rect 310980 217388 311032 217394
rect 310980 217330 311032 217336
rect 311452 216782 311480 220116
rect 311728 220102 311834 220130
rect 311440 216776 311492 216782
rect 311440 216718 311492 216724
rect 310612 216708 310664 216714
rect 310612 216650 310664 216656
rect 311624 216708 311676 216714
rect 311624 216650 311676 216656
rect 311636 8634 311664 216650
rect 311728 8702 311756 220102
rect 312188 217054 312216 220116
rect 312544 217320 312596 217326
rect 312544 217262 312596 217268
rect 312176 217048 312228 217054
rect 312176 216990 312228 216996
rect 311808 216776 311860 216782
rect 311808 216718 311860 216724
rect 311716 8696 311768 8702
rect 311716 8638 311768 8644
rect 311624 8628 311676 8634
rect 311624 8570 311676 8576
rect 311820 5710 311848 216718
rect 311808 5704 311860 5710
rect 311808 5646 311860 5652
rect 310428 5636 310480 5642
rect 310428 5578 310480 5584
rect 311070 4176 311126 4185
rect 311070 4111 311126 4120
rect 311084 4078 311112 4111
rect 310980 4072 311032 4078
rect 310980 4014 311032 4020
rect 311072 4072 311124 4078
rect 311072 4014 311124 4020
rect 309784 3392 309836 3398
rect 309784 3334 309836 3340
rect 309692 3324 309744 3330
rect 309692 3266 309744 3272
rect 308404 3120 308456 3126
rect 308404 3062 308456 3068
rect 308588 3052 308640 3058
rect 308588 2994 308640 3000
rect 308600 400 308628 2994
rect 309796 400 309824 3334
rect 310992 400 311020 4014
rect 312556 3398 312584 217262
rect 312648 216714 312676 220116
rect 313030 220102 313136 220130
rect 312636 216708 312688 216714
rect 312636 216650 312688 216656
rect 313108 8770 313136 220102
rect 313476 217394 313504 220116
rect 313464 217388 313516 217394
rect 313464 217330 313516 217336
rect 313844 217258 313872 220116
rect 314318 220102 314516 220130
rect 313832 217252 313884 217258
rect 313832 217194 313884 217200
rect 313188 216708 313240 216714
rect 313188 216650 313240 216656
rect 313096 8764 313148 8770
rect 313096 8706 313148 8712
rect 313200 5778 313228 216650
rect 314488 8838 314516 220102
rect 314568 217252 314620 217258
rect 314568 217194 314620 217200
rect 314476 8832 314528 8838
rect 314476 8774 314528 8780
rect 314580 5846 314608 217194
rect 314672 217138 314700 220116
rect 314844 217184 314896 217190
rect 314672 217132 314844 217138
rect 314672 217126 314896 217132
rect 314672 217110 314884 217126
rect 315132 216714 315160 220116
rect 315514 220102 315804 220130
rect 315776 219434 315804 220102
rect 315764 219428 315816 219434
rect 315764 219370 315816 219376
rect 315868 218006 315896 220116
rect 315948 219428 316000 219434
rect 315948 219370 316000 219376
rect 315856 218000 315908 218006
rect 315856 217942 315908 217948
rect 315960 217818 315988 219370
rect 315868 217790 315988 217818
rect 315120 216708 315172 216714
rect 315120 216650 315172 216656
rect 315868 205698 315896 217790
rect 316328 216714 316356 220116
rect 316710 220102 317092 220130
rect 316684 217116 316736 217122
rect 316684 217058 316736 217064
rect 315948 216708 316000 216714
rect 315948 216650 316000 216656
rect 316316 216708 316368 216714
rect 316316 216650 316368 216656
rect 315856 205692 315908 205698
rect 315856 205634 315908 205640
rect 315856 202904 315908 202910
rect 315856 202846 315908 202852
rect 315868 196110 315896 202846
rect 315856 196104 315908 196110
rect 315856 196046 315908 196052
rect 315764 191888 315816 191894
rect 315764 191830 315816 191836
rect 315776 191758 315804 191830
rect 315764 191752 315816 191758
rect 315764 191694 315816 191700
rect 315672 182232 315724 182238
rect 315672 182174 315724 182180
rect 315684 174026 315712 182174
rect 315592 173998 315712 174026
rect 315592 173754 315620 173998
rect 315592 173726 315712 173754
rect 315684 164286 315712 173726
rect 315672 164280 315724 164286
rect 315672 164222 315724 164228
rect 315764 164280 315816 164286
rect 315764 164222 315816 164228
rect 315776 157570 315804 164222
rect 315776 157542 315896 157570
rect 315868 153338 315896 157542
rect 315764 153332 315816 153338
rect 315764 153274 315816 153280
rect 315856 153332 315908 153338
rect 315856 153274 315908 153280
rect 315776 147762 315804 153274
rect 315764 147756 315816 147762
rect 315764 147698 315816 147704
rect 315764 147620 315816 147626
rect 315764 147562 315816 147568
rect 315776 143562 315804 147562
rect 315776 143534 315896 143562
rect 315868 142118 315896 143534
rect 315856 142112 315908 142118
rect 315856 142054 315908 142060
rect 315856 132524 315908 132530
rect 315856 132466 315908 132472
rect 315868 118794 315896 132466
rect 315856 118788 315908 118794
rect 315856 118730 315908 118736
rect 315856 114572 315908 114578
rect 315856 114514 315908 114520
rect 315868 109138 315896 114514
rect 315856 109132 315908 109138
rect 315856 109074 315908 109080
rect 315856 104916 315908 104922
rect 315856 104858 315908 104864
rect 315868 104802 315896 104858
rect 315776 104774 315896 104802
rect 315776 96966 315804 104774
rect 315764 96960 315816 96966
rect 315764 96902 315816 96908
rect 315764 87032 315816 87038
rect 315764 86974 315816 86980
rect 315776 58002 315804 86974
rect 315764 57996 315816 58002
rect 315764 57938 315816 57944
rect 315856 57996 315908 58002
rect 315856 57938 315908 57944
rect 315868 22114 315896 57938
rect 315776 22086 315896 22114
rect 315776 21978 315804 22086
rect 315776 21950 315896 21978
rect 315868 8906 315896 21950
rect 315856 8900 315908 8906
rect 315856 8842 315908 8848
rect 315960 5914 315988 216650
rect 315948 5908 316000 5914
rect 315948 5850 316000 5856
rect 314568 5840 314620 5846
rect 314568 5782 314620 5788
rect 313188 5772 313240 5778
rect 313188 5714 313240 5720
rect 316696 4010 316724 217058
rect 317064 217002 317092 220102
rect 317156 217530 317184 220116
rect 317144 217524 317196 217530
rect 317144 217466 317196 217472
rect 317064 216974 317276 217002
rect 317248 205714 317276 216974
rect 317524 216714 317552 220116
rect 317998 220102 318196 220130
rect 318168 217054 318196 220102
rect 318352 217802 318380 220116
rect 318340 217796 318392 217802
rect 318340 217738 318392 217744
rect 318156 217048 318208 217054
rect 318156 216990 318208 216996
rect 318524 217048 318576 217054
rect 318524 216990 318576 216996
rect 317328 216708 317380 216714
rect 317328 216650 317380 216656
rect 317512 216708 317564 216714
rect 317512 216650 317564 216656
rect 317064 205686 317276 205714
rect 317064 205578 317092 205686
rect 317064 205550 317184 205578
rect 317156 186402 317184 205550
rect 317064 186374 317184 186402
rect 317064 186266 317092 186374
rect 317064 186238 317276 186266
rect 317248 173913 317276 186238
rect 317050 173904 317106 173913
rect 317050 173839 317106 173848
rect 317234 173904 317290 173913
rect 317234 173839 317290 173848
rect 317064 167074 317092 173839
rect 317052 167068 317104 167074
rect 317052 167010 317104 167016
rect 317144 167000 317196 167006
rect 317144 166942 317196 166948
rect 317156 162858 317184 166942
rect 317144 162852 317196 162858
rect 317144 162794 317196 162800
rect 317144 157344 317196 157350
rect 317144 157286 317196 157292
rect 317156 153218 317184 157286
rect 317156 153190 317276 153218
rect 317248 147694 317276 153190
rect 317236 147688 317288 147694
rect 317236 147630 317288 147636
rect 317236 143608 317288 143614
rect 317236 143550 317288 143556
rect 317248 135250 317276 143550
rect 317144 135244 317196 135250
rect 317144 135186 317196 135192
rect 317236 135244 317288 135250
rect 317236 135186 317288 135192
rect 317156 128364 317184 135186
rect 317156 128336 317276 128364
rect 317248 109750 317276 128336
rect 317236 109744 317288 109750
rect 317236 109686 317288 109692
rect 317236 96688 317288 96694
rect 317236 96630 317288 96636
rect 317248 67658 317276 96630
rect 317052 67652 317104 67658
rect 317052 67594 317104 67600
rect 317236 67652 317288 67658
rect 317236 67594 317288 67600
rect 317064 67561 317092 67594
rect 316866 67552 316922 67561
rect 316866 67487 316922 67496
rect 317050 67552 317106 67561
rect 317050 67487 317106 67496
rect 316880 58041 316908 67487
rect 316866 58032 316922 58041
rect 316866 57967 316922 57976
rect 317050 57896 317106 57905
rect 317050 57831 317106 57840
rect 317064 50946 317092 57831
rect 317064 50918 317184 50946
rect 317156 46918 317184 50918
rect 317144 46912 317196 46918
rect 317144 46854 317196 46860
rect 317236 37324 317288 37330
rect 317236 37266 317288 37272
rect 317248 29034 317276 37266
rect 317144 29028 317196 29034
rect 317144 28970 317196 28976
rect 317236 29028 317288 29034
rect 317236 28970 317288 28976
rect 317156 28898 317184 28970
rect 317144 28892 317196 28898
rect 317144 28834 317196 28840
rect 317236 19372 317288 19378
rect 317236 19314 317288 19320
rect 317248 12594 317276 19314
rect 317156 12566 317276 12594
rect 317156 12458 317184 12566
rect 317064 12430 317184 12458
rect 317064 9654 317092 12430
rect 317052 9648 317104 9654
rect 317052 9590 317104 9596
rect 317340 5982 317368 216650
rect 318536 205714 318564 216990
rect 318616 216708 318668 216714
rect 318616 216650 318668 216656
rect 318352 205686 318564 205714
rect 318352 205578 318380 205686
rect 318352 205550 318472 205578
rect 318444 186402 318472 205550
rect 318352 186374 318472 186402
rect 318352 186266 318380 186374
rect 318352 186238 318564 186266
rect 318536 169182 318564 186238
rect 318524 169176 318576 169182
rect 318524 169118 318576 169124
rect 318432 164280 318484 164286
rect 318432 164222 318484 164228
rect 318444 162858 318472 164222
rect 318432 162852 318484 162858
rect 318432 162794 318484 162800
rect 318432 157344 318484 157350
rect 318432 157286 318484 157292
rect 318444 153218 318472 157286
rect 318444 153190 318564 153218
rect 318536 147801 318564 153190
rect 318522 147792 318578 147801
rect 318522 147727 318578 147736
rect 318522 143576 318578 143585
rect 318522 143511 318524 143520
rect 318576 143511 318578 143520
rect 318524 143482 318576 143488
rect 318432 134020 318484 134026
rect 318432 133962 318484 133968
rect 318444 133890 318472 133962
rect 318432 133884 318484 133890
rect 318432 133826 318484 133832
rect 318432 125588 318484 125594
rect 318432 125530 318484 125536
rect 318444 124250 318472 125530
rect 318444 124222 318564 124250
rect 318536 124166 318564 124222
rect 318524 124160 318576 124166
rect 318524 124102 318576 124108
rect 318524 114572 318576 114578
rect 318524 114514 318576 114520
rect 318536 109410 318564 114514
rect 318524 109404 318576 109410
rect 318524 109346 318576 109352
rect 318340 104916 318392 104922
rect 318340 104858 318392 104864
rect 318352 96665 318380 104858
rect 318338 96656 318394 96665
rect 318338 96591 318394 96600
rect 318522 96656 318578 96665
rect 318522 96591 318578 96600
rect 318536 77586 318564 96591
rect 318524 77580 318576 77586
rect 318524 77522 318576 77528
rect 318248 75948 318300 75954
rect 318248 75890 318300 75896
rect 318260 70258 318288 75890
rect 318260 70230 318380 70258
rect 318352 67561 318380 70230
rect 318338 67552 318394 67561
rect 318338 67487 318394 67496
rect 318522 67416 318578 67425
rect 318522 67351 318578 67360
rect 318536 57934 318564 67351
rect 318340 57928 318392 57934
rect 318340 57870 318392 57876
rect 318524 57928 318576 57934
rect 318524 57870 318576 57876
rect 318352 56574 318380 57870
rect 318340 56568 318392 56574
rect 318340 56510 318392 56516
rect 318432 46980 318484 46986
rect 318432 46922 318484 46928
rect 318444 46889 318472 46922
rect 318430 46880 318486 46889
rect 318430 46815 318486 46824
rect 318338 46744 318394 46753
rect 318338 46679 318394 46688
rect 318352 41290 318380 46679
rect 318352 41262 318472 41290
rect 318444 33862 318472 41262
rect 318432 33856 318484 33862
rect 318432 33798 318484 33804
rect 318524 33788 318576 33794
rect 318524 33730 318576 33736
rect 318536 12594 318564 33730
rect 318444 12566 318564 12594
rect 318444 12458 318472 12566
rect 318352 12430 318472 12458
rect 318352 9586 318380 12430
rect 318340 9580 318392 9586
rect 318340 9522 318392 9528
rect 318628 6050 318656 216650
rect 318720 6118 318748 220116
rect 319180 216714 319208 220116
rect 319444 217932 319496 217938
rect 319444 217874 319496 217880
rect 319168 216708 319220 216714
rect 319168 216650 319220 216656
rect 318708 6112 318760 6118
rect 318708 6054 318760 6060
rect 318616 6044 318668 6050
rect 318616 5986 318668 5992
rect 317328 5976 317380 5982
rect 317328 5918 317380 5924
rect 316960 4072 317012 4078
rect 316960 4014 317012 4020
rect 314568 4004 314620 4010
rect 314568 3946 314620 3952
rect 316684 4004 316736 4010
rect 316684 3946 316736 3952
rect 312544 3392 312596 3398
rect 312544 3334 312596 3340
rect 313372 3392 313424 3398
rect 313372 3334 313424 3340
rect 312176 2848 312228 2854
rect 312176 2790 312228 2796
rect 312188 400 312216 2790
rect 313384 400 313412 3334
rect 314580 400 314608 3946
rect 315764 2916 315816 2922
rect 315764 2858 315816 2864
rect 315776 400 315804 2858
rect 316972 400 317000 4014
rect 318064 3936 318116 3942
rect 318064 3878 318116 3884
rect 318076 400 318104 3878
rect 319456 3058 319484 217874
rect 319548 217666 319576 220116
rect 320022 220102 320128 220130
rect 319536 217660 319588 217666
rect 319536 217602 319588 217608
rect 319996 216708 320048 216714
rect 319996 216650 320048 216656
rect 320008 9518 320036 216650
rect 319996 9512 320048 9518
rect 319996 9454 320048 9460
rect 320100 6866 320128 220102
rect 320376 216714 320404 220116
rect 320836 217938 320864 220116
rect 321218 220102 321508 220130
rect 320824 217932 320876 217938
rect 320824 217874 320876 217880
rect 320364 216708 320416 216714
rect 320364 216650 320416 216656
rect 321376 216708 321428 216714
rect 321376 216650 321428 216656
rect 321388 9450 321416 216650
rect 321376 9444 321428 9450
rect 321376 9386 321428 9392
rect 320088 6860 320140 6866
rect 320088 6802 320140 6808
rect 321480 6798 321508 220102
rect 321664 217938 321692 220116
rect 321652 217932 321704 217938
rect 321652 217874 321704 217880
rect 322032 216782 322060 220116
rect 322400 217598 322428 220116
rect 322768 220102 322874 220130
rect 322664 217932 322716 217938
rect 322664 217874 322716 217880
rect 322388 217592 322440 217598
rect 322388 217534 322440 217540
rect 322204 217456 322256 217462
rect 322204 217398 322256 217404
rect 322020 216776 322072 216782
rect 322020 216718 322072 216724
rect 321468 6792 321520 6798
rect 321468 6734 321520 6740
rect 320456 4208 320508 4214
rect 320456 4150 320508 4156
rect 319444 3052 319496 3058
rect 319444 2994 319496 3000
rect 319260 2984 319312 2990
rect 319260 2926 319312 2932
rect 319272 400 319300 2926
rect 320468 400 320496 4150
rect 321652 3868 321704 3874
rect 321652 3810 321704 3816
rect 321664 400 321692 3810
rect 322216 2990 322244 217398
rect 322676 9382 322704 217874
rect 322664 9376 322716 9382
rect 322664 9318 322716 9324
rect 322768 9314 322796 220102
rect 322848 217592 322900 217598
rect 322848 217534 322900 217540
rect 322756 9308 322808 9314
rect 322756 9250 322808 9256
rect 322860 6730 322888 217534
rect 323228 217462 323256 220116
rect 323688 217530 323716 220116
rect 324070 220102 324176 220130
rect 323676 217524 323728 217530
rect 323676 217466 323728 217472
rect 323216 217456 323268 217462
rect 323216 217398 323268 217404
rect 323584 216708 323636 216714
rect 323584 216650 323636 216656
rect 322848 6724 322900 6730
rect 322848 6666 322900 6672
rect 322848 3256 322900 3262
rect 322848 3198 322900 3204
rect 322204 2984 322256 2990
rect 322204 2926 322256 2932
rect 322860 400 322888 3198
rect 323596 3126 323624 216650
rect 324148 9246 324176 220102
rect 324516 217530 324544 220116
rect 324884 217598 324912 220116
rect 325266 220102 325556 220130
rect 324872 217592 324924 217598
rect 324872 217534 324924 217540
rect 324228 217524 324280 217530
rect 324228 217466 324280 217472
rect 324504 217524 324556 217530
rect 324504 217466 324556 217472
rect 324136 9240 324188 9246
rect 324136 9182 324188 9188
rect 324240 6662 324268 217466
rect 325528 9178 325556 220102
rect 325608 217592 325660 217598
rect 325608 217534 325660 217540
rect 325516 9172 325568 9178
rect 325516 9114 325568 9120
rect 324228 6656 324280 6662
rect 324228 6598 324280 6604
rect 325620 6594 325648 217534
rect 325712 216714 325740 220116
rect 326080 217598 326108 220116
rect 326554 220102 326660 220130
rect 326068 217592 326120 217598
rect 326068 217534 326120 217540
rect 326344 217320 326396 217326
rect 326344 217262 326396 217268
rect 325700 216708 325752 216714
rect 325700 216650 325752 216656
rect 325608 6588 325660 6594
rect 325608 6530 325660 6536
rect 324044 4276 324096 4282
rect 324044 4218 324096 4224
rect 323584 3120 323636 3126
rect 323584 3062 323636 3068
rect 324056 400 324084 4218
rect 325240 3392 325292 3398
rect 325240 3334 325292 3340
rect 325252 400 325280 3334
rect 326356 3194 326384 217262
rect 326632 217138 326660 220102
rect 326908 217326 326936 220116
rect 327368 217598 327396 220116
rect 327750 220102 328132 220130
rect 326988 217592 327040 217598
rect 326988 217534 327040 217540
rect 327356 217592 327408 217598
rect 327356 217534 327408 217540
rect 326896 217320 326948 217326
rect 326896 217262 326948 217268
rect 326632 217110 326936 217138
rect 326908 196058 326936 217110
rect 326816 196030 326936 196058
rect 326816 195922 326844 196030
rect 326816 195894 326936 195922
rect 326908 167090 326936 195894
rect 326816 167062 326936 167090
rect 326816 166954 326844 167062
rect 326816 166926 326936 166954
rect 326908 147778 326936 166926
rect 326816 147750 326936 147778
rect 326816 147642 326844 147750
rect 326816 147614 326936 147642
rect 326908 128466 326936 147614
rect 326816 128438 326936 128466
rect 326816 128330 326844 128438
rect 326816 128302 326936 128330
rect 326908 109154 326936 128302
rect 326816 109126 326936 109154
rect 326816 109018 326844 109126
rect 326816 108990 326936 109018
rect 326908 89842 326936 108990
rect 326816 89814 326936 89842
rect 326816 89706 326844 89814
rect 326816 89678 326936 89706
rect 326908 70394 326936 89678
rect 326816 70366 326936 70394
rect 326816 70258 326844 70366
rect 326816 70230 326936 70258
rect 326908 51082 326936 70230
rect 326816 51054 326936 51082
rect 326816 50946 326844 51054
rect 326816 50918 326936 50946
rect 326908 31770 326936 50918
rect 326816 31742 326936 31770
rect 326816 31634 326844 31742
rect 326816 31606 326936 31634
rect 326908 12458 326936 31606
rect 326816 12430 326936 12458
rect 326816 9110 326844 12430
rect 326804 9104 326856 9110
rect 326804 9046 326856 9052
rect 327000 6526 327028 217534
rect 327724 217388 327776 217394
rect 327724 217330 327776 217336
rect 326988 6520 327040 6526
rect 326988 6462 327040 6468
rect 327632 4344 327684 4350
rect 327632 4286 327684 4292
rect 326436 3324 326488 3330
rect 326436 3266 326488 3272
rect 326344 3188 326396 3194
rect 326344 3130 326396 3136
rect 326448 400 326476 3266
rect 327644 400 327672 4286
rect 327736 3330 327764 217330
rect 328104 211138 328132 220102
rect 328196 217394 328224 220116
rect 328564 217598 328592 220116
rect 328946 220102 329236 220130
rect 329208 217682 329236 220102
rect 329392 217938 329420 220116
rect 329380 217932 329432 217938
rect 329380 217874 329432 217880
rect 329208 217654 329420 217682
rect 328368 217592 328420 217598
rect 328368 217534 328420 217540
rect 328552 217592 328604 217598
rect 328552 217534 328604 217540
rect 328184 217388 328236 217394
rect 328184 217330 328236 217336
rect 328092 211132 328144 211138
rect 328092 211074 328144 211080
rect 328184 205624 328236 205630
rect 328184 205566 328236 205572
rect 328196 201498 328224 205566
rect 328196 201470 328316 201498
rect 328288 193118 328316 201470
rect 328276 193112 328328 193118
rect 328276 193054 328328 193060
rect 328184 186312 328236 186318
rect 328184 186254 328236 186260
rect 328196 178786 328224 186254
rect 328104 178758 328224 178786
rect 328104 174049 328132 178758
rect 328090 174040 328146 174049
rect 328090 173975 328146 173984
rect 328274 174040 328330 174049
rect 328274 173975 328330 173984
rect 328288 173890 328316 173975
rect 328196 173862 328316 173890
rect 328196 169114 328224 173862
rect 328000 169108 328052 169114
rect 328000 169050 328052 169056
rect 328184 169108 328236 169114
rect 328184 169050 328236 169056
rect 328012 164257 328040 169050
rect 327998 164248 328054 164257
rect 327998 164183 328054 164192
rect 328182 164248 328238 164257
rect 328182 164183 328238 164192
rect 328196 157418 328224 164183
rect 328184 157412 328236 157418
rect 328184 157354 328236 157360
rect 328276 157276 328328 157282
rect 328276 157218 328328 157224
rect 328288 147694 328316 157218
rect 328276 147688 328328 147694
rect 328276 147630 328328 147636
rect 328276 144968 328328 144974
rect 328276 144910 328328 144916
rect 328288 128382 328316 144910
rect 328276 128376 328328 128382
rect 328276 128318 328328 128324
rect 328276 124228 328328 124234
rect 328276 124170 328328 124176
rect 328288 124114 328316 124170
rect 328196 124086 328316 124114
rect 328196 114578 328224 124086
rect 328184 114572 328236 114578
rect 328184 114514 328236 114520
rect 328276 114572 328328 114578
rect 328276 114514 328328 114520
rect 328288 109070 328316 114514
rect 328276 109064 328328 109070
rect 328276 109006 328328 109012
rect 328276 108928 328328 108934
rect 328276 108870 328328 108876
rect 328288 58154 328316 108870
rect 328196 58126 328316 58154
rect 328196 58002 328224 58126
rect 328184 57996 328236 58002
rect 328184 57938 328236 57944
rect 328276 57996 328328 58002
rect 328276 57938 328328 57944
rect 328288 53174 328316 57938
rect 327908 53168 327960 53174
rect 327908 53110 327960 53116
rect 328276 53168 328328 53174
rect 328276 53110 328328 53116
rect 327920 48385 327948 53110
rect 327906 48376 327962 48385
rect 327906 48311 327962 48320
rect 328090 48376 328146 48385
rect 328146 48334 328224 48362
rect 328090 48311 328146 48320
rect 328196 42106 328224 48334
rect 328196 42078 328316 42106
rect 328288 37466 328316 42078
rect 328276 37460 328328 37466
rect 328276 37402 328328 37408
rect 328276 37324 328328 37330
rect 328276 37266 328328 37272
rect 328288 37210 328316 37266
rect 328196 37182 328316 37210
rect 328196 31822 328224 37182
rect 328184 31816 328236 31822
rect 328184 31758 328236 31764
rect 328092 27668 328144 27674
rect 328092 27610 328144 27616
rect 328104 21978 328132 27610
rect 328104 21950 328316 21978
rect 328288 19310 328316 21950
rect 328276 19304 328328 19310
rect 328276 19246 328328 19252
rect 328184 9716 328236 9722
rect 328184 9658 328236 9664
rect 328196 9042 328224 9658
rect 328184 9036 328236 9042
rect 328184 8978 328236 8984
rect 328380 6458 328408 217534
rect 329392 209778 329420 217654
rect 329656 217592 329708 217598
rect 329656 217534 329708 217540
rect 329380 209772 329432 209778
rect 329380 209714 329432 209720
rect 329472 201476 329524 201482
rect 329472 201418 329524 201424
rect 329484 200138 329512 201418
rect 329484 200110 329604 200138
rect 329576 191826 329604 200110
rect 329564 191820 329616 191826
rect 329564 191762 329616 191768
rect 329380 181620 329432 181626
rect 329380 181562 329432 181568
rect 329392 173942 329420 181562
rect 329380 173936 329432 173942
rect 329564 173936 329616 173942
rect 329380 173878 329432 173884
rect 329484 173884 329564 173890
rect 329484 173878 329616 173884
rect 329484 173862 329604 173878
rect 329484 169114 329512 173862
rect 329288 169108 329340 169114
rect 329288 169050 329340 169056
rect 329472 169108 329524 169114
rect 329472 169050 329524 169056
rect 329300 164257 329328 169050
rect 329286 164248 329342 164257
rect 329286 164183 329342 164192
rect 329470 164248 329526 164257
rect 329470 164183 329526 164192
rect 329484 157418 329512 164183
rect 329472 157412 329524 157418
rect 329472 157354 329524 157360
rect 329564 157276 329616 157282
rect 329564 157218 329616 157224
rect 329576 147801 329604 157218
rect 329562 147792 329618 147801
rect 329562 147727 329618 147736
rect 329562 144936 329618 144945
rect 329562 144871 329564 144880
rect 329616 144871 329618 144880
rect 329564 144842 329616 144848
rect 329564 135312 329616 135318
rect 329564 135254 329616 135260
rect 329576 128489 329604 135254
rect 329562 128480 329618 128489
rect 329562 128415 329618 128424
rect 329562 125624 329618 125633
rect 329562 125559 329564 125568
rect 329616 125559 329618 125568
rect 329564 125530 329616 125536
rect 329564 116000 329616 116006
rect 329564 115942 329616 115948
rect 329576 109177 329604 115942
rect 329562 109168 329618 109177
rect 329562 109103 329618 109112
rect 329562 106312 329618 106321
rect 329562 106247 329564 106256
rect 329616 106247 329618 106256
rect 329564 106218 329616 106224
rect 329564 96688 329616 96694
rect 329564 96630 329616 96636
rect 329576 67794 329604 96630
rect 329564 67788 329616 67794
rect 329564 67730 329616 67736
rect 329564 67652 329616 67658
rect 329564 67594 329616 67600
rect 329576 66230 329604 67594
rect 329564 66224 329616 66230
rect 329564 66166 329616 66172
rect 329564 56636 329616 56642
rect 329564 56578 329616 56584
rect 329576 51241 329604 56578
rect 329562 51232 329618 51241
rect 329562 51167 329618 51176
rect 329470 48376 329526 48385
rect 329470 48311 329526 48320
rect 329484 42158 329512 48311
rect 329472 42152 329524 42158
rect 329472 42094 329524 42100
rect 329380 37324 329432 37330
rect 329380 37266 329432 37272
rect 329392 29050 329420 37266
rect 329392 29022 329512 29050
rect 329484 28966 329512 29022
rect 329472 28960 329524 28966
rect 329472 28902 329524 28908
rect 329564 19372 329616 19378
rect 329564 19314 329616 19320
rect 329576 19258 329604 19314
rect 329484 19230 329604 19258
rect 329484 12510 329512 19230
rect 329472 12504 329524 12510
rect 329472 12446 329524 12452
rect 329472 9716 329524 9722
rect 329472 9658 329524 9664
rect 329484 8974 329512 9658
rect 329472 8968 329524 8974
rect 329472 8910 329524 8916
rect 328368 6452 328420 6458
rect 328368 6394 328420 6400
rect 329668 6390 329696 217534
rect 329656 6384 329708 6390
rect 329656 6326 329708 6332
rect 329760 6322 329788 220116
rect 330220 217598 330248 220116
rect 330484 218068 330536 218074
rect 330484 218010 330536 218016
rect 330208 217592 330260 217598
rect 330208 217534 330260 217540
rect 329748 6316 329800 6322
rect 329748 6258 329800 6264
rect 330024 4412 330076 4418
rect 330024 4354 330076 4360
rect 328828 4004 328880 4010
rect 328828 3946 328880 3952
rect 327724 3324 327776 3330
rect 327724 3266 327776 3272
rect 328840 400 328868 3946
rect 330036 400 330064 4354
rect 330496 4010 330524 218010
rect 330588 216782 330616 220116
rect 331062 220102 331168 220130
rect 331036 217592 331088 217598
rect 331036 217534 331088 217540
rect 330576 216776 330628 216782
rect 330576 216718 330628 216724
rect 331048 8945 331076 217534
rect 331034 8936 331090 8945
rect 331034 8871 331090 8880
rect 331140 6254 331168 220102
rect 331310 217832 331366 217841
rect 331310 217767 331366 217776
rect 331324 217734 331352 217767
rect 331416 217734 331444 220116
rect 331312 217728 331364 217734
rect 331312 217670 331364 217676
rect 331404 217728 331456 217734
rect 331404 217670 331456 217676
rect 331784 217297 331812 220116
rect 332258 220102 332548 220130
rect 332416 217728 332468 217734
rect 332416 217670 332468 217676
rect 331770 217288 331826 217297
rect 331770 217223 331826 217232
rect 332428 12442 332456 217670
rect 332416 12436 332468 12442
rect 332416 12378 332468 12384
rect 331128 6248 331180 6254
rect 331128 6190 331180 6196
rect 332520 6186 332548 220102
rect 332612 217462 332640 220116
rect 333086 220102 333376 220130
rect 332600 217456 332652 217462
rect 332600 217398 332652 217404
rect 333348 214606 333376 220102
rect 333440 217734 333468 220116
rect 333624 220102 333914 220130
rect 334282 220102 334664 220130
rect 333428 217728 333480 217734
rect 333428 217670 333480 217676
rect 333336 214600 333388 214606
rect 333336 214542 333388 214548
rect 333624 12714 333652 220102
rect 334636 218210 334664 220102
rect 334624 218204 334676 218210
rect 334624 218146 334676 218152
rect 334624 218068 334676 218074
rect 334624 218010 334676 218016
rect 333796 217728 333848 217734
rect 333796 217670 333848 217676
rect 333704 217456 333756 217462
rect 333704 217398 333756 217404
rect 333612 12708 333664 12714
rect 333612 12650 333664 12656
rect 333716 12374 333744 217398
rect 333704 12368 333756 12374
rect 333704 12310 333756 12316
rect 333808 6225 333836 217670
rect 333888 214600 333940 214606
rect 333888 214542 333940 214548
rect 333794 6216 333850 6225
rect 332508 6180 332560 6186
rect 333794 6151 333850 6160
rect 332508 6122 332560 6128
rect 331220 4548 331272 4554
rect 331220 4490 331272 4496
rect 330484 4004 330536 4010
rect 330484 3946 330536 3952
rect 331232 400 331260 4490
rect 333612 4480 333664 4486
rect 333612 4422 333664 4428
rect 332414 3360 332470 3369
rect 332414 3295 332470 3304
rect 332428 400 332456 3295
rect 333624 400 333652 4422
rect 333900 3874 333928 214542
rect 333888 3868 333940 3874
rect 333888 3810 333940 3816
rect 334636 2922 334664 218010
rect 334728 217734 334756 220116
rect 335110 220102 335216 220130
rect 334716 217728 334768 217734
rect 334716 217670 334768 217676
rect 335188 12782 335216 220102
rect 335464 217870 335492 220116
rect 335452 217864 335504 217870
rect 335452 217806 335504 217812
rect 335924 217734 335952 220116
rect 336306 220102 336504 220130
rect 335268 217728 335320 217734
rect 335268 217670 335320 217676
rect 335912 217728 335964 217734
rect 335912 217670 335964 217676
rect 335176 12776 335228 12782
rect 335176 12718 335228 12724
rect 335280 12306 335308 217670
rect 335268 12300 335320 12306
rect 335268 12242 335320 12248
rect 336476 12238 336504 220102
rect 336752 217870 336780 220116
rect 336648 217864 336700 217870
rect 336648 217806 336700 217812
rect 336740 217864 336792 217870
rect 336740 217806 336792 217812
rect 336556 217728 336608 217734
rect 336556 217670 336608 217676
rect 336464 12232 336516 12238
rect 336464 12174 336516 12180
rect 336568 10878 336596 217670
rect 336556 10872 336608 10878
rect 336556 10814 336608 10820
rect 334716 4616 334768 4622
rect 334716 4558 334768 4564
rect 334624 2916 334676 2922
rect 334624 2858 334676 2864
rect 334728 400 334756 4558
rect 336660 3806 336688 217806
rect 337120 217462 337148 220116
rect 337580 217734 337608 220116
rect 337856 220102 337962 220130
rect 337752 217864 337804 217870
rect 337752 217806 337804 217812
rect 337568 217728 337620 217734
rect 337568 217670 337620 217676
rect 337108 217456 337160 217462
rect 337108 217398 337160 217404
rect 337384 216776 337436 216782
rect 337384 216718 337436 216724
rect 337108 4684 337160 4690
rect 337108 4626 337160 4632
rect 335912 3800 335964 3806
rect 335912 3742 335964 3748
rect 336648 3800 336700 3806
rect 336648 3742 336700 3748
rect 335924 400 335952 3742
rect 337120 400 337148 4626
rect 337396 3942 337424 216718
rect 337764 12850 337792 217806
rect 337856 12918 337884 220102
rect 338316 217734 338344 220116
rect 337936 217728 337988 217734
rect 337936 217670 337988 217676
rect 338304 217728 338356 217734
rect 338304 217670 338356 217676
rect 337844 12912 337896 12918
rect 337844 12854 337896 12860
rect 337752 12844 337804 12850
rect 337752 12786 337804 12792
rect 337948 12170 337976 217670
rect 338028 217456 338080 217462
rect 338028 217398 338080 217404
rect 337936 12164 337988 12170
rect 337936 12106 337988 12112
rect 338040 10810 338068 217398
rect 338776 217394 338804 220116
rect 339158 220102 339264 220130
rect 338764 217388 338816 217394
rect 338764 217330 338816 217336
rect 338210 40624 338266 40633
rect 338210 40559 338266 40568
rect 338224 40225 338252 40559
rect 338210 40216 338266 40225
rect 338210 40151 338266 40160
rect 339236 12986 339264 220102
rect 339408 217728 339460 217734
rect 339408 217670 339460 217676
rect 339316 217388 339368 217394
rect 339316 217330 339368 217336
rect 339224 12980 339276 12986
rect 339224 12922 339276 12928
rect 339328 12102 339356 217330
rect 339316 12096 339368 12102
rect 339316 12038 339368 12044
rect 338028 10804 338080 10810
rect 338028 10746 338080 10752
rect 339420 10742 339448 217670
rect 339604 216782 339632 220116
rect 339972 217462 340000 220116
rect 340446 220102 340552 220130
rect 340144 218136 340196 218142
rect 340144 218078 340196 218084
rect 339960 217456 340012 217462
rect 339960 217398 340012 217404
rect 339592 216776 339644 216782
rect 339592 216718 339644 216724
rect 339408 10736 339460 10742
rect 339408 10678 339460 10684
rect 338304 4752 338356 4758
rect 338304 4694 338356 4700
rect 337384 3936 337436 3942
rect 337384 3878 337436 3884
rect 338316 400 338344 4694
rect 339500 3732 339552 3738
rect 339500 3674 339552 3680
rect 339512 400 339540 3674
rect 340156 3262 340184 218078
rect 340524 13054 340552 220102
rect 340708 220102 340814 220130
rect 340604 217456 340656 217462
rect 340604 217398 340656 217404
rect 340512 13048 340564 13054
rect 340512 12990 340564 12996
rect 340616 12034 340644 217398
rect 340604 12028 340656 12034
rect 340604 11970 340656 11976
rect 340708 10606 340736 220102
rect 340788 217864 340840 217870
rect 340786 217832 340788 217841
rect 340840 217832 340842 217841
rect 340786 217767 340842 217776
rect 341168 217734 341196 220116
rect 341642 220102 341932 220130
rect 342010 220102 342208 220130
rect 341064 217728 341116 217734
rect 341064 217670 341116 217676
rect 341156 217728 341208 217734
rect 341156 217670 341208 217676
rect 341076 216782 341104 217670
rect 340788 216776 340840 216782
rect 340788 216718 340840 216724
rect 341064 216776 341116 216782
rect 341064 216718 341116 216724
rect 341524 216776 341576 216782
rect 341524 216718 341576 216724
rect 340800 10674 340828 216718
rect 340788 10668 340840 10674
rect 340788 10610 340840 10616
rect 340696 10600 340748 10606
rect 340696 10542 340748 10548
rect 340696 5432 340748 5438
rect 340696 5374 340748 5380
rect 340144 3256 340196 3262
rect 340144 3198 340196 3204
rect 340708 400 340736 5374
rect 341536 3398 341564 216718
rect 341904 215234 341932 220102
rect 342076 217728 342128 217734
rect 342076 217670 342128 217676
rect 341904 215206 342024 215234
rect 341996 211138 342024 215206
rect 341800 211132 341852 211138
rect 341800 211074 341852 211080
rect 341984 211132 342036 211138
rect 341984 211074 342036 211080
rect 341812 201521 341840 211074
rect 341798 201512 341854 201521
rect 341798 201447 341854 201456
rect 341982 201512 342038 201521
rect 341982 201447 342038 201456
rect 341996 196058 342024 201447
rect 341904 196030 342024 196058
rect 341904 195922 341932 196030
rect 341904 195894 342024 195922
rect 341996 167090 342024 195894
rect 341904 167062 342024 167090
rect 341904 166954 341932 167062
rect 341904 166926 342024 166954
rect 341996 162858 342024 166926
rect 341984 162852 342036 162858
rect 341984 162794 342036 162800
rect 341984 153264 342036 153270
rect 341984 153206 342036 153212
rect 341996 142186 342024 153206
rect 341984 142180 342036 142186
rect 341984 142122 342036 142128
rect 341984 140820 342036 140826
rect 341984 140762 342036 140768
rect 341996 139398 342024 140762
rect 341984 139392 342036 139398
rect 341984 139334 342036 139340
rect 341708 129804 341760 129810
rect 341708 129746 341760 129752
rect 341720 122754 341748 129746
rect 341720 122726 341840 122754
rect 341812 113218 341840 122726
rect 341800 113212 341852 113218
rect 341800 113154 341852 113160
rect 341892 113212 341944 113218
rect 341892 113154 341944 113160
rect 341904 113082 341932 113154
rect 341892 113076 341944 113082
rect 341892 113018 341944 113024
rect 341984 103556 342036 103562
rect 341984 103498 342036 103504
rect 341996 84386 342024 103498
rect 341984 84380 342036 84386
rect 341984 84322 342036 84328
rect 341984 84244 342036 84250
rect 341984 84186 342036 84192
rect 341996 74662 342024 84186
rect 341984 74656 342036 74662
rect 341984 74598 342036 74604
rect 341984 73296 342036 73302
rect 341904 73244 341984 73250
rect 341904 73238 342036 73244
rect 341904 73222 342024 73238
rect 341904 64938 341932 73222
rect 341892 64932 341944 64938
rect 341892 64874 341944 64880
rect 341984 64796 342036 64802
rect 341984 64738 342036 64744
rect 341996 63510 342024 64738
rect 341984 63504 342036 63510
rect 341984 63446 342036 63452
rect 341892 63436 341944 63442
rect 341892 63378 341944 63384
rect 341904 62121 341932 63378
rect 341706 62112 341762 62121
rect 341706 62047 341762 62056
rect 341890 62112 341946 62121
rect 341890 62047 341946 62056
rect 341720 53530 341748 62047
rect 341720 53502 341932 53530
rect 341904 45626 341932 53502
rect 341892 45620 341944 45626
rect 341892 45562 341944 45568
rect 341892 45484 341944 45490
rect 341892 45426 341944 45432
rect 341904 18426 341932 45426
rect 341892 18420 341944 18426
rect 341892 18362 341944 18368
rect 342088 11966 342116 217670
rect 342076 11960 342128 11966
rect 342076 11902 342128 11908
rect 342180 10538 342208 220102
rect 342456 217734 342484 220116
rect 342838 220102 343220 220130
rect 343298 220102 343588 220130
rect 342444 217728 342496 217734
rect 342444 217670 342496 217676
rect 343192 215234 343220 220102
rect 343456 217728 343508 217734
rect 343456 217670 343508 217676
rect 343192 215206 343312 215234
rect 343284 211138 343312 215206
rect 343272 211132 343324 211138
rect 343272 211074 343324 211080
rect 343272 205624 343324 205630
rect 343272 205566 343324 205572
rect 343284 201498 343312 205566
rect 343284 201470 343404 201498
rect 343376 193225 343404 201470
rect 343178 193216 343234 193225
rect 343178 193151 343234 193160
rect 343362 193216 343418 193225
rect 343362 193151 343418 193160
rect 343192 191826 343220 193151
rect 342996 191820 343048 191826
rect 342996 191762 343048 191768
rect 343180 191820 343232 191826
rect 343180 191762 343232 191768
rect 343008 182209 343036 191762
rect 342994 182200 343050 182209
rect 342994 182135 343050 182144
rect 343178 182200 343234 182209
rect 343178 182135 343234 182144
rect 343192 172553 343220 182135
rect 343178 172544 343234 172553
rect 343178 172479 343234 172488
rect 343362 172544 343418 172553
rect 343362 172479 343418 172488
rect 343376 169726 343404 172479
rect 343272 169720 343324 169726
rect 343272 169662 343324 169668
rect 343364 169720 343416 169726
rect 343364 169662 343416 169668
rect 343284 160313 343312 169662
rect 343270 160304 343326 160313
rect 343270 160239 343326 160248
rect 343270 160168 343326 160177
rect 343270 160103 343326 160112
rect 343284 158710 343312 160103
rect 343272 158704 343324 158710
rect 343272 158646 343324 158652
rect 343364 140820 343416 140826
rect 343364 140762 343416 140768
rect 343376 132530 343404 140762
rect 343272 132524 343324 132530
rect 343272 132466 343324 132472
rect 343364 132524 343416 132530
rect 343364 132466 343416 132472
rect 343284 131102 343312 132466
rect 343272 131096 343324 131102
rect 343272 131038 343324 131044
rect 343272 121508 343324 121514
rect 343272 121450 343324 121456
rect 343284 118130 343312 121450
rect 343192 118102 343312 118130
rect 343192 103442 343220 118102
rect 343100 103414 343220 103442
rect 343100 93906 343128 103414
rect 343088 93900 343140 93906
rect 343088 93842 343140 93848
rect 343180 93900 343232 93906
rect 343180 93842 343232 93848
rect 343192 86986 343220 93842
rect 343192 86958 343312 86986
rect 343284 84182 343312 86958
rect 343272 84176 343324 84182
rect 343272 84118 343324 84124
rect 343364 74588 343416 74594
rect 343364 74530 343416 74536
rect 343376 65113 343404 74530
rect 343362 65104 343418 65113
rect 343362 65039 343418 65048
rect 343178 64968 343234 64977
rect 343178 64903 343234 64912
rect 343192 63510 343220 64903
rect 343180 63504 343232 63510
rect 343180 63446 343232 63452
rect 343364 63504 343416 63510
rect 343364 63446 343416 63452
rect 343376 37330 343404 63446
rect 343364 37324 343416 37330
rect 343364 37266 343416 37272
rect 343364 28484 343416 28490
rect 343364 28426 343416 28432
rect 343376 27606 343404 28426
rect 343364 27600 343416 27606
rect 343364 27542 343416 27548
rect 343468 11898 343496 217670
rect 343456 11892 343508 11898
rect 343456 11834 343508 11840
rect 342168 10532 342220 10538
rect 342168 10474 342220 10480
rect 343560 10470 343588 220102
rect 343652 216782 343680 220116
rect 344126 220102 344324 220130
rect 344494 220102 344784 220130
rect 344862 220102 344968 220130
rect 344296 217682 344324 220102
rect 344756 217682 344784 220102
rect 344296 217654 344508 217682
rect 344756 217654 344876 217682
rect 343640 216776 343692 216782
rect 343640 216718 343692 216724
rect 344480 215234 344508 217654
rect 344744 216776 344796 216782
rect 344744 216718 344796 216724
rect 344480 215206 344600 215234
rect 344572 211138 344600 215206
rect 344560 211132 344612 211138
rect 344560 211074 344612 211080
rect 344560 205624 344612 205630
rect 344560 205566 344612 205572
rect 344572 201498 344600 205566
rect 344572 201470 344692 201498
rect 344664 193225 344692 201470
rect 344374 193216 344430 193225
rect 344374 193151 344430 193160
rect 344650 193216 344706 193225
rect 344650 193151 344706 193160
rect 344388 183666 344416 193151
rect 344376 183660 344428 183666
rect 344376 183602 344428 183608
rect 344560 183660 344612 183666
rect 344560 183602 344612 183608
rect 344572 176662 344600 183602
rect 344560 176656 344612 176662
rect 344560 176598 344612 176604
rect 344468 176588 344520 176594
rect 344468 176530 344520 176536
rect 344480 172553 344508 176530
rect 344466 172544 344522 172553
rect 344466 172479 344522 172488
rect 344650 172544 344706 172553
rect 344650 172479 344706 172488
rect 344664 167550 344692 172479
rect 344652 167544 344704 167550
rect 344652 167486 344704 167492
rect 344560 162920 344612 162926
rect 344560 162862 344612 162868
rect 344572 151842 344600 162862
rect 344468 151836 344520 151842
rect 344468 151778 344520 151784
rect 344560 151836 344612 151842
rect 344560 151778 344612 151784
rect 344480 142202 344508 151778
rect 344388 142174 344508 142202
rect 344388 140826 344416 142174
rect 344284 140820 344336 140826
rect 344284 140762 344336 140768
rect 344376 140820 344428 140826
rect 344376 140762 344428 140768
rect 344296 132394 344324 140762
rect 344284 132388 344336 132394
rect 344284 132330 344336 132336
rect 344560 132388 344612 132394
rect 344560 132330 344612 132336
rect 344572 122806 344600 132330
rect 344468 122800 344520 122806
rect 344468 122742 344520 122748
rect 344560 122800 344612 122806
rect 344560 122742 344612 122748
rect 344480 109698 344508 122742
rect 344480 109670 344600 109698
rect 344572 103494 344600 109670
rect 344560 103488 344612 103494
rect 344560 103430 344612 103436
rect 344468 93900 344520 93906
rect 344468 93842 344520 93848
rect 344480 86986 344508 93842
rect 344480 86958 344600 86986
rect 344572 79354 344600 86958
rect 344560 79348 344612 79354
rect 344560 79290 344612 79296
rect 344560 67652 344612 67658
rect 344560 67594 344612 67600
rect 344572 64870 344600 67594
rect 344560 64864 344612 64870
rect 344560 64806 344612 64812
rect 344468 55276 344520 55282
rect 344468 55218 344520 55224
rect 344480 51814 344508 55218
rect 344468 51808 344520 51814
rect 344468 51750 344520 51756
rect 344560 41132 344612 41138
rect 344560 41074 344612 41080
rect 344572 38706 344600 41074
rect 344572 38678 344692 38706
rect 344664 38622 344692 38678
rect 344652 38616 344704 38622
rect 344652 38558 344704 38564
rect 344652 29028 344704 29034
rect 344652 28970 344704 28976
rect 344664 27606 344692 28970
rect 344652 27600 344704 27606
rect 344652 27542 344704 27548
rect 344756 11830 344784 216718
rect 344744 11824 344796 11830
rect 344744 11766 344796 11772
rect 343548 10464 343600 10470
rect 343548 10406 343600 10412
rect 344848 10402 344876 217654
rect 344836 10396 344888 10402
rect 344836 10338 344888 10344
rect 344940 7002 344968 220102
rect 345308 217734 345336 220116
rect 345676 217870 345704 220116
rect 346150 220102 346256 220130
rect 345572 217864 345624 217870
rect 345572 217806 345624 217812
rect 345664 217864 345716 217870
rect 345664 217806 345716 217812
rect 345296 217728 345348 217734
rect 345296 217670 345348 217676
rect 345584 217682 345612 217806
rect 346124 217728 346176 217734
rect 345584 217654 345796 217682
rect 346124 217670 346176 217676
rect 345664 216708 345716 216714
rect 345664 216650 345716 216656
rect 345676 196058 345704 216650
rect 345584 196030 345704 196058
rect 345584 195922 345612 196030
rect 345584 195894 345704 195922
rect 345676 172514 345704 195894
rect 345480 172508 345532 172514
rect 345480 172450 345532 172456
rect 345664 172508 345716 172514
rect 345664 172450 345716 172456
rect 345492 162897 345520 172450
rect 345478 162888 345534 162897
rect 345478 162823 345534 162832
rect 345662 162888 345718 162897
rect 345662 162823 345718 162832
rect 345676 161430 345704 162823
rect 345664 161424 345716 161430
rect 345664 161366 345716 161372
rect 345664 151836 345716 151842
rect 345664 151778 345716 151784
rect 345676 148322 345704 151778
rect 345584 148294 345704 148322
rect 345584 138106 345612 148294
rect 345572 138100 345624 138106
rect 345572 138042 345624 138048
rect 345662 132560 345718 132569
rect 345584 132518 345662 132546
rect 345584 132462 345612 132518
rect 345662 132495 345718 132504
rect 345572 132456 345624 132462
rect 345572 132398 345624 132404
rect 345572 122868 345624 122874
rect 345572 122810 345624 122816
rect 345584 122754 345612 122810
rect 345492 122726 345612 122754
rect 345492 114458 345520 122726
rect 345492 114430 345612 114458
rect 345584 104802 345612 114430
rect 345584 104774 345704 104802
rect 345676 86986 345704 104774
rect 345584 86958 345704 86986
rect 345584 84182 345612 86958
rect 345572 84176 345624 84182
rect 345572 84118 345624 84124
rect 345664 74588 345716 74594
rect 345664 74530 345716 74536
rect 345676 64818 345704 74530
rect 345584 64790 345704 64818
rect 345584 60042 345612 64790
rect 345572 60036 345624 60042
rect 345572 59978 345624 59984
rect 345664 46980 345716 46986
rect 345664 46922 345716 46928
rect 345676 27606 345704 46922
rect 345664 27600 345716 27606
rect 345664 27542 345716 27548
rect 345664 18012 345716 18018
rect 345664 17954 345716 17960
rect 344928 6996 344980 7002
rect 344928 6938 344980 6944
rect 341892 5500 341944 5506
rect 341892 5442 341944 5448
rect 341524 3392 341576 3398
rect 341524 3334 341576 3340
rect 341904 400 341932 5442
rect 345480 5364 345532 5370
rect 345480 5306 345532 5312
rect 344284 5296 344336 5302
rect 344284 5238 344336 5244
rect 343088 3664 343140 3670
rect 343088 3606 343140 3612
rect 343100 400 343128 3606
rect 344296 400 344324 5238
rect 345492 400 345520 5306
rect 345676 4078 345704 17954
rect 345664 4072 345716 4078
rect 345664 4014 345716 4020
rect 345768 2854 345796 217654
rect 345848 138100 345900 138106
rect 345848 138042 345900 138048
rect 345860 132569 345888 138042
rect 345846 132560 345902 132569
rect 345846 132495 345902 132504
rect 346136 13598 346164 217670
rect 346124 13592 346176 13598
rect 346124 13534 346176 13540
rect 346228 7070 346256 220102
rect 346504 217870 346532 220116
rect 346308 217864 346360 217870
rect 346308 217806 346360 217812
rect 346492 217864 346544 217870
rect 346492 217806 346544 217812
rect 346216 7064 346268 7070
rect 346216 7006 346268 7012
rect 346320 4214 346348 217806
rect 346964 210458 346992 220116
rect 347346 220102 347636 220130
rect 347504 217864 347556 217870
rect 347504 217806 347556 217812
rect 347412 217728 347464 217734
rect 347412 217670 347464 217676
rect 346952 210452 347004 210458
rect 346952 210394 347004 210400
rect 347424 13530 347452 217670
rect 347412 13524 347464 13530
rect 347412 13466 347464 13472
rect 347516 10334 347544 217806
rect 347504 10328 347556 10334
rect 347504 10270 347556 10276
rect 346676 8084 346728 8090
rect 346676 8026 346728 8032
rect 346308 4208 346360 4214
rect 346308 4150 346360 4156
rect 345756 2848 345808 2854
rect 345756 2790 345808 2796
rect 346688 400 346716 8026
rect 347608 7138 347636 220102
rect 347700 217734 347728 220116
rect 348160 217870 348188 220116
rect 348148 217864 348200 217870
rect 348148 217806 348200 217812
rect 348528 217734 348556 220116
rect 348896 220102 349002 220130
rect 347688 217728 347740 217734
rect 347688 217670 347740 217676
rect 348516 217728 348568 217734
rect 348516 217670 348568 217676
rect 347688 210452 347740 210458
rect 347688 210394 347740 210400
rect 347596 7132 347648 7138
rect 347596 7074 347648 7080
rect 347700 4282 347728 210394
rect 348896 13462 348924 220102
rect 349356 218006 349384 220116
rect 349344 218000 349396 218006
rect 349344 217942 349396 217948
rect 349068 217864 349120 217870
rect 349068 217806 349120 217812
rect 348976 217728 349028 217734
rect 348976 217670 349028 217676
rect 348884 13456 348936 13462
rect 348884 13398 348936 13404
rect 348988 9874 349016 217670
rect 348804 9846 349016 9874
rect 348804 7206 348832 9846
rect 349080 8242 349108 217806
rect 349816 217734 349844 220116
rect 350198 220102 350304 220130
rect 349804 217728 349856 217734
rect 349804 217670 349856 217676
rect 350276 13394 350304 220102
rect 350448 218000 350500 218006
rect 350448 217942 350500 217948
rect 350356 217728 350408 217734
rect 350356 217670 350408 217676
rect 350264 13388 350316 13394
rect 350264 13330 350316 13336
rect 348988 8214 349108 8242
rect 348792 7200 348844 7206
rect 348792 7142 348844 7148
rect 347872 5228 347924 5234
rect 347872 5170 347924 5176
rect 347688 4276 347740 4282
rect 347688 4218 347740 4224
rect 347884 400 347912 5170
rect 348988 4350 349016 8214
rect 349068 8016 349120 8022
rect 349068 7958 349120 7964
rect 348976 4344 349028 4350
rect 348976 4286 349028 4292
rect 349080 400 349108 7958
rect 350368 7274 350396 217670
rect 350356 7268 350408 7274
rect 350356 7210 350408 7216
rect 350460 4418 350488 217942
rect 350644 217802 350672 220116
rect 350632 217796 350684 217802
rect 350632 217738 350684 217744
rect 351012 217734 351040 220116
rect 351394 220102 351592 220130
rect 351000 217728 351052 217734
rect 351000 217670 351052 217676
rect 351564 13326 351592 220102
rect 351748 220102 351854 220130
rect 351644 217728 351696 217734
rect 351644 217670 351696 217676
rect 351552 13320 351604 13326
rect 351552 13262 351604 13268
rect 351656 7342 351684 217670
rect 351644 7336 351696 7342
rect 351644 7278 351696 7284
rect 351368 5160 351420 5166
rect 351368 5102 351420 5108
rect 350448 4412 350500 4418
rect 350448 4354 350500 4360
rect 350264 3596 350316 3602
rect 350264 3538 350316 3544
rect 350276 400 350304 3538
rect 351380 400 351408 5102
rect 351748 4554 351776 220102
rect 351828 217796 351880 217802
rect 351828 217738 351880 217744
rect 351736 4548 351788 4554
rect 351736 4490 351788 4496
rect 351840 4486 351868 217738
rect 352208 217734 352236 220116
rect 352682 220102 352972 220130
rect 353050 220102 353248 220130
rect 352564 217864 352616 217870
rect 352564 217806 352616 217812
rect 352196 217728 352248 217734
rect 352196 217670 352248 217676
rect 352576 8242 352604 217806
rect 352944 215234 352972 220102
rect 353116 217728 353168 217734
rect 353116 217670 353168 217676
rect 352944 215206 353064 215234
rect 353036 212537 353064 215206
rect 352838 212528 352894 212537
rect 352838 212463 352894 212472
rect 353022 212528 353078 212537
rect 353022 212463 353078 212472
rect 352852 202910 352880 212463
rect 352840 202904 352892 202910
rect 352840 202846 352892 202852
rect 353024 202904 353076 202910
rect 353024 202846 353076 202852
rect 353036 196058 353064 202846
rect 352944 196030 353064 196058
rect 352944 195922 352972 196030
rect 352944 195894 353064 195922
rect 353036 167090 353064 195894
rect 352944 167062 353064 167090
rect 352944 166954 352972 167062
rect 352944 166926 353064 166954
rect 353036 147778 353064 166926
rect 352944 147750 353064 147778
rect 352944 147642 352972 147750
rect 352944 147614 353064 147642
rect 353036 128466 353064 147614
rect 352944 128438 353064 128466
rect 352944 128330 352972 128438
rect 352944 128302 353064 128330
rect 353036 109154 353064 128302
rect 352944 109126 353064 109154
rect 352944 109018 352972 109126
rect 352944 108990 353064 109018
rect 353036 89842 353064 108990
rect 352944 89814 353064 89842
rect 352944 89706 352972 89814
rect 352944 89678 353064 89706
rect 353036 70394 353064 89678
rect 352944 70366 353064 70394
rect 352944 70258 352972 70366
rect 352944 70230 353064 70258
rect 353036 51082 353064 70230
rect 352944 51054 353064 51082
rect 352944 50946 352972 51054
rect 352944 50918 353064 50946
rect 353036 31770 353064 50918
rect 352944 31742 353064 31770
rect 352944 19310 352972 31742
rect 352932 19304 352984 19310
rect 352932 19246 352984 19252
rect 352484 8214 352604 8242
rect 351828 4480 351880 4486
rect 351828 4422 351880 4428
rect 352484 4146 352512 8214
rect 352564 7948 352616 7954
rect 352564 7890 352616 7896
rect 352472 4140 352524 4146
rect 352472 4082 352524 4088
rect 352576 400 352604 7890
rect 353128 7410 353156 217670
rect 353116 7404 353168 7410
rect 353116 7346 353168 7352
rect 353220 4622 353248 220102
rect 353496 217734 353524 220116
rect 353878 220102 354076 220130
rect 354246 220102 354628 220130
rect 353484 217728 353536 217734
rect 354048 217716 354076 220102
rect 354496 217728 354548 217734
rect 354048 217688 354260 217716
rect 353484 217670 353536 217676
rect 354232 215234 354260 217688
rect 354496 217670 354548 217676
rect 354232 215206 354352 215234
rect 354324 212514 354352 215206
rect 354232 212486 354352 212514
rect 354232 211138 354260 212486
rect 354128 211132 354180 211138
rect 354128 211074 354180 211080
rect 354220 211132 354272 211138
rect 354220 211074 354272 211080
rect 354140 201521 354168 211074
rect 354126 201512 354182 201521
rect 354126 201447 354182 201456
rect 354402 201512 354458 201521
rect 354402 201447 354458 201456
rect 354416 193225 354444 201447
rect 354218 193216 354274 193225
rect 354218 193151 354274 193160
rect 354402 193216 354458 193225
rect 354402 193151 354458 193160
rect 354232 191826 354260 193151
rect 354220 191820 354272 191826
rect 354220 191762 354272 191768
rect 354220 183524 354272 183530
rect 354220 183466 354272 183472
rect 354232 182186 354260 183466
rect 354232 182170 354352 182186
rect 354232 182164 354364 182170
rect 354232 182158 354312 182164
rect 354312 182106 354364 182112
rect 354404 176588 354456 176594
rect 354404 176530 354456 176536
rect 354416 164286 354444 176530
rect 354312 164280 354364 164286
rect 354312 164222 354364 164228
rect 354404 164280 354456 164286
rect 354404 164222 354456 164228
rect 354324 162858 354352 164222
rect 354312 162852 354364 162858
rect 354312 162794 354364 162800
rect 354312 157344 354364 157350
rect 354312 157286 354364 157292
rect 354324 153218 354352 157286
rect 354324 153190 354444 153218
rect 354416 147830 354444 153190
rect 354404 147824 354456 147830
rect 354404 147766 354456 147772
rect 354404 147688 354456 147694
rect 354404 147630 354456 147636
rect 354416 128382 354444 147630
rect 354404 128376 354456 128382
rect 354404 128318 354456 128324
rect 354404 124228 354456 124234
rect 354404 124170 354456 124176
rect 354416 114646 354444 124170
rect 354404 114640 354456 114646
rect 354404 114582 354456 114588
rect 354220 113212 354272 113218
rect 354220 113154 354272 113160
rect 354232 109750 354260 113154
rect 354220 109744 354272 109750
rect 354220 109686 354272 109692
rect 354404 96688 354456 96694
rect 354404 96630 354456 96636
rect 354416 58206 354444 96630
rect 354404 58200 354456 58206
rect 354404 58142 354456 58148
rect 354404 58064 354456 58070
rect 354404 58006 354456 58012
rect 354416 57934 354444 58006
rect 354404 57928 354456 57934
rect 354404 57870 354456 57876
rect 354312 48408 354364 48414
rect 354312 48350 354364 48356
rect 354324 48278 354352 48350
rect 354312 48272 354364 48278
rect 354312 48214 354364 48220
rect 354312 41132 354364 41138
rect 354312 41074 354364 41080
rect 354324 38706 354352 41074
rect 354324 38678 354444 38706
rect 354416 27606 354444 38678
rect 354404 27600 354456 27606
rect 354404 27542 354456 27548
rect 354312 18012 354364 18018
rect 354312 17954 354364 17960
rect 354324 13258 354352 17954
rect 354312 13252 354364 13258
rect 354312 13194 354364 13200
rect 354508 7478 354536 217670
rect 354496 7472 354548 7478
rect 354496 7414 354548 7420
rect 354600 4690 354628 220102
rect 354692 217802 354720 220116
rect 355060 217870 355088 220116
rect 355048 217864 355100 217870
rect 355048 217806 355100 217812
rect 354680 217796 354732 217802
rect 354680 217738 354732 217744
rect 355520 217734 355548 220116
rect 355796 220102 355902 220130
rect 355600 217864 355652 217870
rect 355600 217806 355652 217812
rect 355508 217728 355560 217734
rect 355508 217670 355560 217676
rect 355612 211138 355640 217806
rect 355416 211132 355468 211138
rect 355416 211074 355468 211080
rect 355600 211132 355652 211138
rect 355600 211074 355652 211080
rect 355428 201521 355456 211074
rect 355414 201512 355470 201521
rect 355414 201447 355470 201456
rect 355690 201512 355746 201521
rect 355690 201447 355746 201456
rect 355704 193225 355732 201447
rect 355414 193216 355470 193225
rect 355414 193151 355470 193160
rect 355690 193216 355746 193225
rect 355690 193151 355746 193160
rect 355428 191826 355456 193151
rect 355416 191820 355468 191826
rect 355416 191762 355468 191768
rect 355508 191820 355560 191826
rect 355508 191762 355560 191768
rect 355520 182186 355548 191762
rect 355520 182170 355640 182186
rect 355520 182164 355652 182170
rect 355520 182158 355600 182164
rect 355600 182106 355652 182112
rect 355600 176656 355652 176662
rect 355600 176598 355652 176604
rect 355612 172530 355640 176598
rect 355612 172502 355732 172530
rect 355704 167074 355732 172502
rect 355692 167068 355744 167074
rect 355692 167010 355744 167016
rect 355600 164280 355652 164286
rect 355600 164222 355652 164228
rect 355612 162858 355640 164222
rect 355600 162852 355652 162858
rect 355600 162794 355652 162800
rect 355508 153264 355560 153270
rect 355508 153206 355560 153212
rect 355520 144945 355548 153206
rect 355506 144936 355562 144945
rect 355506 144871 355562 144880
rect 355690 144936 355746 144945
rect 355690 144871 355746 144880
rect 355704 128382 355732 144871
rect 355692 128376 355744 128382
rect 355692 128318 355744 128324
rect 355796 125594 355824 220102
rect 355876 217796 355928 217802
rect 355876 217738 355928 217744
rect 355784 125588 355836 125594
rect 355784 125530 355836 125536
rect 355784 125452 355836 125458
rect 355784 125394 355836 125400
rect 355692 124228 355744 124234
rect 355692 124170 355744 124176
rect 355704 114458 355732 124170
rect 355612 114430 355732 114458
rect 355612 113150 355640 114430
rect 355600 113144 355652 113150
rect 355600 113086 355652 113092
rect 355692 103556 355744 103562
rect 355692 103498 355744 103504
rect 355704 93838 355732 103498
rect 355692 93832 355744 93838
rect 355692 93774 355744 93780
rect 355692 84244 355744 84250
rect 355692 84186 355744 84192
rect 355704 79506 355732 84186
rect 355612 79478 355732 79506
rect 355612 71074 355640 79478
rect 355796 75750 355824 125394
rect 355888 75818 355916 217738
rect 356348 217734 356376 220116
rect 356716 217802 356744 220116
rect 357190 220102 357296 220130
rect 356704 217796 356756 217802
rect 356704 217738 356756 217744
rect 355968 217728 356020 217734
rect 355968 217670 356020 217676
rect 356336 217728 356388 217734
rect 356336 217670 356388 217676
rect 357164 217728 357216 217734
rect 357164 217670 357216 217676
rect 355980 75886 356008 217670
rect 355968 75880 356020 75886
rect 355968 75822 356020 75828
rect 355876 75812 355928 75818
rect 355876 75754 355928 75760
rect 355784 75744 355836 75750
rect 355784 75686 355836 75692
rect 355876 75676 355928 75682
rect 355876 75618 355928 75624
rect 355784 75608 355836 75614
rect 355784 75550 355836 75556
rect 355612 71046 355732 71074
rect 355704 64870 355732 71046
rect 355692 64864 355744 64870
rect 355692 64806 355744 64812
rect 355600 48340 355652 48346
rect 355600 48282 355652 48288
rect 355612 38706 355640 48282
rect 355612 38678 355732 38706
rect 355704 27606 355732 38678
rect 355692 27600 355744 27606
rect 355692 27542 355744 27548
rect 355508 18012 355560 18018
rect 355508 17954 355560 17960
rect 355520 13190 355548 17954
rect 355508 13184 355560 13190
rect 355508 13126 355560 13132
rect 355796 8294 355824 75550
rect 355784 8288 355836 8294
rect 355784 8230 355836 8236
rect 355888 7546 355916 75618
rect 355968 67380 356020 67386
rect 355968 67322 356020 67328
rect 355876 7540 355928 7546
rect 355876 7482 355928 7488
rect 354956 5092 355008 5098
rect 354956 5034 355008 5040
rect 354588 4684 354640 4690
rect 354588 4626 354640 4632
rect 353208 4616 353260 4622
rect 353208 4558 353260 4564
rect 353760 3528 353812 3534
rect 353760 3470 353812 3476
rect 353772 400 353800 3470
rect 354968 400 354996 5034
rect 355980 4758 356008 67322
rect 357176 13122 357204 217670
rect 357164 13116 357216 13122
rect 357164 13058 357216 13064
rect 357268 8226 357296 220102
rect 357348 217796 357400 217802
rect 357348 217738 357400 217744
rect 357256 8220 357308 8226
rect 357256 8162 357308 8168
rect 356152 7880 356204 7886
rect 356152 7822 356204 7828
rect 355968 4752 356020 4758
rect 355968 4694 356020 4700
rect 356164 400 356192 7822
rect 357360 5506 357388 217738
rect 357544 217734 357572 220116
rect 357912 217802 357940 220116
rect 358386 220102 358676 220130
rect 358084 217932 358136 217938
rect 358084 217874 358136 217880
rect 357900 217796 357952 217802
rect 357900 217738 357952 217744
rect 357532 217728 357584 217734
rect 357532 217670 357584 217676
rect 357348 5500 357400 5506
rect 357348 5442 357400 5448
rect 358096 3466 358124 217874
rect 358544 217728 358596 217734
rect 358544 217670 358596 217676
rect 358556 14482 358584 217670
rect 358544 14476 358596 14482
rect 358544 14418 358596 14424
rect 358648 8158 358676 220102
rect 358740 218006 358768 220116
rect 358728 218000 358780 218006
rect 358728 217942 358780 217948
rect 358728 217796 358780 217802
rect 358728 217738 358780 217744
rect 358636 8152 358688 8158
rect 358636 8094 358688 8100
rect 358740 5438 358768 217738
rect 359200 217734 359228 220116
rect 359582 220102 359964 220130
rect 360042 220102 360148 220130
rect 359188 217728 359240 217734
rect 359188 217670 359240 217676
rect 359936 8090 359964 220102
rect 360016 217728 360068 217734
rect 360016 217670 360068 217676
rect 359924 8084 359976 8090
rect 359924 8026 359976 8032
rect 359740 7812 359792 7818
rect 359740 7754 359792 7760
rect 358728 5432 358780 5438
rect 358728 5374 358780 5380
rect 358544 5024 358596 5030
rect 358544 4966 358596 4972
rect 357348 3460 357400 3466
rect 357348 3402 357400 3408
rect 358084 3460 358136 3466
rect 358084 3402 358136 3408
rect 357360 400 357388 3402
rect 358556 400 358584 4966
rect 359752 400 359780 7754
rect 360028 5370 360056 217670
rect 360016 5364 360068 5370
rect 360016 5306 360068 5312
rect 360120 3738 360148 220102
rect 360396 217734 360424 220116
rect 360384 217728 360436 217734
rect 360384 217670 360436 217676
rect 360764 212566 360792 220116
rect 361224 216782 361252 220116
rect 361592 217802 361620 220116
rect 362052 217870 362080 220116
rect 362040 217864 362092 217870
rect 362040 217806 362092 217812
rect 361580 217796 361632 217802
rect 361580 217738 361632 217744
rect 362420 217734 362448 220116
rect 362696 220102 362894 220130
rect 362592 217864 362644 217870
rect 362592 217806 362644 217812
rect 361488 217728 361540 217734
rect 361488 217670 361540 217676
rect 362408 217728 362460 217734
rect 362408 217670 362460 217676
rect 361212 216776 361264 216782
rect 361212 216718 361264 216724
rect 360752 212560 360804 212566
rect 360752 212502 360804 212508
rect 361304 212560 361356 212566
rect 361304 212502 361356 212508
rect 361316 196058 361344 212502
rect 361224 196030 361344 196058
rect 361224 186130 361252 196030
rect 361224 186102 361344 186130
rect 361316 183546 361344 186102
rect 361224 183518 361344 183546
rect 361224 182170 361252 183518
rect 360936 182164 360988 182170
rect 360936 182106 360988 182112
rect 361212 182164 361264 182170
rect 361212 182106 361264 182112
rect 360948 172553 360976 182106
rect 360934 172544 360990 172553
rect 360934 172479 360990 172488
rect 361118 172544 361174 172553
rect 361118 172479 361120 172488
rect 361172 172479 361174 172488
rect 361396 172508 361448 172514
rect 361120 172450 361172 172456
rect 361396 172450 361448 172456
rect 361408 161514 361436 172450
rect 361224 161486 361436 161514
rect 361224 160070 361252 161486
rect 361212 160064 361264 160070
rect 361212 160006 361264 160012
rect 361304 150476 361356 150482
rect 361304 150418 361356 150424
rect 361316 143426 361344 150418
rect 361316 143398 361436 143426
rect 361408 142118 361436 143398
rect 361396 142112 361448 142118
rect 361396 142054 361448 142060
rect 361396 132524 361448 132530
rect 361396 132466 361448 132472
rect 361408 124234 361436 132466
rect 361304 124228 361356 124234
rect 361304 124170 361356 124176
rect 361396 124228 361448 124234
rect 361396 124170 361448 124176
rect 361316 116006 361344 124170
rect 361212 116000 361264 116006
rect 361212 115942 361264 115948
rect 361304 116000 361356 116006
rect 361304 115942 361356 115948
rect 361224 106457 361252 115942
rect 361210 106448 361266 106457
rect 361210 106383 361266 106392
rect 361302 106312 361358 106321
rect 361302 106247 361358 106256
rect 361316 99906 361344 106247
rect 361224 99878 361344 99906
rect 361224 93838 361252 99878
rect 361212 93832 361264 93838
rect 361212 93774 361264 93780
rect 361212 85536 361264 85542
rect 361212 85478 361264 85484
rect 361224 84266 361252 85478
rect 361224 84238 361344 84266
rect 361316 84182 361344 84238
rect 361304 84176 361356 84182
rect 361304 84118 361356 84124
rect 361396 79348 361448 79354
rect 361396 79290 361448 79296
rect 361408 70258 361436 79290
rect 361316 70230 361436 70258
rect 361316 58018 361344 70230
rect 361224 57990 361344 58018
rect 361224 53122 361252 57990
rect 361224 53094 361436 53122
rect 361408 50946 361436 53094
rect 361316 50918 361436 50946
rect 361316 41426 361344 50918
rect 361316 41398 361436 41426
rect 361408 31822 361436 41398
rect 361396 31816 361448 31822
rect 361396 31758 361448 31764
rect 361304 29028 361356 29034
rect 361304 28970 361356 28976
rect 361316 27606 361344 28970
rect 361304 27600 361356 27606
rect 361304 27542 361356 27548
rect 361212 18012 361264 18018
rect 361212 17954 361264 17960
rect 361224 12322 361252 17954
rect 361224 12294 361344 12322
rect 361316 8022 361344 12294
rect 361304 8016 361356 8022
rect 361304 7958 361356 7964
rect 361500 5302 361528 217670
rect 362604 201482 362632 217806
rect 362592 201476 362644 201482
rect 362592 201418 362644 201424
rect 362500 191888 362552 191894
rect 362500 191830 362552 191836
rect 362512 183546 362540 191830
rect 362512 183518 362632 183546
rect 362604 182170 362632 183518
rect 362592 182164 362644 182170
rect 362592 182106 362644 182112
rect 362316 171216 362368 171222
rect 362368 171164 362448 171170
rect 362316 171158 362448 171164
rect 362328 171142 362448 171158
rect 362420 171086 362448 171142
rect 362408 171080 362460 171086
rect 362408 171022 362460 171028
rect 362408 161492 362460 161498
rect 362408 161434 362460 161440
rect 362420 156670 362448 161434
rect 362408 156664 362460 156670
rect 362408 156606 362460 156612
rect 362408 144900 362460 144906
rect 362408 144842 362460 144848
rect 362420 143562 362448 144842
rect 362420 143534 362540 143562
rect 362512 137850 362540 143534
rect 362328 137822 362540 137850
rect 362328 127702 362356 137822
rect 362316 127696 362368 127702
rect 362316 127638 362368 127644
rect 362592 127696 362644 127702
rect 362592 127638 362644 127644
rect 362604 122913 362632 127638
rect 362314 122904 362370 122913
rect 362314 122839 362370 122848
rect 362590 122904 362646 122913
rect 362590 122839 362646 122848
rect 362328 121446 362356 122839
rect 362316 121440 362368 121446
rect 362316 121382 362368 121388
rect 362316 115932 362368 115938
rect 362316 115874 362368 115880
rect 362328 85610 362356 115874
rect 362316 85604 362368 85610
rect 362316 85546 362368 85552
rect 362500 85604 362552 85610
rect 362500 85546 362552 85552
rect 362512 84182 362540 85546
rect 362500 84176 362552 84182
rect 362500 84118 362552 84124
rect 362316 67652 362368 67658
rect 362316 67594 362368 67600
rect 362328 67522 362356 67594
rect 362224 67516 362276 67522
rect 362224 67458 362276 67464
rect 362316 67516 362368 67522
rect 362316 67458 362368 67464
rect 362236 67130 362264 67458
rect 362236 67102 362356 67130
rect 362328 57934 362356 67102
rect 362316 57928 362368 57934
rect 362316 57870 362368 57876
rect 362500 48340 362552 48346
rect 362500 48282 362552 48288
rect 362512 41426 362540 48282
rect 362512 41398 362632 41426
rect 362604 31890 362632 41398
rect 362592 31884 362644 31890
rect 362592 31826 362644 31832
rect 362408 29028 362460 29034
rect 362408 28970 362460 28976
rect 362420 22114 362448 28970
rect 362420 22086 362632 22114
rect 362604 19310 362632 22086
rect 362592 19304 362644 19310
rect 362592 19246 362644 19252
rect 362500 9716 362552 9722
rect 362500 9658 362552 9664
rect 362512 9625 362540 9658
rect 362498 9616 362554 9625
rect 362498 9551 362554 9560
rect 361488 5296 361540 5302
rect 361488 5238 361540 5244
rect 362696 5166 362724 220102
rect 362776 217796 362828 217802
rect 362776 217738 362828 217744
rect 362788 5234 362816 217738
rect 363248 217734 363276 220116
rect 363708 217870 363736 220116
rect 364090 220102 364288 220130
rect 363696 217864 363748 217870
rect 363696 217806 363748 217812
rect 362868 217728 362920 217734
rect 362868 217670 362920 217676
rect 363236 217728 363288 217734
rect 363236 217670 363288 217676
rect 364156 217728 364208 217734
rect 364156 217670 364208 217676
rect 362776 5228 362828 5234
rect 362776 5170 362828 5176
rect 362684 5160 362736 5166
rect 362684 5102 362736 5108
rect 362132 4956 362184 4962
rect 362132 4898 362184 4904
rect 360108 3732 360160 3738
rect 360108 3674 360160 3680
rect 360936 3052 360988 3058
rect 360936 2994 360988 3000
rect 360948 400 360976 2994
rect 362144 400 362172 4898
rect 362880 3670 362908 217670
rect 363602 9480 363658 9489
rect 363602 9415 363658 9424
rect 363616 7954 363644 9415
rect 363604 7948 363656 7954
rect 363604 7890 363656 7896
rect 364168 7886 364196 217670
rect 364156 7880 364208 7886
rect 364156 7822 364208 7828
rect 363328 7744 363380 7750
rect 363328 7686 363380 7692
rect 362868 3664 362920 3670
rect 362868 3606 362920 3612
rect 363340 400 363368 7686
rect 364260 5098 364288 220102
rect 364444 217734 364472 220116
rect 364904 217802 364932 220116
rect 365286 220102 365576 220130
rect 364892 217796 364944 217802
rect 364892 217738 364944 217744
rect 364432 217728 364484 217734
rect 364432 217670 364484 217676
rect 365444 217728 365496 217734
rect 365444 217670 365496 217676
rect 365456 7818 365484 217670
rect 365444 7812 365496 7818
rect 365444 7754 365496 7760
rect 364524 7608 364576 7614
rect 364524 7550 364576 7556
rect 364248 5092 364300 5098
rect 364248 5034 364300 5040
rect 364536 400 364564 7550
rect 365548 5030 365576 220102
rect 365732 217802 365760 220116
rect 366100 217938 366128 220116
rect 366088 217932 366140 217938
rect 366088 217874 366140 217880
rect 365628 217796 365680 217802
rect 365628 217738 365680 217744
rect 365720 217796 365772 217802
rect 365720 217738 365772 217744
rect 365536 5024 365588 5030
rect 365536 4966 365588 4972
rect 365640 3602 365668 217738
rect 366560 217734 366588 220116
rect 366824 217796 366876 217802
rect 366824 217738 366876 217744
rect 366548 217728 366600 217734
rect 366548 217670 366600 217676
rect 366732 11076 366784 11082
rect 366732 11018 366784 11024
rect 366744 4962 366772 11018
rect 366836 7750 366864 217738
rect 366928 10010 366956 220116
rect 367296 217802 367324 220116
rect 367284 217796 367336 217802
rect 367284 217738 367336 217744
rect 367756 217734 367784 220116
rect 368138 220102 368244 220130
rect 367008 217728 367060 217734
rect 367008 217670 367060 217676
rect 367744 217728 367796 217734
rect 367744 217670 367796 217676
rect 367020 11082 367048 217670
rect 367098 40352 367154 40361
rect 367098 40287 367100 40296
rect 367152 40287 367154 40296
rect 367100 40258 367152 40264
rect 367100 14748 367152 14754
rect 367100 14690 367152 14696
rect 367008 11076 367060 11082
rect 367008 11018 367060 11024
rect 366928 9982 367048 10010
rect 366824 7744 366876 7750
rect 366824 7686 366876 7692
rect 367020 7682 367048 9982
rect 366916 7676 366968 7682
rect 366916 7618 366968 7624
rect 367008 7676 367060 7682
rect 367008 7618 367060 7624
rect 366732 4956 366784 4962
rect 366732 4898 366784 4904
rect 365720 4888 365772 4894
rect 365720 4830 365772 4836
rect 365628 3596 365680 3602
rect 365628 3538 365680 3544
rect 365732 400 365760 4830
rect 366928 400 366956 7618
rect 367112 542 367140 14690
rect 368216 7614 368244 220102
rect 368584 217802 368612 220116
rect 368388 217796 368440 217802
rect 368388 217738 368440 217744
rect 368572 217796 368624 217802
rect 368572 217738 368624 217744
rect 368296 217728 368348 217734
rect 368296 217670 368348 217676
rect 368204 7608 368256 7614
rect 368204 7550 368256 7556
rect 368308 4894 368336 217670
rect 368296 4888 368348 4894
rect 368296 4830 368348 4836
rect 368400 3534 368428 217738
rect 368952 217734 368980 220116
rect 369426 220102 369624 220130
rect 368940 217728 368992 217734
rect 368940 217670 368992 217676
rect 369596 7585 369624 220102
rect 369676 217728 369728 217734
rect 369676 217670 369728 217676
rect 369582 7576 369638 7585
rect 369582 7511 369638 7520
rect 369688 4826 369716 217670
rect 369216 4820 369268 4826
rect 369216 4762 369268 4768
rect 369676 4820 369728 4826
rect 369676 4762 369728 4768
rect 368388 3528 368440 3534
rect 368388 3470 368440 3476
rect 367100 536 367152 542
rect 367100 478 367152 484
rect 368020 536 368072 542
rect 368020 478 368072 484
rect 368032 400 368060 478
rect 369228 400 369256 4762
rect 369780 3466 369808 220116
rect 369952 40316 370004 40322
rect 369952 40258 370004 40264
rect 369964 40089 369992 40258
rect 369950 40080 370006 40089
rect 369950 40015 370006 40024
rect 370516 30326 370544 522543
rect 370596 520668 370648 520674
rect 370596 520610 370648 520616
rect 370608 393310 370636 520610
rect 370688 519580 370740 519586
rect 370688 519522 370740 519528
rect 370700 405686 370728 519522
rect 370792 416770 370820 522854
rect 370964 520804 371016 520810
rect 370964 520746 371016 520752
rect 370872 520736 370924 520742
rect 370872 520678 370924 520684
rect 370884 440230 370912 520678
rect 370976 452606 371004 520746
rect 371068 463690 371096 522922
rect 376024 522844 376076 522850
rect 376024 522786 376076 522792
rect 372066 518936 372122 518945
rect 372066 518871 372122 518880
rect 371882 518392 371938 518401
rect 371882 518327 371938 518336
rect 371896 518129 371924 518327
rect 372080 518129 372108 518871
rect 375286 518800 375342 518809
rect 375286 518735 375342 518744
rect 375300 518702 375328 518735
rect 375288 518696 375340 518702
rect 375288 518638 375340 518644
rect 371882 518120 371938 518129
rect 371882 518055 371938 518064
rect 372066 518120 372122 518129
rect 372066 518055 372122 518064
rect 371146 517984 371202 517993
rect 371146 517919 371202 517928
rect 371160 499526 371188 517919
rect 371148 499520 371200 499526
rect 371148 499462 371200 499468
rect 371882 486432 371938 486441
rect 371882 486367 371938 486376
rect 371896 485897 371924 486367
rect 371882 485888 371938 485897
rect 371882 485823 371938 485832
rect 371056 463684 371108 463690
rect 371056 463626 371108 463632
rect 370964 452600 371016 452606
rect 370964 452542 371016 452548
rect 370872 440224 370924 440230
rect 370872 440166 370924 440172
rect 370780 416764 370832 416770
rect 370780 416706 370832 416712
rect 370688 405680 370740 405686
rect 370688 405622 370740 405628
rect 370596 393304 370648 393310
rect 370596 393246 370648 393252
rect 376036 171086 376064 522786
rect 580814 522200 580870 522209
rect 580814 522135 580870 522144
rect 580630 522064 580686 522073
rect 580630 521999 580686 522008
rect 580446 521928 580502 521937
rect 580446 521863 580502 521872
rect 580262 521792 580318 521801
rect 580262 521727 580318 521736
rect 379426 518800 379482 518809
rect 379426 518735 379482 518744
rect 405752 518758 405872 518786
rect 379440 518650 379468 518735
rect 405752 518673 405780 518758
rect 379610 518664 379666 518673
rect 379440 518622 379610 518650
rect 379610 518599 379666 518608
rect 386418 518664 386474 518673
rect 386418 518599 386474 518608
rect 399298 518664 399354 518673
rect 399298 518599 399354 518608
rect 405738 518664 405794 518673
rect 405738 518599 405794 518608
rect 386432 517857 386460 518599
rect 399312 517857 399340 518599
rect 405844 517993 405872 518758
rect 425072 518758 425192 518786
rect 425072 518673 425100 518758
rect 418066 518664 418122 518673
rect 418066 518599 418122 518608
rect 425058 518664 425114 518673
rect 425058 518599 425114 518608
rect 418080 517993 418108 518599
rect 425164 517993 425192 518758
rect 444392 518758 444512 518786
rect 444392 518673 444420 518758
rect 437386 518664 437442 518673
rect 437386 518599 437442 518608
rect 444378 518664 444434 518673
rect 444378 518599 444434 518608
rect 437400 517993 437428 518599
rect 444484 517993 444512 518758
rect 463712 518758 463832 518786
rect 463712 518673 463740 518758
rect 456706 518664 456762 518673
rect 456706 518599 456762 518608
rect 463698 518664 463754 518673
rect 463698 518599 463754 518608
rect 456720 517993 456748 518599
rect 463804 517993 463832 518758
rect 483032 518758 483152 518786
rect 483032 518673 483060 518758
rect 476026 518664 476082 518673
rect 476026 518599 476082 518608
rect 483018 518664 483074 518673
rect 483018 518599 483074 518608
rect 476040 517993 476068 518599
rect 483124 517993 483152 518758
rect 502352 518758 502472 518786
rect 502352 518673 502380 518758
rect 495346 518664 495402 518673
rect 495346 518599 495402 518608
rect 502338 518664 502394 518673
rect 502338 518599 502394 518608
rect 495360 517993 495388 518599
rect 502444 517993 502472 518758
rect 514666 518664 514722 518673
rect 514666 518599 514722 518608
rect 553398 518664 553454 518673
rect 553398 518599 553454 518608
rect 562966 518664 563022 518673
rect 562966 518599 563022 518608
rect 580078 518664 580134 518673
rect 580078 518599 580134 518608
rect 514680 517993 514708 518599
rect 553412 517993 553440 518599
rect 562980 517993 563008 518599
rect 579802 518528 579858 518537
rect 579802 518463 579858 518472
rect 579618 518392 579674 518401
rect 579618 518327 579674 518336
rect 405830 517984 405886 517993
rect 405830 517919 405886 517928
rect 418066 517984 418122 517993
rect 418066 517919 418122 517928
rect 425150 517984 425206 517993
rect 425150 517919 425206 517928
rect 437386 517984 437442 517993
rect 437386 517919 437442 517928
rect 444470 517984 444526 517993
rect 444470 517919 444526 517928
rect 456706 517984 456762 517993
rect 456706 517919 456762 517928
rect 463790 517984 463846 517993
rect 463790 517919 463846 517928
rect 476026 517984 476082 517993
rect 476026 517919 476082 517928
rect 483110 517984 483166 517993
rect 483110 517919 483166 517928
rect 495346 517984 495402 517993
rect 495346 517919 495402 517928
rect 502430 517984 502486 517993
rect 502430 517919 502486 517928
rect 514666 517984 514722 517993
rect 514666 517919 514722 517928
rect 553398 517984 553454 517993
rect 553398 517919 553454 517928
rect 562966 517984 563022 517993
rect 562966 517919 563022 517928
rect 386418 517848 386474 517857
rect 386418 517783 386474 517792
rect 399298 517848 399354 517857
rect 399298 517783 399354 517792
rect 576858 486976 576914 486985
rect 576858 486911 576914 486920
rect 394606 486296 394662 486305
rect 394606 486231 394662 486240
rect 379610 486024 379666 486033
rect 379440 485982 379610 486010
rect 379440 485897 379468 485982
rect 379610 485959 379666 485968
rect 394620 485897 394648 486231
rect 405646 486160 405702 486169
rect 405646 486095 405702 486104
rect 405660 486062 405688 486095
rect 398748 486056 398800 486062
rect 398746 486024 398748 486033
rect 405648 486056 405700 486062
rect 398800 486024 398802 486033
rect 405648 485998 405700 486004
rect 398746 485959 398802 485968
rect 576872 485897 576900 486911
rect 379426 485888 379482 485897
rect 379426 485823 379482 485832
rect 394606 485888 394662 485897
rect 394606 485823 394662 485832
rect 576858 485888 576914 485897
rect 576858 485823 576914 485832
rect 576858 299296 576914 299305
rect 576858 299231 576914 299240
rect 576872 298217 576900 299231
rect 576858 298208 576914 298217
rect 576858 298143 576914 298152
rect 579632 275777 579660 518327
rect 579710 518120 579766 518129
rect 579710 518055 579766 518064
rect 579724 510270 579752 518055
rect 579712 510264 579764 510270
rect 579712 510206 579764 510212
rect 579618 275768 579674 275777
rect 579618 275703 579674 275712
rect 579816 263945 579844 518463
rect 579988 510604 580040 510610
rect 579988 510546 580040 510552
rect 580000 510377 580028 510546
rect 579986 510368 580042 510377
rect 579986 510303 580042 510312
rect 579988 510264 580040 510270
rect 579988 510206 580040 510212
rect 579896 499520 579948 499526
rect 579896 499462 579948 499468
rect 579908 498681 579936 499462
rect 579894 498672 579950 498681
rect 579894 498607 579950 498616
rect 579896 463684 579948 463690
rect 579896 463626 579948 463632
rect 579908 463457 579936 463626
rect 579894 463448 579950 463457
rect 579894 463383 579950 463392
rect 579896 452600 579948 452606
rect 579896 452542 579948 452548
rect 579908 451761 579936 452542
rect 579894 451752 579950 451761
rect 579894 451687 579950 451696
rect 579896 440224 579948 440230
rect 579896 440166 579948 440172
rect 579908 439929 579936 440166
rect 579894 439920 579950 439929
rect 579894 439855 579950 439864
rect 579896 416764 579948 416770
rect 579896 416706 579948 416712
rect 579908 416537 579936 416706
rect 579894 416528 579950 416537
rect 579894 416463 579950 416472
rect 579896 405680 579948 405686
rect 579896 405622 579948 405628
rect 579908 404841 579936 405622
rect 579894 404832 579950 404841
rect 579894 404767 579950 404776
rect 579896 393304 579948 393310
rect 579896 393246 579948 393252
rect 579908 393009 579936 393246
rect 579894 393000 579950 393009
rect 579894 392935 579950 392944
rect 579896 369844 579948 369850
rect 579896 369786 579948 369792
rect 579908 369617 579936 369786
rect 579894 369608 579950 369617
rect 579894 369543 579950 369552
rect 579802 263936 579858 263945
rect 579802 263871 579858 263880
rect 576858 252376 576914 252385
rect 576858 252311 576914 252320
rect 576872 251297 576900 252311
rect 576858 251288 576914 251297
rect 576858 251223 576914 251232
rect 580000 228857 580028 510206
rect 580092 357921 580120 518599
rect 580170 518256 580226 518265
rect 580170 518191 580226 518200
rect 580078 357912 580134 357921
rect 580078 357847 580134 357856
rect 580080 346384 580132 346390
rect 580080 346326 580132 346332
rect 580092 346089 580120 346326
rect 580078 346080 580134 346089
rect 580078 346015 580134 346024
rect 580080 322924 580132 322930
rect 580080 322866 580132 322872
rect 580092 322697 580120 322866
rect 580078 322688 580134 322697
rect 580078 322623 580134 322632
rect 579986 228848 580042 228857
rect 579986 228783 580042 228792
rect 469864 218000 469916 218006
rect 469864 217942 469916 217948
rect 434720 217660 434772 217666
rect 434720 217602 434772 217608
rect 427820 217252 427872 217258
rect 427820 217194 427872 217200
rect 420920 217184 420972 217190
rect 420920 217126 420972 217132
rect 414020 217116 414072 217122
rect 414020 217058 414072 217064
rect 407120 217048 407172 217054
rect 407120 216990 407172 216996
rect 400220 216980 400272 216986
rect 400220 216922 400272 216928
rect 391940 216912 391992 216918
rect 391940 216854 391992 216860
rect 385040 216844 385092 216850
rect 385040 216786 385092 216792
rect 376024 171080 376076 171086
rect 376024 171022 376076 171028
rect 379610 40216 379666 40225
rect 379440 40174 379610 40202
rect 379440 40089 379468 40174
rect 379610 40151 379666 40160
rect 379426 40080 379482 40089
rect 379426 40015 379482 40024
rect 370504 30320 370556 30326
rect 370504 30262 370556 30268
rect 371240 14680 371292 14686
rect 371240 14622 371292 14628
rect 369860 11280 369912 11286
rect 369860 11222 369912 11228
rect 369768 3460 369820 3466
rect 369768 3402 369820 3408
rect 369872 490 369900 11222
rect 371252 490 371280 14622
rect 375196 14612 375248 14618
rect 375196 14554 375248 14560
rect 374092 11348 374144 11354
rect 374092 11290 374144 11296
rect 372802 4856 372858 4865
rect 372802 4791 372858 4800
rect 369872 462 370452 490
rect 371252 462 371648 490
rect 370424 400 370452 462
rect 371620 400 371648 462
rect 372816 400 372844 4791
rect 374104 1578 374132 11290
rect 374012 1550 374132 1578
rect 374012 400 374040 1550
rect 375208 400 375236 14554
rect 378140 14544 378192 14550
rect 378140 14486 378192 14492
rect 376760 11416 376812 11422
rect 376760 11358 376812 11364
rect 375380 9920 375432 9926
rect 375380 9862 375432 9868
rect 375392 542 375420 9862
rect 376772 542 376800 11358
rect 375380 536 375432 542
rect 375380 478 375432 484
rect 376392 536 376444 542
rect 376392 478 376444 484
rect 376760 536 376812 542
rect 376760 478 376812 484
rect 377588 536 377640 542
rect 377588 478 377640 484
rect 378152 490 378180 14486
rect 383660 11552 383712 11558
rect 383660 11494 383712 11500
rect 380900 11484 380952 11490
rect 380900 11426 380952 11432
rect 379520 9988 379572 9994
rect 379520 9930 379572 9936
rect 379532 490 379560 9930
rect 380912 490 380940 11426
rect 382372 10056 382424 10062
rect 382372 9998 382424 10004
rect 382384 2922 382412 9998
rect 382280 2916 382332 2922
rect 382280 2858 382332 2864
rect 382372 2916 382424 2922
rect 382372 2858 382424 2864
rect 383568 2916 383620 2922
rect 383568 2858 383620 2864
rect 382292 2802 382320 2858
rect 382292 2774 382412 2802
rect 376404 400 376432 478
rect 377600 400 377628 478
rect 378152 462 378824 490
rect 379532 462 380020 490
rect 380912 462 381216 490
rect 378796 400 378824 462
rect 379992 400 380020 462
rect 381188 400 381216 462
rect 382384 400 382412 2774
rect 383580 400 383608 2858
rect 383672 542 383700 11494
rect 385052 542 385080 216786
rect 390560 11688 390612 11694
rect 390560 11630 390612 11636
rect 387800 11620 387852 11626
rect 387800 11562 387852 11568
rect 386420 10124 386472 10130
rect 386420 10066 386472 10072
rect 383660 536 383712 542
rect 383660 478 383712 484
rect 384672 536 384724 542
rect 384672 478 384724 484
rect 385040 536 385092 542
rect 385040 478 385092 484
rect 385868 536 385920 542
rect 385868 478 385920 484
rect 386432 490 386460 10066
rect 387812 490 387840 11562
rect 390572 2922 390600 11630
rect 390652 10192 390704 10198
rect 390652 10134 390704 10140
rect 390560 2916 390612 2922
rect 390560 2858 390612 2864
rect 389456 2848 389508 2854
rect 389456 2790 389508 2796
rect 384684 400 384712 478
rect 385880 400 385908 478
rect 386432 462 387104 490
rect 387812 462 388300 490
rect 387076 400 387104 462
rect 388272 400 388300 462
rect 389468 400 389496 2790
rect 390664 400 390692 10134
rect 391848 2916 391900 2922
rect 391848 2858 391900 2864
rect 391860 400 391888 2858
rect 391952 542 391980 216854
rect 394606 40488 394662 40497
rect 394606 40423 394662 40432
rect 394620 40089 394648 40423
rect 398748 40248 398800 40254
rect 398746 40216 398748 40225
rect 398800 40216 398802 40225
rect 398746 40151 398802 40160
rect 394606 40080 394662 40089
rect 394606 40015 394662 40024
rect 397460 11008 397512 11014
rect 397460 10950 397512 10956
rect 393320 10260 393372 10266
rect 393320 10202 393372 10208
rect 393332 3346 393360 10202
rect 395436 8356 395488 8362
rect 395436 8298 395488 8304
rect 393332 3318 394280 3346
rect 391940 536 391992 542
rect 391940 478 391992 484
rect 393044 536 393096 542
rect 393044 478 393096 484
rect 393056 400 393084 478
rect 394252 400 394280 3318
rect 395448 400 395476 8298
rect 397472 3346 397500 10950
rect 399024 8424 399076 8430
rect 399024 8366 399076 8372
rect 397472 3318 397868 3346
rect 396632 2984 396684 2990
rect 396632 2926 396684 2932
rect 396644 400 396672 2926
rect 397840 400 397868 3318
rect 399036 400 399064 8366
rect 400232 400 400260 216922
rect 405646 40352 405702 40361
rect 405646 40287 405702 40296
rect 405660 40254 405688 40287
rect 405648 40248 405700 40254
rect 405648 40190 405700 40196
rect 400312 10940 400364 10946
rect 400312 10882 400364 10888
rect 400324 3346 400352 10882
rect 406108 8560 406160 8566
rect 406108 8502 406160 8508
rect 402520 8492 402572 8498
rect 402520 8434 402572 8440
rect 400324 3318 401364 3346
rect 401336 400 401364 3318
rect 402532 400 402560 8434
rect 404912 5568 404964 5574
rect 404912 5510 404964 5516
rect 403716 3120 403768 3126
rect 403716 3062 403768 3068
rect 403728 400 403756 3062
rect 404924 400 404952 5510
rect 406120 400 406148 8502
rect 407132 3346 407160 216990
rect 413284 8696 413336 8702
rect 413284 8638 413336 8644
rect 409696 8628 409748 8634
rect 409696 8570 409748 8576
rect 408500 5636 408552 5642
rect 408500 5578 408552 5584
rect 407132 3318 407344 3346
rect 407316 400 407344 3318
rect 408512 400 408540 5578
rect 409708 400 409736 8570
rect 412088 5704 412140 5710
rect 412088 5646 412140 5652
rect 410892 3188 410944 3194
rect 410892 3130 410944 3136
rect 410904 400 410932 3130
rect 412100 400 412128 5646
rect 413296 400 413324 8638
rect 414032 3346 414060 217058
rect 420368 8832 420420 8838
rect 420368 8774 420420 8780
rect 416872 8764 416924 8770
rect 416872 8706 416924 8712
rect 415676 5772 415728 5778
rect 415676 5714 415728 5720
rect 414032 3318 414520 3346
rect 414492 400 414520 3318
rect 415688 400 415716 5714
rect 416884 400 416912 8706
rect 419172 5840 419224 5846
rect 419172 5782 419224 5788
rect 417976 3324 418028 3330
rect 417976 3266 418028 3272
rect 417988 400 418016 3266
rect 419184 400 419212 5782
rect 420380 400 420408 8774
rect 420932 3346 420960 217126
rect 427544 9648 427596 9654
rect 427544 9590 427596 9596
rect 423956 8900 424008 8906
rect 423956 8842 424008 8848
rect 422760 5908 422812 5914
rect 422760 5850 422812 5856
rect 420932 3318 421604 3346
rect 421576 400 421604 3318
rect 422772 400 422800 5850
rect 423968 400 423996 8842
rect 426348 5976 426400 5982
rect 426348 5918 426400 5924
rect 425152 3256 425204 3262
rect 425152 3198 425204 3204
rect 425164 400 425192 3198
rect 426360 400 426388 5918
rect 427556 400 427584 9590
rect 427832 3346 427860 217194
rect 431132 9580 431184 9586
rect 431132 9522 431184 9528
rect 429936 6044 429988 6050
rect 429936 5986 429988 5992
rect 427832 3318 428780 3346
rect 428752 400 428780 3318
rect 429948 400 429976 5986
rect 431144 400 431172 9522
rect 434628 9512 434680 9518
rect 434628 9454 434680 9460
rect 433524 6112 433576 6118
rect 433524 6054 433576 6060
rect 432328 3052 432380 3058
rect 432328 2994 432380 3000
rect 432340 400 432368 2994
rect 433536 400 433564 6054
rect 434640 400 434668 9454
rect 434732 3346 434760 217602
rect 443000 217592 443052 217598
rect 443000 217534 443052 217540
rect 438216 9444 438268 9450
rect 438216 9386 438268 9392
rect 437020 6860 437072 6866
rect 437020 6802 437072 6808
rect 434732 3318 435864 3346
rect 435836 400 435864 3318
rect 437032 400 437060 6802
rect 438228 400 438256 9386
rect 441804 9376 441856 9382
rect 441804 9318 441856 9324
rect 440608 6792 440660 6798
rect 440608 6734 440660 6740
rect 439412 4004 439464 4010
rect 439412 3946 439464 3952
rect 439424 400 439452 3946
rect 440620 400 440648 6734
rect 441816 400 441844 9318
rect 443012 400 443040 217534
rect 449900 217524 449952 217530
rect 449900 217466 449952 217472
rect 445392 9308 445444 9314
rect 445392 9250 445444 9256
rect 444196 6724 444248 6730
rect 444196 6666 444248 6672
rect 444208 400 444236 6666
rect 445404 400 445432 9250
rect 448980 9240 449032 9246
rect 448980 9182 449032 9188
rect 447784 6656 447836 6662
rect 447784 6598 447836 6604
rect 446588 3392 446640 3398
rect 446588 3334 446640 3340
rect 446600 400 446628 3334
rect 447796 400 447824 6598
rect 448992 400 449020 9182
rect 449912 3482 449940 217466
rect 456800 217456 456852 217462
rect 456800 217398 456852 217404
rect 452476 9172 452528 9178
rect 452476 9114 452528 9120
rect 451280 6588 451332 6594
rect 451280 6530 451332 6536
rect 449912 3454 450216 3482
rect 450188 400 450216 3454
rect 451292 400 451320 6530
rect 452488 400 452516 9114
rect 456064 9104 456116 9110
rect 456064 9046 456116 9052
rect 454868 6520 454920 6526
rect 454868 6462 454920 6468
rect 453672 4072 453724 4078
rect 453672 4014 453724 4020
rect 453684 400 453712 4014
rect 454880 400 454908 6462
rect 456076 400 456104 9046
rect 456812 3346 456840 217398
rect 463700 217388 463752 217394
rect 463700 217330 463752 217336
rect 459652 9036 459704 9042
rect 459652 8978 459704 8984
rect 458456 6452 458508 6458
rect 458456 6394 458508 6400
rect 456812 3318 457300 3346
rect 457272 400 457300 3318
rect 458468 400 458496 6394
rect 459664 400 459692 8978
rect 463240 8968 463292 8974
rect 463240 8910 463292 8916
rect 462044 6384 462096 6390
rect 462044 6326 462096 6332
rect 460848 4140 460900 4146
rect 460848 4082 460900 4088
rect 460860 400 460888 4082
rect 462056 400 462084 6326
rect 463252 400 463280 8910
rect 463712 542 463740 217330
rect 469220 12436 469272 12442
rect 469220 12378 469272 12384
rect 466826 8936 466882 8945
rect 466826 8871 466882 8880
rect 465632 6316 465684 6322
rect 465632 6258 465684 6264
rect 463700 536 463752 542
rect 463700 478 463752 484
rect 464436 536 464488 542
rect 464436 478 464488 484
rect 464448 400 464476 478
rect 465644 400 465672 6258
rect 466840 400 466868 8871
rect 469128 6248 469180 6254
rect 469128 6190 469180 6196
rect 467932 3936 467984 3942
rect 467932 3878 467984 3884
rect 467944 400 467972 3878
rect 469140 400 469168 6190
rect 469232 3346 469260 12378
rect 469876 4146 469904 217942
rect 478144 217932 478196 217938
rect 478144 217874 478196 217880
rect 475384 217864 475436 217870
rect 475384 217806 475436 217812
rect 474004 217728 474056 217734
rect 474004 217670 474056 217676
rect 470598 217288 470654 217297
rect 470598 217223 470654 217232
rect 469864 4140 469916 4146
rect 469864 4082 469916 4088
rect 469232 3318 470364 3346
rect 470336 400 470364 3318
rect 470612 490 470640 217223
rect 473360 12368 473412 12374
rect 473360 12310 473412 12316
rect 472716 6180 472768 6186
rect 472716 6122 472768 6128
rect 470612 462 471560 490
rect 471532 400 471560 462
rect 472728 400 472756 6122
rect 473372 490 473400 12310
rect 474016 4078 474044 217670
rect 474004 4072 474056 4078
rect 474004 4014 474056 4020
rect 475396 4010 475424 217806
rect 477500 217320 477552 217326
rect 477500 217262 477552 217268
rect 476302 6216 476358 6225
rect 476302 6151 476358 6160
rect 475384 4004 475436 4010
rect 475384 3946 475436 3952
rect 475108 3868 475160 3874
rect 475108 3810 475160 3816
rect 473372 462 473952 490
rect 473924 400 473952 462
rect 475120 400 475148 3810
rect 476316 400 476344 6151
rect 477512 3874 477540 217262
rect 477592 12708 477644 12714
rect 477592 12650 477644 12656
rect 477500 3868 477552 3874
rect 477500 3810 477552 3816
rect 477604 3482 477632 12650
rect 478156 3942 478184 217874
rect 480904 217796 480956 217802
rect 480904 217738 480956 217744
rect 480260 12776 480312 12782
rect 480260 12718 480312 12724
rect 478880 12300 478932 12306
rect 478880 12242 478932 12248
rect 478144 3936 478196 3942
rect 478144 3878 478196 3884
rect 478696 3868 478748 3874
rect 478696 3810 478748 3816
rect 477512 3454 477632 3482
rect 477512 400 477540 3454
rect 478708 400 478736 3810
rect 478892 542 478920 12242
rect 480272 3346 480300 12718
rect 480916 3874 480944 217738
rect 580184 217025 580212 518191
rect 580170 217016 580226 217025
rect 580170 216951 580226 216960
rect 576858 205456 576914 205465
rect 576858 205391 576914 205400
rect 576872 204377 576900 205391
rect 576858 204368 576914 204377
rect 576858 204303 576914 204312
rect 580172 171080 580224 171086
rect 580172 171022 580224 171028
rect 580184 170105 580212 171022
rect 580170 170096 580226 170105
rect 580170 170031 580226 170040
rect 580276 64569 580304 521727
rect 580356 518220 580408 518226
rect 580356 518162 580408 518168
rect 580368 76265 580396 518162
rect 580460 87961 580488 521863
rect 580540 520328 580592 520334
rect 580540 520270 580592 520276
rect 580552 134881 580580 520270
rect 580538 134872 580594 134881
rect 580538 134807 580594 134816
rect 580644 111489 580672 521999
rect 580724 521688 580776 521694
rect 580724 521630 580776 521636
rect 580736 158409 580764 521630
rect 580722 158400 580778 158409
rect 580722 158335 580778 158344
rect 580828 123185 580856 522135
rect 580908 520396 580960 520402
rect 580908 520338 580960 520344
rect 580920 181937 580948 520338
rect 583390 486976 583446 486985
rect 583390 486911 583446 486920
rect 583404 486849 583432 486911
rect 583390 486840 583446 486849
rect 583390 486775 583446 486784
rect 583390 310856 583446 310865
rect 583390 310791 583446 310800
rect 583404 310729 583432 310791
rect 583390 310720 583446 310729
rect 583390 310655 583446 310664
rect 583390 299296 583446 299305
rect 583390 299231 583446 299240
rect 583404 299169 583432 299231
rect 583390 299160 583446 299169
rect 583390 299095 583446 299104
rect 583390 252376 583446 252385
rect 583390 252311 583446 252320
rect 583404 252249 583432 252311
rect 583390 252240 583446 252249
rect 583390 252175 583446 252184
rect 583390 205456 583446 205465
rect 583390 205391 583446 205400
rect 583404 205329 583432 205391
rect 583390 205320 583446 205329
rect 583390 205255 583446 205264
rect 580906 181928 580962 181937
rect 580906 181863 580962 181872
rect 580814 123176 580870 123185
rect 580814 123111 580870 123120
rect 580630 111480 580686 111489
rect 580630 111415 580686 111424
rect 580446 87952 580502 87961
rect 580446 87887 580502 87896
rect 580354 76256 580410 76265
rect 580354 76191 580410 76200
rect 580262 64560 580318 64569
rect 580262 64495 580318 64504
rect 576858 41168 576914 41177
rect 576858 41103 576914 41112
rect 583390 41168 583446 41177
rect 583390 41103 583446 41112
rect 576872 40089 576900 41103
rect 583404 41041 583432 41103
rect 583390 41032 583446 41041
rect 583390 40967 583446 40976
rect 576858 40080 576914 40089
rect 576858 40015 576914 40024
rect 580264 30320 580316 30326
rect 580264 30262 580316 30268
rect 580276 29345 580304 30262
rect 580262 29336 580318 29345
rect 580262 29271 580318 29280
rect 579620 17944 579672 17950
rect 579620 17886 579672 17892
rect 579632 17649 579660 17886
rect 579618 17640 579674 17649
rect 579618 17575 579674 17584
rect 546500 14476 546552 14482
rect 546500 14418 546552 14424
rect 499580 13796 499632 13802
rect 499580 13738 499632 13744
rect 495440 13048 495492 13054
rect 495440 12990 495492 12996
rect 492680 12980 492732 12986
rect 492680 12922 492732 12928
rect 488540 12912 488592 12918
rect 488540 12854 488592 12860
rect 485780 12844 485832 12850
rect 485780 12786 485832 12792
rect 484400 12232 484452 12238
rect 484400 12174 484452 12180
rect 483020 10872 483072 10878
rect 483020 10814 483072 10820
rect 480904 3868 480956 3874
rect 480904 3810 480956 3816
rect 482284 3800 482336 3806
rect 482284 3742 482336 3748
rect 480272 3318 481128 3346
rect 478880 536 478932 542
rect 478880 478 478932 484
rect 479892 536 479944 542
rect 479892 478 479944 484
rect 479904 400 479932 478
rect 481100 400 481128 3318
rect 482296 400 482324 3742
rect 483032 490 483060 10814
rect 484412 490 484440 12174
rect 483032 462 483520 490
rect 484412 462 484624 490
rect 483492 400 483520 462
rect 484596 400 484624 462
rect 485792 400 485820 12786
rect 487160 12164 487212 12170
rect 487160 12106 487212 12112
rect 485872 10804 485924 10810
rect 485872 10746 485924 10752
rect 485884 542 485912 10746
rect 487172 542 487200 12106
rect 485872 536 485924 542
rect 485872 478 485924 484
rect 486976 536 487028 542
rect 486976 478 487028 484
rect 487160 536 487212 542
rect 487160 478 487212 484
rect 488172 536 488224 542
rect 488172 478 488224 484
rect 488552 490 488580 12854
rect 491300 12096 491352 12102
rect 491300 12038 491352 12044
rect 489920 10736 489972 10742
rect 489920 10678 489972 10684
rect 489932 542 489960 10678
rect 489920 536 489972 542
rect 486988 400 487016 478
rect 488184 400 488212 478
rect 488552 462 489408 490
rect 489920 478 489972 484
rect 490564 536 490616 542
rect 490564 478 490616 484
rect 491312 490 491340 12038
rect 492692 490 492720 12922
rect 494060 12028 494112 12034
rect 494060 11970 494112 11976
rect 494072 3398 494100 11970
rect 494152 10668 494204 10674
rect 494152 10610 494204 10616
rect 494060 3392 494112 3398
rect 494060 3334 494112 3340
rect 489380 400 489408 462
rect 490576 400 490604 478
rect 491312 462 491800 490
rect 492692 462 492996 490
rect 491772 400 491800 462
rect 492968 400 492996 462
rect 494164 400 494192 10610
rect 495348 3392 495400 3398
rect 495348 3334 495400 3340
rect 495360 400 495388 3334
rect 495452 542 495480 12990
rect 498200 11960 498252 11966
rect 498200 11902 498252 11908
rect 496820 10600 496872 10606
rect 496820 10542 496872 10548
rect 496832 542 496860 10542
rect 495440 536 495492 542
rect 495440 478 495492 484
rect 496544 536 496596 542
rect 496544 478 496596 484
rect 496820 536 496872 542
rect 496820 478 496872 484
rect 497740 536 497792 542
rect 497740 478 497792 484
rect 498212 490 498240 11902
rect 499592 3346 499620 13738
rect 502340 13728 502392 13734
rect 502340 13670 502392 13676
rect 500960 10532 501012 10538
rect 500960 10474 501012 10480
rect 500972 3346 501000 10474
rect 502352 3398 502380 13670
rect 506480 13660 506532 13666
rect 506480 13602 506532 13608
rect 502432 11892 502484 11898
rect 502432 11834 502484 11840
rect 502340 3392 502392 3398
rect 499592 3318 500172 3346
rect 500972 3318 501276 3346
rect 502340 3334 502392 3340
rect 496556 400 496584 478
rect 497752 400 497780 478
rect 498212 462 498976 490
rect 498948 400 498976 462
rect 500144 400 500172 3318
rect 501248 400 501276 3318
rect 502444 400 502472 11834
rect 505100 11824 505152 11830
rect 505100 11766 505152 11772
rect 503720 10464 503772 10470
rect 503720 10406 503772 10412
rect 503628 3392 503680 3398
rect 503628 3334 503680 3340
rect 503732 3346 503760 10406
rect 505112 3346 505140 11766
rect 506492 3346 506520 13602
rect 510620 13592 510672 13598
rect 510620 13534 510672 13540
rect 507860 10396 507912 10402
rect 507860 10338 507912 10344
rect 507872 3346 507900 10338
rect 509608 6996 509660 7002
rect 509608 6938 509660 6944
rect 503640 400 503668 3334
rect 503732 3318 504864 3346
rect 505112 3318 506060 3346
rect 506492 3318 507256 3346
rect 507872 3318 508452 3346
rect 504836 400 504864 3318
rect 506032 400 506060 3318
rect 507228 400 507256 3318
rect 508424 400 508452 3318
rect 509620 400 509648 6938
rect 510632 3482 510660 13534
rect 517520 13524 517572 13530
rect 517520 13466 517572 13472
rect 513380 10328 513432 10334
rect 513380 10270 513432 10276
rect 513196 7064 513248 7070
rect 513196 7006 513248 7012
rect 512000 4208 512052 4214
rect 512000 4150 512052 4156
rect 510632 3454 510844 3482
rect 510816 400 510844 3454
rect 512012 400 512040 4150
rect 513208 400 513236 7006
rect 513392 3482 513420 10270
rect 516784 7132 516836 7138
rect 516784 7074 516836 7080
rect 515588 4276 515640 4282
rect 515588 4218 515640 4224
rect 513392 3454 514432 3482
rect 514404 400 514432 3454
rect 515600 400 515628 4218
rect 516796 400 516824 7074
rect 517532 3482 517560 13466
rect 520280 13456 520332 13462
rect 520280 13398 520332 13404
rect 519084 4344 519136 4350
rect 519084 4286 519136 4292
rect 517532 3454 517928 3482
rect 517900 400 517928 3454
rect 519096 400 519124 4286
rect 520292 3806 520320 13398
rect 524420 13388 524472 13394
rect 524420 13330 524472 13336
rect 523868 7268 523920 7274
rect 523868 7210 523920 7216
rect 520372 7200 520424 7206
rect 520372 7142 520424 7148
rect 520280 3800 520332 3806
rect 520280 3742 520332 3748
rect 520384 3482 520412 7142
rect 522672 4412 522724 4418
rect 522672 4354 522724 4360
rect 521476 3800 521528 3806
rect 521476 3742 521528 3748
rect 520292 3454 520412 3482
rect 520292 400 520320 3454
rect 521488 400 521516 3742
rect 522684 400 522712 4354
rect 523880 400 523908 7210
rect 524432 490 524460 13330
rect 528560 13320 528612 13326
rect 528560 13262 528612 13268
rect 527456 7336 527508 7342
rect 527456 7278 527508 7284
rect 526260 4480 526312 4486
rect 526260 4422 526312 4428
rect 524432 462 525104 490
rect 525076 400 525104 462
rect 526272 400 526300 4422
rect 527468 400 527496 7278
rect 528572 490 528600 13262
rect 535460 13252 535512 13258
rect 535460 13194 535512 13200
rect 531320 11756 531372 11762
rect 531320 11698 531372 11704
rect 531044 7404 531096 7410
rect 531044 7346 531096 7352
rect 529848 4548 529900 4554
rect 529848 4490 529900 4496
rect 528572 462 528692 490
rect 528664 400 528692 462
rect 529860 400 529888 4490
rect 531056 400 531084 7346
rect 531332 490 531360 11698
rect 534540 7472 534592 7478
rect 534540 7414 534592 7420
rect 533436 4616 533488 4622
rect 533436 4558 533488 4564
rect 531332 462 532280 490
rect 532252 400 532280 462
rect 533448 400 533476 4558
rect 534552 400 534580 7414
rect 535472 490 535500 13194
rect 538220 13184 538272 13190
rect 538220 13126 538272 13132
rect 538128 7540 538180 7546
rect 538128 7482 538180 7488
rect 536932 4684 536984 4690
rect 536932 4626 536984 4632
rect 535472 462 535776 490
rect 535748 400 535776 462
rect 536944 400 536972 4626
rect 538140 400 538168 7482
rect 538232 542 538260 13126
rect 542360 13116 542412 13122
rect 542360 13058 542412 13064
rect 541716 8288 541768 8294
rect 541716 8230 541768 8236
rect 540520 4752 540572 4758
rect 540520 4694 540572 4700
rect 538220 536 538272 542
rect 538220 478 538272 484
rect 539324 536 539376 542
rect 539324 478 539376 484
rect 539336 400 539364 478
rect 540532 400 540560 4694
rect 541728 400 541756 8230
rect 542372 490 542400 13058
rect 545304 8220 545356 8226
rect 545304 8162 545356 8168
rect 544108 5500 544160 5506
rect 544108 5442 544160 5448
rect 542372 462 542952 490
rect 542924 400 542952 462
rect 544120 400 544148 5442
rect 545316 400 545344 8162
rect 546512 400 546540 14418
rect 548892 8152 548944 8158
rect 548892 8094 548944 8100
rect 547696 5432 547748 5438
rect 547696 5374 547748 5380
rect 547708 400 547736 5374
rect 548904 400 548932 8094
rect 552388 8084 552440 8090
rect 552388 8026 552440 8032
rect 551192 5364 551244 5370
rect 551192 5306 551244 5312
rect 550088 4140 550140 4146
rect 550088 4082 550140 4088
rect 550100 400 550128 4082
rect 551204 400 551232 5306
rect 552400 400 552428 8026
rect 555976 8016 556028 8022
rect 555976 7958 556028 7964
rect 554780 5296 554832 5302
rect 554780 5238 554832 5244
rect 553584 3732 553636 3738
rect 553584 3674 553636 3680
rect 553596 400 553624 3674
rect 554792 400 554820 5238
rect 555988 400 556016 7958
rect 559564 7948 559616 7954
rect 559564 7890 559616 7896
rect 558368 5228 558420 5234
rect 558368 5170 558420 5176
rect 557172 4072 557224 4078
rect 557172 4014 557224 4020
rect 557184 400 557212 4014
rect 558380 400 558408 5170
rect 559576 400 559604 7890
rect 563152 7880 563204 7886
rect 563152 7822 563204 7828
rect 561956 5160 562008 5166
rect 561956 5102 562008 5108
rect 560760 3664 560812 3670
rect 560760 3606 560812 3612
rect 560772 400 560800 3606
rect 561968 400 561996 5102
rect 563164 400 563192 7822
rect 566740 7812 566792 7818
rect 566740 7754 566792 7760
rect 565544 5092 565596 5098
rect 565544 5034 565596 5040
rect 564348 4004 564400 4010
rect 564348 3946 564400 3952
rect 564360 400 564388 3946
rect 565556 400 565584 5034
rect 566752 400 566780 7754
rect 570236 7744 570288 7750
rect 570236 7686 570288 7692
rect 569040 5024 569092 5030
rect 569040 4966 569092 4972
rect 567844 3596 567896 3602
rect 567844 3538 567896 3544
rect 567856 400 567884 3538
rect 569052 400 569080 4966
rect 570248 400 570276 7686
rect 573824 7676 573876 7682
rect 573824 7618 573876 7624
rect 572628 4956 572680 4962
rect 572628 4898 572680 4904
rect 571432 3936 571484 3942
rect 571432 3878 571484 3884
rect 571444 400 571472 3878
rect 572640 400 572668 4898
rect 573836 400 573864 7618
rect 577412 7608 577464 7614
rect 577412 7550 577464 7556
rect 580998 7576 581054 7585
rect 576216 4888 576268 4894
rect 576216 4830 576268 4836
rect 575020 3528 575072 3534
rect 575020 3470 575072 3476
rect 575032 400 575060 3470
rect 576228 400 576256 4830
rect 577424 400 577452 7550
rect 580998 7511 581054 7520
rect 579804 4820 579856 4826
rect 579804 4762 579856 4768
rect 578608 3868 578660 3874
rect 578608 3810 578660 3816
rect 578620 400 578648 3810
rect 579816 400 579844 4762
rect 581012 400 581040 7511
rect 582196 3460 582248 3466
rect 582196 3402 582248 3408
rect 582208 400 582236 3402
rect 542 -800 654 400
rect 1646 -800 1758 400
rect 2842 -800 2954 400
rect 4038 -800 4150 400
rect 5234 -800 5346 400
rect 6430 -800 6542 400
rect 7626 -800 7738 400
rect 8822 -800 8934 400
rect 10018 -800 10130 400
rect 11214 -800 11326 400
rect 12410 -800 12522 400
rect 13606 -800 13718 400
rect 14802 -800 14914 400
rect 15998 -800 16110 400
rect 17194 -800 17306 400
rect 18298 -800 18410 400
rect 19494 -800 19606 400
rect 20690 -800 20802 400
rect 21886 -800 21998 400
rect 23082 -800 23194 400
rect 24278 -800 24390 400
rect 25474 -800 25586 400
rect 26670 -800 26782 400
rect 27866 -800 27978 400
rect 29062 -800 29174 400
rect 30258 -800 30370 400
rect 31454 -800 31566 400
rect 32650 -800 32762 400
rect 33846 -800 33958 400
rect 34950 -800 35062 400
rect 36146 -800 36258 400
rect 37342 -800 37454 400
rect 38538 -800 38650 400
rect 39734 -800 39846 400
rect 40930 -800 41042 400
rect 42126 -800 42238 400
rect 43322 -800 43434 400
rect 44518 -800 44630 400
rect 45714 -800 45826 400
rect 46910 -800 47022 400
rect 48106 -800 48218 400
rect 49302 -800 49414 400
rect 50498 -800 50610 400
rect 51602 -800 51714 400
rect 52798 -800 52910 400
rect 53994 -800 54106 400
rect 55190 -800 55302 400
rect 56386 -800 56498 400
rect 57582 -800 57694 400
rect 58778 -800 58890 400
rect 59974 -800 60086 400
rect 61170 -800 61282 400
rect 62366 -800 62478 400
rect 63562 -800 63674 400
rect 64758 -800 64870 400
rect 65954 -800 66066 400
rect 67150 -800 67262 400
rect 68254 -800 68366 400
rect 69450 -800 69562 400
rect 70646 -800 70758 400
rect 71842 -800 71954 400
rect 73038 -800 73150 400
rect 74234 -800 74346 400
rect 75430 -800 75542 400
rect 76626 -800 76738 400
rect 77822 -800 77934 400
rect 79018 -800 79130 400
rect 80214 -800 80326 400
rect 81410 -800 81522 400
rect 82606 -800 82718 400
rect 83802 -800 83914 400
rect 84906 -800 85018 400
rect 86102 -800 86214 400
rect 87298 -800 87410 400
rect 88494 -800 88606 400
rect 89690 -800 89802 400
rect 90886 -800 90998 400
rect 92082 -800 92194 400
rect 93278 -800 93390 400
rect 94474 -800 94586 400
rect 95670 -800 95782 400
rect 96866 -800 96978 400
rect 98062 -800 98174 400
rect 99258 -800 99370 400
rect 100454 -800 100566 400
rect 101558 -800 101670 400
rect 102754 -800 102866 400
rect 103950 -800 104062 400
rect 105146 -800 105258 400
rect 106342 -800 106454 400
rect 107538 -800 107650 400
rect 108734 -800 108846 400
rect 109930 -800 110042 400
rect 111126 -800 111238 400
rect 112322 -800 112434 400
rect 113518 -800 113630 400
rect 114714 -800 114826 400
rect 115910 -800 116022 400
rect 117106 -800 117218 400
rect 118210 -800 118322 400
rect 119406 -800 119518 400
rect 120602 -800 120714 400
rect 121798 -800 121910 400
rect 122994 -800 123106 400
rect 124190 -800 124302 400
rect 125386 -800 125498 400
rect 126582 -800 126694 400
rect 127778 -800 127890 400
rect 128974 -800 129086 400
rect 130170 -800 130282 400
rect 131366 -800 131478 400
rect 132562 -800 132674 400
rect 133758 -800 133870 400
rect 134862 -800 134974 400
rect 136058 -800 136170 400
rect 137254 -800 137366 400
rect 138450 -800 138562 400
rect 139646 -800 139758 400
rect 140842 -800 140954 400
rect 142038 -800 142150 400
rect 143234 -800 143346 400
rect 144430 -800 144542 400
rect 145626 -800 145738 400
rect 146822 -800 146934 400
rect 148018 -800 148130 400
rect 149214 -800 149326 400
rect 150410 -800 150522 400
rect 151514 -800 151626 400
rect 152710 -800 152822 400
rect 153906 -800 154018 400
rect 155102 -800 155214 400
rect 156298 -800 156410 400
rect 157494 -800 157606 400
rect 158690 -800 158802 400
rect 159886 -800 159998 400
rect 161082 -800 161194 400
rect 162278 -800 162390 400
rect 163474 -800 163586 400
rect 164670 -800 164782 400
rect 165866 -800 165978 400
rect 167062 -800 167174 400
rect 168166 -800 168278 400
rect 169362 -800 169474 400
rect 170558 -800 170670 400
rect 171754 -800 171866 400
rect 172950 -800 173062 400
rect 174146 -800 174258 400
rect 175342 -800 175454 400
rect 176538 -800 176650 400
rect 177734 -800 177846 400
rect 178930 -800 179042 400
rect 180126 -800 180238 400
rect 181322 -800 181434 400
rect 182518 -800 182630 400
rect 183714 -800 183826 400
rect 184818 -800 184930 400
rect 186014 -800 186126 400
rect 187210 -800 187322 400
rect 188406 -800 188518 400
rect 189602 -800 189714 400
rect 190798 -800 190910 400
rect 191994 -800 192106 400
rect 193190 -800 193302 400
rect 194386 -800 194498 400
rect 195582 -800 195694 400
rect 196778 -800 196890 400
rect 197974 -800 198086 400
rect 199170 -800 199282 400
rect 200366 -800 200478 400
rect 201470 -800 201582 400
rect 202666 -800 202778 400
rect 203862 -800 203974 400
rect 205058 -800 205170 400
rect 206254 -800 206366 400
rect 207450 -800 207562 400
rect 208646 -800 208758 400
rect 209842 -800 209954 400
rect 211038 -800 211150 400
rect 212234 -800 212346 400
rect 213430 -800 213542 400
rect 214626 -800 214738 400
rect 215822 -800 215934 400
rect 217018 -800 217130 400
rect 218122 -800 218234 400
rect 219318 -800 219430 400
rect 220514 -800 220626 400
rect 221710 -800 221822 400
rect 222906 -800 223018 400
rect 224102 -800 224214 400
rect 225298 -800 225410 400
rect 226494 -800 226606 400
rect 227690 -800 227802 400
rect 228886 -800 228998 400
rect 230082 -800 230194 400
rect 231278 -800 231390 400
rect 232474 -800 232586 400
rect 233670 -800 233782 400
rect 234774 -800 234886 400
rect 235970 -800 236082 400
rect 237166 -800 237278 400
rect 238362 -800 238474 400
rect 239558 -800 239670 400
rect 240754 -800 240866 400
rect 241950 -800 242062 400
rect 243146 -800 243258 400
rect 244342 -800 244454 400
rect 245538 -800 245650 400
rect 246734 -800 246846 400
rect 247930 -800 248042 400
rect 249126 -800 249238 400
rect 250322 -800 250434 400
rect 251426 -800 251538 400
rect 252622 -800 252734 400
rect 253818 -800 253930 400
rect 255014 -800 255126 400
rect 256210 -800 256322 400
rect 257406 -800 257518 400
rect 258602 -800 258714 400
rect 259798 -800 259910 400
rect 260994 -800 261106 400
rect 262190 -800 262302 400
rect 263386 -800 263498 400
rect 264582 -800 264694 400
rect 265778 -800 265890 400
rect 266974 -800 267086 400
rect 268078 -800 268190 400
rect 269274 -800 269386 400
rect 270470 -800 270582 400
rect 271666 -800 271778 400
rect 272862 -800 272974 400
rect 274058 -800 274170 400
rect 275254 -800 275366 400
rect 276450 -800 276562 400
rect 277646 -800 277758 400
rect 278842 -800 278954 400
rect 280038 -800 280150 400
rect 281234 -800 281346 400
rect 282430 -800 282542 400
rect 283626 -800 283738 400
rect 284730 -800 284842 400
rect 285926 -800 286038 400
rect 287122 -800 287234 400
rect 288318 -800 288430 400
rect 289514 -800 289626 400
rect 290710 -800 290822 400
rect 291906 -800 292018 400
rect 293102 -800 293214 400
rect 294298 -800 294410 400
rect 295494 -800 295606 400
rect 296690 -800 296802 400
rect 297886 -800 297998 400
rect 299082 -800 299194 400
rect 300278 -800 300390 400
rect 301382 -800 301494 400
rect 302578 -800 302690 400
rect 303774 -800 303886 400
rect 304970 -800 305082 400
rect 306166 -800 306278 400
rect 307362 -800 307474 400
rect 308558 -800 308670 400
rect 309754 -800 309866 400
rect 310950 -800 311062 400
rect 312146 -800 312258 400
rect 313342 -800 313454 400
rect 314538 -800 314650 400
rect 315734 -800 315846 400
rect 316930 -800 317042 400
rect 318034 -800 318146 400
rect 319230 -800 319342 400
rect 320426 -800 320538 400
rect 321622 -800 321734 400
rect 322818 -800 322930 400
rect 324014 -800 324126 400
rect 325210 -800 325322 400
rect 326406 -800 326518 400
rect 327602 -800 327714 400
rect 328798 -800 328910 400
rect 329994 -800 330106 400
rect 331190 -800 331302 400
rect 332386 -800 332498 400
rect 333582 -800 333694 400
rect 334686 -800 334798 400
rect 335882 -800 335994 400
rect 337078 -800 337190 400
rect 338274 -800 338386 400
rect 339470 -800 339582 400
rect 340666 -800 340778 400
rect 341862 -800 341974 400
rect 343058 -800 343170 400
rect 344254 -800 344366 400
rect 345450 -800 345562 400
rect 346646 -800 346758 400
rect 347842 -800 347954 400
rect 349038 -800 349150 400
rect 350234 -800 350346 400
rect 351338 -800 351450 400
rect 352534 -800 352646 400
rect 353730 -800 353842 400
rect 354926 -800 355038 400
rect 356122 -800 356234 400
rect 357318 -800 357430 400
rect 358514 -800 358626 400
rect 359710 -800 359822 400
rect 360906 -800 361018 400
rect 362102 -800 362214 400
rect 363298 -800 363410 400
rect 364494 -800 364606 400
rect 365690 -800 365802 400
rect 366886 -800 366998 400
rect 367990 -800 368102 400
rect 369186 -800 369298 400
rect 370382 -800 370494 400
rect 371578 -800 371690 400
rect 372774 -800 372886 400
rect 373970 -800 374082 400
rect 375166 -800 375278 400
rect 376362 -800 376474 400
rect 377558 -800 377670 400
rect 378754 -800 378866 400
rect 379950 -800 380062 400
rect 381146 -800 381258 400
rect 382342 -800 382454 400
rect 383538 -800 383650 400
rect 384642 -800 384754 400
rect 385838 -800 385950 400
rect 387034 -800 387146 400
rect 388230 -800 388342 400
rect 389426 -800 389538 400
rect 390622 -800 390734 400
rect 391818 -800 391930 400
rect 393014 -800 393126 400
rect 394210 -800 394322 400
rect 395406 -800 395518 400
rect 396602 -800 396714 400
rect 397798 -800 397910 400
rect 398994 -800 399106 400
rect 400190 -800 400302 400
rect 401294 -800 401406 400
rect 402490 -800 402602 400
rect 403686 -800 403798 400
rect 404882 -800 404994 400
rect 406078 -800 406190 400
rect 407274 -800 407386 400
rect 408470 -800 408582 400
rect 409666 -800 409778 400
rect 410862 -800 410974 400
rect 412058 -800 412170 400
rect 413254 -800 413366 400
rect 414450 -800 414562 400
rect 415646 -800 415758 400
rect 416842 -800 416954 400
rect 417946 -800 418058 400
rect 419142 -800 419254 400
rect 420338 -800 420450 400
rect 421534 -800 421646 400
rect 422730 -800 422842 400
rect 423926 -800 424038 400
rect 425122 -800 425234 400
rect 426318 -800 426430 400
rect 427514 -800 427626 400
rect 428710 -800 428822 400
rect 429906 -800 430018 400
rect 431102 -800 431214 400
rect 432298 -800 432410 400
rect 433494 -800 433606 400
rect 434598 -800 434710 400
rect 435794 -800 435906 400
rect 436990 -800 437102 400
rect 438186 -800 438298 400
rect 439382 -800 439494 400
rect 440578 -800 440690 400
rect 441774 -800 441886 400
rect 442970 -800 443082 400
rect 444166 -800 444278 400
rect 445362 -800 445474 400
rect 446558 -800 446670 400
rect 447754 -800 447866 400
rect 448950 -800 449062 400
rect 450146 -800 450258 400
rect 451250 -800 451362 400
rect 452446 -800 452558 400
rect 453642 -800 453754 400
rect 454838 -800 454950 400
rect 456034 -800 456146 400
rect 457230 -800 457342 400
rect 458426 -800 458538 400
rect 459622 -800 459734 400
rect 460818 -800 460930 400
rect 462014 -800 462126 400
rect 463210 -800 463322 400
rect 464406 -800 464518 400
rect 465602 -800 465714 400
rect 466798 -800 466910 400
rect 467902 -800 468014 400
rect 469098 -800 469210 400
rect 470294 -800 470406 400
rect 471490 -800 471602 400
rect 472686 -800 472798 400
rect 473882 -800 473994 400
rect 475078 -800 475190 400
rect 476274 -800 476386 400
rect 477470 -800 477582 400
rect 478666 -800 478778 400
rect 479862 -800 479974 400
rect 481058 -800 481170 400
rect 482254 -800 482366 400
rect 483450 -800 483562 400
rect 484554 -800 484666 400
rect 485750 -800 485862 400
rect 486946 -800 487058 400
rect 488142 -800 488254 400
rect 489338 -800 489450 400
rect 490534 -800 490646 400
rect 491730 -800 491842 400
rect 492926 -800 493038 400
rect 494122 -800 494234 400
rect 495318 -800 495430 400
rect 496514 -800 496626 400
rect 497710 -800 497822 400
rect 498906 -800 499018 400
rect 500102 -800 500214 400
rect 501206 -800 501318 400
rect 502402 -800 502514 400
rect 503598 -800 503710 400
rect 504794 -800 504906 400
rect 505990 -800 506102 400
rect 507186 -800 507298 400
rect 508382 -800 508494 400
rect 509578 -800 509690 400
rect 510774 -800 510886 400
rect 511970 -800 512082 400
rect 513166 -800 513278 400
rect 514362 -800 514474 400
rect 515558 -800 515670 400
rect 516754 -800 516866 400
rect 517858 -800 517970 400
rect 519054 -800 519166 400
rect 520250 -800 520362 400
rect 521446 -800 521558 400
rect 522642 -800 522754 400
rect 523838 -800 523950 400
rect 525034 -800 525146 400
rect 526230 -800 526342 400
rect 527426 -800 527538 400
rect 528622 -800 528734 400
rect 529818 -800 529930 400
rect 531014 -800 531126 400
rect 532210 -800 532322 400
rect 533406 -800 533518 400
rect 534510 -800 534622 400
rect 535706 -800 535818 400
rect 536902 -800 537014 400
rect 538098 -800 538210 400
rect 539294 -800 539406 400
rect 540490 -800 540602 400
rect 541686 -800 541798 400
rect 542882 -800 542994 400
rect 544078 -800 544190 400
rect 545274 -800 545386 400
rect 546470 -800 546582 400
rect 547666 -800 547778 400
rect 548862 -800 548974 400
rect 550058 -800 550170 400
rect 551162 -800 551274 400
rect 552358 -800 552470 400
rect 553554 -800 553666 400
rect 554750 -800 554862 400
rect 555946 -800 556058 400
rect 557142 -800 557254 400
rect 558338 -800 558450 400
rect 559534 -800 559646 400
rect 560730 -800 560842 400
rect 561926 -800 562038 400
rect 563122 -800 563234 400
rect 564318 -800 564430 400
rect 565514 -800 565626 400
rect 566710 -800 566822 400
rect 567814 -800 567926 400
rect 569010 -800 569122 400
rect 570206 -800 570318 400
rect 571402 -800 571514 400
rect 572598 -800 572710 400
rect 573794 -800 573906 400
rect 574990 -800 575102 400
rect 576186 -800 576298 400
rect 577382 -800 577494 400
rect 578578 -800 578690 400
rect 579774 -800 579886 400
rect 580970 -800 581082 400
rect 582166 -800 582278 400
rect 583362 -800 583474 400
<< via2 >>
rect 3514 682216 3570 682272
rect 3422 667956 3478 667992
rect 3422 667936 3424 667956
rect 3424 667936 3476 667956
rect 3476 667936 3478 667956
rect 3054 653520 3110 653576
rect 3422 624824 3478 624880
rect 3422 610408 3478 610464
rect 3238 595992 3294 596048
rect 3422 567296 3478 567352
rect 3146 553016 3202 553072
rect 3422 538600 3478 538656
rect 196806 522960 196862 523016
rect 209686 522960 209742 523016
rect 184846 522688 184902 522744
rect 2962 509904 3018 509960
rect 2778 495524 2780 495544
rect 2780 495524 2832 495544
rect 2832 495524 2834 495544
rect 2778 495488 2834 495524
rect 3054 481072 3110 481128
rect 3054 452412 3056 452432
rect 3056 452412 3108 452432
rect 3108 452412 3110 452432
rect 3054 452376 3110 452412
rect 3146 437960 3202 438016
rect 3146 423680 3202 423736
rect 3238 394984 3294 395040
rect 2778 380604 2780 380624
rect 2780 380604 2832 380624
rect 2832 380604 2834 380624
rect 2778 380568 2834 380604
rect 2778 366152 2834 366208
rect 3330 337456 3386 337512
rect 3146 323040 3202 323096
rect 3330 280100 3332 280120
rect 3332 280100 3384 280120
rect 3384 280100 3386 280120
rect 3330 280064 3386 280100
rect 2778 265648 2834 265704
rect 3330 236952 3386 237008
rect 3146 193840 3202 193896
rect 2778 165008 2834 165064
rect 3330 150728 3386 150784
rect 2778 136312 2834 136368
rect 2778 122032 2834 122088
rect 3330 107616 3386 107672
rect 3606 518744 3662 518800
rect 174542 522552 174598 522608
rect 28262 522416 28318 522472
rect 4894 522280 4950 522336
rect 4066 308760 4122 308816
rect 3974 294344 4030 294400
rect 3882 251232 3938 251288
rect 3790 222536 3846 222592
rect 3698 208120 3754 208176
rect 3606 179424 3662 179480
rect 3514 93200 3570 93256
rect 3422 78920 3478 78976
rect 754 64776 810 64832
rect 754 64504 810 64560
rect 2778 50124 2780 50144
rect 2780 50124 2832 50144
rect 2832 50124 2834 50144
rect 2778 50088 2834 50124
rect 6274 517520 6330 517576
rect 12530 517656 12586 517712
rect 12346 517520 12402 517576
rect 10322 217232 10378 217288
rect 2778 35844 2780 35864
rect 2780 35844 2832 35864
rect 2832 35844 2834 35864
rect 2778 35808 2834 35844
rect 478 21936 534 21992
rect 478 21392 534 21448
rect 2962 10240 3018 10296
rect 2962 7112 3018 7168
rect 570 4800 626 4856
rect 5262 3304 5318 3360
rect 22006 517656 22062 517712
rect 22190 517520 22246 517576
rect 27618 517556 27620 517576
rect 27620 517556 27672 517576
rect 27672 517556 27674 517576
rect 27618 517520 27674 517556
rect 21914 6160 21970 6216
rect 181350 522008 181406 522064
rect 177946 521872 178002 521928
rect 176198 521736 176254 521792
rect 190642 522688 190698 522744
rect 190642 522144 190698 522200
rect 191654 520240 191710 520296
rect 201958 522824 202014 522880
rect 222014 522960 222070 523016
rect 209686 522688 209742 522744
rect 252374 700304 252430 700360
rect 267462 645768 267518 645824
rect 267554 640192 267610 640248
rect 267370 578176 267426 578232
rect 267554 578176 267610 578232
rect 269118 578176 269174 578232
rect 269302 578176 269358 578232
rect 267370 568520 267426 568576
rect 267554 568520 267610 568576
rect 269302 540912 269358 540968
rect 269486 540912 269542 540968
rect 267002 531256 267058 531312
rect 267186 531292 267188 531312
rect 267188 531292 267240 531312
rect 267240 531292 267242 531312
rect 267186 531256 267242 531292
rect 276018 550604 276020 550624
rect 276020 550604 276072 550624
rect 276072 550604 276074 550624
rect 276018 550568 276074 550604
rect 276478 550568 276534 550624
rect 287058 550604 287060 550624
rect 287060 550604 287112 550624
rect 287112 550604 287114 550624
rect 287058 550568 287114 550604
rect 287242 550568 287298 550624
rect 287058 549208 287114 549264
rect 287242 549208 287298 549264
rect 291106 549208 291162 549264
rect 291290 549208 291346 549264
rect 293314 531292 293316 531312
rect 293316 531292 293368 531312
rect 293368 531292 293370 531312
rect 293314 531256 293370 531292
rect 293498 531292 293500 531312
rect 293500 531292 293552 531312
rect 293552 531292 293554 531312
rect 293498 531256 293554 531292
rect 543462 700304 543518 700360
rect 579894 697992 579950 698048
rect 494886 686024 494942 686080
rect 494242 685888 494298 685944
rect 580078 686296 580134 686352
rect 580262 674600 580318 674656
rect 579894 651072 579950 651128
rect 580078 639376 580134 639432
rect 580262 627680 580318 627736
rect 299662 540912 299718 540968
rect 299846 540912 299902 540968
rect 579894 604152 579950 604208
rect 580078 592456 580134 592512
rect 493874 579672 493930 579728
rect 494058 579672 494114 579728
rect 580262 580760 580318 580816
rect 494150 560224 494206 560280
rect 494334 560224 494390 560280
rect 579894 557232 579950 557288
rect 580078 545536 580134 545592
rect 494150 540912 494206 540968
rect 494334 540912 494390 540968
rect 580262 533840 580318 533896
rect 311806 522144 311862 522200
rect 311990 522144 312046 522200
rect 370502 522552 370558 522608
rect 353482 522416 353538 522472
rect 325698 522144 325754 522200
rect 335266 522144 335322 522200
rect 345018 522180 345020 522200
rect 345020 522180 345072 522200
rect 345072 522180 345074 522200
rect 345018 522144 345074 522180
rect 356794 522280 356850 522336
rect 354586 522180 354588 522200
rect 354588 522180 354640 522200
rect 354640 522180 354642 522200
rect 354586 522144 354642 522180
rect 37186 517928 37242 517984
rect 57886 517928 57942 517984
rect 77206 517928 77262 517984
rect 96526 517928 96582 517984
rect 115846 517928 115902 517984
rect 135166 517928 135222 517984
rect 154486 517928 154542 517984
rect 166998 517928 167054 517984
rect 50986 517828 50988 517848
rect 50988 517828 51040 517848
rect 51040 517828 51042 517848
rect 50986 517792 51042 517828
rect 70306 517828 70308 517848
rect 70308 517828 70360 517848
rect 70360 517828 70362 517848
rect 70306 517792 70362 517828
rect 89626 517828 89628 517848
rect 89628 517828 89680 517848
rect 89680 517828 89682 517848
rect 89626 517792 89682 517828
rect 108946 517828 108948 517848
rect 108948 517828 109000 517848
rect 109000 517828 109002 517848
rect 108946 517792 109002 517828
rect 128266 517828 128268 517848
rect 128268 517828 128320 517848
rect 128320 517828 128322 517848
rect 128266 517792 128322 517828
rect 147586 517828 147588 517848
rect 147588 517828 147640 517848
rect 147640 517828 147642 517848
rect 147586 517792 147642 517828
rect 166906 517792 166962 517848
rect 52826 7520 52882 7576
rect 172886 519288 172942 519344
rect 193126 519288 193182 519344
rect 195058 519288 195114 519344
rect 198370 519288 198426 519344
rect 199934 519288 199990 519344
rect 205178 519288 205234 519344
rect 210330 519288 210386 519344
rect 225786 519288 225842 519344
rect 315762 519288 315818 519344
rect 341614 519288 341670 519344
rect 359002 519288 359058 519344
rect 361946 519288 362002 519344
rect 363602 519288 363658 519344
rect 370318 518644 370320 518664
rect 370320 518644 370372 518664
rect 370372 518644 370374 518664
rect 370318 518608 370374 518644
rect 170034 4800 170090 4856
rect 172242 217232 172298 217288
rect 171414 154536 171470 154592
rect 171598 154536 171654 154592
rect 171414 135224 171470 135280
rect 171598 135224 171654 135280
rect 171138 3304 171194 3360
rect 173254 212508 173256 212528
rect 173256 212508 173308 212528
rect 173308 212508 173310 212528
rect 173254 212472 173310 212508
rect 173438 212472 173494 212528
rect 173070 154536 173126 154592
rect 173254 154536 173310 154592
rect 173070 135224 173126 135280
rect 173254 135224 173310 135280
rect 178038 63416 178094 63472
rect 178314 63416 178370 63472
rect 176842 6160 176898 6216
rect 184018 191800 184074 191856
rect 184294 191800 184350 191856
rect 187882 7520 187938 7576
rect 189446 116048 189502 116104
rect 189354 115932 189410 115968
rect 189354 115912 189356 115932
rect 189356 115912 189408 115932
rect 189408 115912 189410 115932
rect 191102 154672 191158 154728
rect 191102 154536 191158 154592
rect 191102 106392 191158 106448
rect 191010 106256 191066 106312
rect 191102 65048 191158 65104
rect 191010 64912 191066 64968
rect 191102 54032 191158 54088
rect 191102 53896 191158 53952
rect 190918 53760 190974 53816
rect 191102 53760 191158 53816
rect 194966 154672 195022 154728
rect 194966 154536 195022 154592
rect 194966 143520 195022 143576
rect 194966 142160 195022 142216
rect 194966 66136 195022 66192
rect 194874 57840 194930 57896
rect 195150 37304 195206 37360
rect 194874 37168 194930 37224
rect 200394 154672 200450 154728
rect 200394 154536 200450 154592
rect 200394 135360 200450 135416
rect 200394 135224 200450 135280
rect 200394 96600 200450 96656
rect 200578 96600 200634 96656
rect 201498 39924 201500 39944
rect 201500 39924 201552 39944
rect 201552 39924 201554 39944
rect 201498 39888 201554 39924
rect 201866 154672 201922 154728
rect 201866 154536 201922 154592
rect 201866 135360 201922 135416
rect 201866 135224 201922 135280
rect 201866 96600 201922 96656
rect 202050 96600 202106 96656
rect 201866 40024 201922 40080
rect 203154 87080 203210 87136
rect 203062 86944 203118 87000
rect 212354 212608 212410 212664
rect 211894 212506 211950 212562
rect 212170 212472 212226 212528
rect 212354 212508 212356 212528
rect 212356 212508 212408 212528
rect 212408 212508 212410 212528
rect 212354 212472 212410 212508
rect 211894 58112 211950 58168
rect 211986 57840 212042 57896
rect 212446 40060 212448 40080
rect 212448 40060 212500 40080
rect 212500 40060 212502 40080
rect 212446 40024 212502 40060
rect 216678 202816 216734 202872
rect 216678 183504 216734 183560
rect 217046 211132 217102 211168
rect 217046 211112 217048 211132
rect 217048 211112 217100 211132
rect 217100 211112 217102 211132
rect 217966 211112 218022 211168
rect 216954 202816 217010 202872
rect 216954 183504 217010 183560
rect 219530 93744 219586 93800
rect 219714 193160 219770 193216
rect 219990 193160 220046 193216
rect 219806 133864 219862 133920
rect 219990 133864 220046 133920
rect 219714 93744 219770 93800
rect 220726 40160 220782 40216
rect 224038 133864 224094 133920
rect 224222 133864 224278 133920
rect 225142 200096 225198 200152
rect 225326 200096 225382 200152
rect 225234 180784 225290 180840
rect 225510 180784 225566 180840
rect 225326 140664 225382 140720
rect 225510 140664 225566 140720
rect 229374 212472 229430 212528
rect 229558 212472 229614 212528
rect 228270 139304 228326 139360
rect 228454 139304 228510 139360
rect 229282 182164 229338 182200
rect 229282 182144 229284 182164
rect 229284 182144 229336 182164
rect 229336 182144 229338 182164
rect 229558 182144 229614 182200
rect 229374 125704 229430 125760
rect 229282 125568 229338 125624
rect 229282 86964 229338 87000
rect 229282 86944 229284 86964
rect 229284 86944 229336 86964
rect 229336 86944 229338 86964
rect 229466 86944 229522 87000
rect 230846 190440 230902 190496
rect 231030 190440 231086 190496
rect 230938 154536 230994 154592
rect 231214 154536 231270 154592
rect 231766 143520 231822 143576
rect 232042 212472 232098 212528
rect 232318 212472 232374 212528
rect 232042 193160 232098 193216
rect 232226 193160 232282 193216
rect 232042 143520 232098 143576
rect 235078 183540 235080 183560
rect 235080 183540 235132 183560
rect 235132 183540 235134 183560
rect 235078 183504 235134 183540
rect 235354 183504 235410 183560
rect 235170 164328 235226 164384
rect 235078 164212 235134 164248
rect 235078 164192 235080 164212
rect 235080 164192 235132 164212
rect 235132 164192 235134 164212
rect 234986 137944 235042 138000
rect 235262 137944 235318 138000
rect 235170 125704 235226 125760
rect 235078 125588 235134 125624
rect 235078 125568 235080 125588
rect 235080 125568 235132 125588
rect 235132 125568 235134 125588
rect 235170 106392 235226 106448
rect 235078 106276 235134 106312
rect 235078 106256 235080 106276
rect 235080 106256 235132 106276
rect 235132 106256 235134 106276
rect 235078 86964 235134 87000
rect 235078 86944 235080 86964
rect 235080 86944 235132 86964
rect 235132 86944 235134 86964
rect 235354 86944 235410 87000
rect 234986 41384 235042 41440
rect 235354 41384 235410 41440
rect 236366 48456 236422 48512
rect 236274 48320 236330 48376
rect 258170 77152 258226 77208
rect 258354 77152 258410 77208
rect 261114 172488 261170 172544
rect 261298 172488 261354 172544
rect 260930 67632 260986 67688
rect 261114 67632 261170 67688
rect 262310 154536 262366 154592
rect 262586 154536 262642 154592
rect 262310 135224 262366 135280
rect 262586 135224 262642 135280
rect 262310 115912 262366 115968
rect 262586 115912 262642 115968
rect 262310 96600 262366 96656
rect 262586 96600 262642 96656
rect 266542 191800 266598 191856
rect 266726 191800 266782 191856
rect 268750 29144 268806 29200
rect 268750 29008 268806 29064
rect 270498 40196 270500 40216
rect 270500 40196 270552 40216
rect 270552 40196 270554 40216
rect 270498 40160 270554 40196
rect 272982 172624 273038 172680
rect 273074 172488 273130 172544
rect 275466 219544 275522 219600
rect 275834 219408 275890 219464
rect 275926 217912 275982 217968
rect 275926 217640 275982 217696
rect 275742 40196 275744 40216
rect 275744 40196 275796 40216
rect 275796 40196 275798 40216
rect 275742 40160 275798 40196
rect 276938 201456 276994 201512
rect 277214 201456 277270 201512
rect 277030 162832 277086 162888
rect 277122 153196 277178 153232
rect 277122 153176 277124 153196
rect 277124 153176 277176 153196
rect 277176 153176 277178 153196
rect 277030 143520 277086 143576
rect 277214 143520 277270 143576
rect 277214 3032 277270 3088
rect 282458 211112 282514 211168
rect 282642 211112 282698 211168
rect 282734 183540 282736 183560
rect 282736 183540 282788 183560
rect 282788 183540 282790 183560
rect 282734 183504 282790 183540
rect 282918 183540 282920 183560
rect 282920 183540 282972 183560
rect 282972 183540 282974 183560
rect 282918 183504 282974 183540
rect 282642 164192 282698 164248
rect 282826 164192 282882 164248
rect 280434 3052 280490 3088
rect 280434 3032 280436 3052
rect 280436 3032 280488 3052
rect 280488 3032 280490 3052
rect 283838 201456 283894 201512
rect 284022 201456 284078 201512
rect 283838 182144 283894 182200
rect 284022 182144 284078 182200
rect 283838 162832 283894 162888
rect 284022 162832 284078 162888
rect 284022 106256 284078 106312
rect 285218 191936 285274 191992
rect 285310 191800 285366 191856
rect 284298 124208 284354 124264
rect 286506 202816 286562 202872
rect 286690 202816 286746 202872
rect 286598 183540 286600 183560
rect 286600 183540 286652 183560
rect 286652 183540 286654 183560
rect 286598 183504 286654 183540
rect 286506 183368 286562 183424
rect 286414 106256 286470 106312
rect 286598 106256 286654 106312
rect 284206 3304 284262 3360
rect 289174 212472 289230 212528
rect 289358 212508 289360 212528
rect 289360 212508 289412 212528
rect 289412 212508 289414 212528
rect 289358 212472 289414 212508
rect 289266 202816 289322 202872
rect 289450 202852 289452 202872
rect 289452 202852 289504 202872
rect 289504 202852 289506 202872
rect 289450 202816 289506 202852
rect 289266 193196 289268 193216
rect 289268 193196 289320 193216
rect 289320 193196 289322 193216
rect 289266 193160 289322 193196
rect 289450 193196 289452 193216
rect 289452 193196 289504 193216
rect 289504 193196 289506 193216
rect 289450 193160 289506 193196
rect 289266 183540 289268 183560
rect 289268 183540 289320 183560
rect 289320 183540 289322 183560
rect 289266 183504 289322 183540
rect 289450 183540 289452 183560
rect 289452 183540 289504 183560
rect 289504 183540 289506 183560
rect 289450 183504 289506 183540
rect 289266 153176 289322 153232
rect 289450 153176 289506 153232
rect 289174 106256 289230 106312
rect 289358 106256 289414 106312
rect 289266 17992 289322 18048
rect 289266 17856 289322 17912
rect 289910 40296 289966 40352
rect 289818 40160 289874 40216
rect 291658 193160 291714 193216
rect 291842 193160 291898 193216
rect 291842 134000 291898 134056
rect 291934 133884 291990 133920
rect 291934 133864 291936 133884
rect 291936 133864 291988 133884
rect 291988 133864 291990 133884
rect 291750 124208 291806 124264
rect 291934 124208 291990 124264
rect 297914 4800 297970 4856
rect 298926 86944 298982 87000
rect 299202 86944 299258 87000
rect 306378 4140 306434 4176
rect 306378 4120 306380 4140
rect 306380 4120 306432 4140
rect 306432 4120 306434 4140
rect 311070 4120 311126 4176
rect 317050 173848 317106 173904
rect 317234 173848 317290 173904
rect 316866 67496 316922 67552
rect 317050 67496 317106 67552
rect 316866 57976 316922 58032
rect 317050 57840 317106 57896
rect 318522 147736 318578 147792
rect 318522 143540 318578 143576
rect 318522 143520 318524 143540
rect 318524 143520 318576 143540
rect 318576 143520 318578 143540
rect 318338 96600 318394 96656
rect 318522 96600 318578 96656
rect 318338 67496 318394 67552
rect 318522 67360 318578 67416
rect 318430 46824 318486 46880
rect 318338 46688 318394 46744
rect 328090 173984 328146 174040
rect 328274 173984 328330 174040
rect 327998 164192 328054 164248
rect 328182 164192 328238 164248
rect 327906 48320 327962 48376
rect 328090 48320 328146 48376
rect 329286 164192 329342 164248
rect 329470 164192 329526 164248
rect 329562 147736 329618 147792
rect 329562 144900 329618 144936
rect 329562 144880 329564 144900
rect 329564 144880 329616 144900
rect 329616 144880 329618 144900
rect 329562 128424 329618 128480
rect 329562 125588 329618 125624
rect 329562 125568 329564 125588
rect 329564 125568 329616 125588
rect 329616 125568 329618 125588
rect 329562 109112 329618 109168
rect 329562 106276 329618 106312
rect 329562 106256 329564 106276
rect 329564 106256 329616 106276
rect 329616 106256 329618 106276
rect 329562 51176 329618 51232
rect 329470 48320 329526 48376
rect 331034 8880 331090 8936
rect 331310 217776 331366 217832
rect 331770 217232 331826 217288
rect 333794 6160 333850 6216
rect 332414 3304 332470 3360
rect 338210 40568 338266 40624
rect 338210 40160 338266 40216
rect 340786 217812 340788 217832
rect 340788 217812 340840 217832
rect 340840 217812 340842 217832
rect 340786 217776 340842 217812
rect 341798 201456 341854 201512
rect 341982 201456 342038 201512
rect 341706 62056 341762 62112
rect 341890 62056 341946 62112
rect 343178 193160 343234 193216
rect 343362 193160 343418 193216
rect 342994 182144 343050 182200
rect 343178 182144 343234 182200
rect 343178 172488 343234 172544
rect 343362 172488 343418 172544
rect 343270 160248 343326 160304
rect 343270 160112 343326 160168
rect 343362 65048 343418 65104
rect 343178 64912 343234 64968
rect 344374 193160 344430 193216
rect 344650 193160 344706 193216
rect 344466 172488 344522 172544
rect 344650 172488 344706 172544
rect 345478 162832 345534 162888
rect 345662 162832 345718 162888
rect 345662 132504 345718 132560
rect 345846 132504 345902 132560
rect 352838 212472 352894 212528
rect 353022 212472 353078 212528
rect 354126 201456 354182 201512
rect 354402 201456 354458 201512
rect 354218 193160 354274 193216
rect 354402 193160 354458 193216
rect 355414 201456 355470 201512
rect 355690 201456 355746 201512
rect 355414 193160 355470 193216
rect 355690 193160 355746 193216
rect 355506 144880 355562 144936
rect 355690 144880 355746 144936
rect 360934 172488 360990 172544
rect 361118 172508 361174 172544
rect 361118 172488 361120 172508
rect 361120 172488 361172 172508
rect 361172 172488 361174 172508
rect 361210 106392 361266 106448
rect 361302 106256 361358 106312
rect 362314 122848 362370 122904
rect 362590 122848 362646 122904
rect 362498 9560 362554 9616
rect 363602 9424 363658 9480
rect 367098 40316 367154 40352
rect 367098 40296 367100 40316
rect 367100 40296 367152 40316
rect 367152 40296 367154 40316
rect 369582 7520 369638 7576
rect 369950 40024 370006 40080
rect 372066 518880 372122 518936
rect 371882 518336 371938 518392
rect 375286 518744 375342 518800
rect 371882 518064 371938 518120
rect 372066 518064 372122 518120
rect 371146 517928 371202 517984
rect 371882 486376 371938 486432
rect 371882 485832 371938 485888
rect 580814 522144 580870 522200
rect 580630 522008 580686 522064
rect 580446 521872 580502 521928
rect 580262 521736 580318 521792
rect 379426 518744 379482 518800
rect 379610 518608 379666 518664
rect 386418 518608 386474 518664
rect 399298 518608 399354 518664
rect 405738 518608 405794 518664
rect 418066 518608 418122 518664
rect 425058 518608 425114 518664
rect 437386 518608 437442 518664
rect 444378 518608 444434 518664
rect 456706 518608 456762 518664
rect 463698 518608 463754 518664
rect 476026 518608 476082 518664
rect 483018 518608 483074 518664
rect 495346 518608 495402 518664
rect 502338 518608 502394 518664
rect 514666 518608 514722 518664
rect 553398 518608 553454 518664
rect 562966 518608 563022 518664
rect 580078 518608 580134 518664
rect 579802 518472 579858 518528
rect 579618 518336 579674 518392
rect 405830 517928 405886 517984
rect 418066 517928 418122 517984
rect 425150 517928 425206 517984
rect 437386 517928 437442 517984
rect 444470 517928 444526 517984
rect 456706 517928 456762 517984
rect 463790 517928 463846 517984
rect 476026 517928 476082 517984
rect 483110 517928 483166 517984
rect 495346 517928 495402 517984
rect 502430 517928 502486 517984
rect 514666 517928 514722 517984
rect 553398 517928 553454 517984
rect 562966 517928 563022 517984
rect 386418 517792 386474 517848
rect 399298 517792 399354 517848
rect 576858 486920 576914 486976
rect 394606 486240 394662 486296
rect 379610 485968 379666 486024
rect 405646 486104 405702 486160
rect 398746 486004 398748 486024
rect 398748 486004 398800 486024
rect 398800 486004 398802 486024
rect 398746 485968 398802 486004
rect 379426 485832 379482 485888
rect 394606 485832 394662 485888
rect 576858 485832 576914 485888
rect 576858 299240 576914 299296
rect 576858 298152 576914 298208
rect 579710 518064 579766 518120
rect 579618 275712 579674 275768
rect 579986 510312 580042 510368
rect 579894 498616 579950 498672
rect 579894 463392 579950 463448
rect 579894 451696 579950 451752
rect 579894 439864 579950 439920
rect 579894 416472 579950 416528
rect 579894 404776 579950 404832
rect 579894 392944 579950 393000
rect 579894 369552 579950 369608
rect 579802 263880 579858 263936
rect 576858 252320 576914 252376
rect 576858 251232 576914 251288
rect 580170 518200 580226 518256
rect 580078 357856 580134 357912
rect 580078 346024 580134 346080
rect 580078 322632 580134 322688
rect 579986 228792 580042 228848
rect 379610 40160 379666 40216
rect 379426 40024 379482 40080
rect 372802 4800 372858 4856
rect 394606 40432 394662 40488
rect 398746 40196 398748 40216
rect 398748 40196 398800 40216
rect 398800 40196 398802 40216
rect 398746 40160 398802 40196
rect 394606 40024 394662 40080
rect 405646 40296 405702 40352
rect 466826 8880 466882 8936
rect 470598 217232 470654 217288
rect 476302 6160 476358 6216
rect 580170 216960 580226 217016
rect 576858 205400 576914 205456
rect 576858 204312 576914 204368
rect 580170 170040 580226 170096
rect 580538 134816 580594 134872
rect 580722 158344 580778 158400
rect 583390 486920 583446 486976
rect 583390 486784 583446 486840
rect 583390 310800 583446 310856
rect 583390 310664 583446 310720
rect 583390 299240 583446 299296
rect 583390 299104 583446 299160
rect 583390 252320 583446 252376
rect 583390 252184 583446 252240
rect 583390 205400 583446 205456
rect 583390 205264 583446 205320
rect 580906 181872 580962 181928
rect 580814 123120 580870 123176
rect 580630 111424 580686 111480
rect 580446 87896 580502 87952
rect 580354 76200 580410 76256
rect 580262 64504 580318 64560
rect 576858 41112 576914 41168
rect 583390 41112 583446 41168
rect 583390 40976 583446 41032
rect 576858 40024 576914 40080
rect 580262 29280 580318 29336
rect 579618 17584 579674 17640
rect 580998 7520 581054 7576
<< metal3 >>
rect 252369 700362 252435 700365
rect 543457 700362 543523 700365
rect 252369 700360 543523 700362
rect 252369 700304 252374 700360
rect 252430 700304 543462 700360
rect 543518 700304 543523 700360
rect 252369 700302 543523 700304
rect 252369 700299 252435 700302
rect 543457 700299 543523 700302
rect 579889 698050 579955 698053
rect 583600 698050 584800 698140
rect 579889 698048 584800 698050
rect 579889 697992 579894 698048
rect 579950 697992 584800 698048
rect 579889 697990 584800 697992
rect 579889 697987 579955 697990
rect 583600 697900 584800 697990
rect -800 696540 400 696780
rect 580073 686354 580139 686357
rect 583600 686354 584800 686444
rect 580073 686352 584800 686354
rect 580073 686296 580078 686352
rect 580134 686296 584800 686352
rect 580073 686294 584800 686296
rect 580073 686291 580139 686294
rect 583600 686204 584800 686294
rect 494881 686082 494947 686085
rect 494102 686080 494947 686082
rect 494102 686024 494886 686080
rect 494942 686024 494947 686080
rect 494102 686022 494947 686024
rect 494102 685946 494162 686022
rect 494881 686019 494947 686022
rect 494237 685946 494303 685949
rect 494102 685944 494303 685946
rect 494102 685888 494242 685944
rect 494298 685888 494303 685944
rect 494102 685886 494303 685888
rect 494237 685883 494303 685886
rect -800 682274 400 682364
rect 3509 682274 3575 682277
rect -800 682272 3575 682274
rect -800 682216 3514 682272
rect 3570 682216 3575 682272
rect -800 682214 3575 682216
rect -800 682124 400 682214
rect 3509 682211 3575 682214
rect 580257 674658 580323 674661
rect 583600 674658 584800 674748
rect 580257 674656 584800 674658
rect 580257 674600 580262 674656
rect 580318 674600 584800 674656
rect 580257 674598 584800 674600
rect 580257 674595 580323 674598
rect 583600 674508 584800 674598
rect -800 667994 400 668084
rect 3417 667994 3483 667997
rect -800 667992 3483 667994
rect -800 667936 3422 667992
rect 3478 667936 3483 667992
rect -800 667934 3483 667936
rect -800 667844 400 667934
rect 3417 667931 3483 667934
rect 583600 662676 584800 662916
rect -800 653578 400 653668
rect 3049 653578 3115 653581
rect -800 653576 3115 653578
rect -800 653520 3054 653576
rect 3110 653520 3115 653576
rect -800 653518 3115 653520
rect -800 653428 400 653518
rect 3049 653515 3115 653518
rect 579889 651130 579955 651133
rect 583600 651130 584800 651220
rect 579889 651128 584800 651130
rect 579889 651072 579894 651128
rect 579950 651072 584800 651128
rect 579889 651070 584800 651072
rect 579889 651067 579955 651070
rect 583600 650980 584800 651070
rect 267457 645828 267523 645829
rect 267406 645764 267412 645828
rect 267476 645826 267523 645828
rect 267476 645824 267568 645826
rect 267518 645768 267568 645824
rect 267476 645766 267568 645768
rect 267476 645764 267523 645766
rect 267457 645763 267523 645764
rect 267406 640188 267412 640252
rect 267476 640250 267482 640252
rect 267549 640250 267615 640253
rect 267476 640248 267615 640250
rect 267476 640192 267554 640248
rect 267610 640192 267615 640248
rect 267476 640190 267615 640192
rect 267476 640188 267482 640190
rect 267549 640187 267615 640190
rect 580073 639434 580139 639437
rect 583600 639434 584800 639524
rect 580073 639432 584800 639434
rect 580073 639376 580078 639432
rect 580134 639376 584800 639432
rect 580073 639374 584800 639376
rect 580073 639371 580139 639374
rect 583600 639284 584800 639374
rect -800 639012 400 639252
rect 580257 627738 580323 627741
rect 583600 627738 584800 627828
rect 580257 627736 584800 627738
rect 580257 627680 580262 627736
rect 580318 627680 584800 627736
rect 580257 627678 584800 627680
rect 580257 627675 580323 627678
rect 583600 627588 584800 627678
rect -800 624882 400 624972
rect 3417 624882 3483 624885
rect -800 624880 3483 624882
rect -800 624824 3422 624880
rect 3478 624824 3483 624880
rect -800 624822 3483 624824
rect -800 624732 400 624822
rect 3417 624819 3483 624822
rect 583600 615756 584800 615996
rect -800 610466 400 610556
rect 3417 610466 3483 610469
rect -800 610464 3483 610466
rect -800 610408 3422 610464
rect 3478 610408 3483 610464
rect -800 610406 3483 610408
rect -800 610316 400 610406
rect 3417 610403 3483 610406
rect 579889 604210 579955 604213
rect 583600 604210 584800 604300
rect 579889 604208 584800 604210
rect 579889 604152 579894 604208
rect 579950 604152 584800 604208
rect 579889 604150 584800 604152
rect 579889 604147 579955 604150
rect 583600 604060 584800 604150
rect -800 596050 400 596140
rect 3233 596050 3299 596053
rect -800 596048 3299 596050
rect -800 595992 3238 596048
rect 3294 595992 3299 596048
rect -800 595990 3299 595992
rect -800 595900 400 595990
rect 3233 595987 3299 595990
rect 580073 592514 580139 592517
rect 583600 592514 584800 592604
rect 580073 592512 584800 592514
rect 580073 592456 580078 592512
rect 580134 592456 584800 592512
rect 580073 592454 584800 592456
rect 580073 592451 580139 592454
rect 583600 592364 584800 592454
rect -800 581620 400 581860
rect 580257 580818 580323 580821
rect 583600 580818 584800 580908
rect 580257 580816 584800 580818
rect 580257 580760 580262 580816
rect 580318 580760 584800 580816
rect 580257 580758 584800 580760
rect 580257 580755 580323 580758
rect 583600 580668 584800 580758
rect 493869 579730 493935 579733
rect 494053 579730 494119 579733
rect 493869 579728 494119 579730
rect 493869 579672 493874 579728
rect 493930 579672 494058 579728
rect 494114 579672 494119 579728
rect 493869 579670 494119 579672
rect 493869 579667 493935 579670
rect 494053 579667 494119 579670
rect 267365 578234 267431 578237
rect 267549 578234 267615 578237
rect 267365 578232 267615 578234
rect 267365 578176 267370 578232
rect 267426 578176 267554 578232
rect 267610 578176 267615 578232
rect 267365 578174 267615 578176
rect 267365 578171 267431 578174
rect 267549 578171 267615 578174
rect 269113 578234 269179 578237
rect 269297 578234 269363 578237
rect 269113 578232 269363 578234
rect 269113 578176 269118 578232
rect 269174 578176 269302 578232
rect 269358 578176 269363 578232
rect 269113 578174 269363 578176
rect 269113 578171 269179 578174
rect 269297 578171 269363 578174
rect 583600 568836 584800 569076
rect 267365 568578 267431 568581
rect 267549 568578 267615 568581
rect 267365 568576 267615 568578
rect 267365 568520 267370 568576
rect 267426 568520 267554 568576
rect 267610 568520 267615 568576
rect 267365 568518 267615 568520
rect 267365 568515 267431 568518
rect 267549 568515 267615 568518
rect -800 567354 400 567444
rect 3417 567354 3483 567357
rect -800 567352 3483 567354
rect -800 567296 3422 567352
rect 3478 567296 3483 567352
rect -800 567294 3483 567296
rect -800 567204 400 567294
rect 3417 567291 3483 567294
rect 494145 560282 494211 560285
rect 494329 560282 494395 560285
rect 494145 560280 494395 560282
rect 494145 560224 494150 560280
rect 494206 560224 494334 560280
rect 494390 560224 494395 560280
rect 494145 560222 494395 560224
rect 494145 560219 494211 560222
rect 494329 560219 494395 560222
rect 579889 557290 579955 557293
rect 583600 557290 584800 557380
rect 579889 557288 584800 557290
rect 579889 557232 579894 557288
rect 579950 557232 584800 557288
rect 579889 557230 584800 557232
rect 579889 557227 579955 557230
rect 583600 557140 584800 557230
rect -800 553074 400 553164
rect 3141 553074 3207 553077
rect -800 553072 3207 553074
rect -800 553016 3146 553072
rect 3202 553016 3207 553072
rect -800 553014 3207 553016
rect -800 552924 400 553014
rect 3141 553011 3207 553014
rect 276013 550626 276079 550629
rect 276473 550626 276539 550629
rect 276013 550624 276539 550626
rect 276013 550568 276018 550624
rect 276074 550568 276478 550624
rect 276534 550568 276539 550624
rect 276013 550566 276539 550568
rect 276013 550563 276079 550566
rect 276473 550563 276539 550566
rect 287053 550626 287119 550629
rect 287237 550626 287303 550629
rect 287053 550624 287303 550626
rect 287053 550568 287058 550624
rect 287114 550568 287242 550624
rect 287298 550568 287303 550624
rect 287053 550566 287303 550568
rect 287053 550563 287119 550566
rect 287237 550563 287303 550566
rect 287053 549266 287119 549269
rect 287237 549266 287303 549269
rect 287053 549264 287303 549266
rect 287053 549208 287058 549264
rect 287114 549208 287242 549264
rect 287298 549208 287303 549264
rect 287053 549206 287303 549208
rect 287053 549203 287119 549206
rect 287237 549203 287303 549206
rect 291101 549266 291167 549269
rect 291285 549266 291351 549269
rect 291101 549264 291351 549266
rect 291101 549208 291106 549264
rect 291162 549208 291290 549264
rect 291346 549208 291351 549264
rect 291101 549206 291351 549208
rect 291101 549203 291167 549206
rect 291285 549203 291351 549206
rect 580073 545594 580139 545597
rect 583600 545594 584800 545684
rect 580073 545592 584800 545594
rect 580073 545536 580078 545592
rect 580134 545536 584800 545592
rect 580073 545534 584800 545536
rect 580073 545531 580139 545534
rect 583600 545444 584800 545534
rect 269297 540970 269363 540973
rect 269481 540970 269547 540973
rect 269297 540968 269547 540970
rect 269297 540912 269302 540968
rect 269358 540912 269486 540968
rect 269542 540912 269547 540968
rect 269297 540910 269547 540912
rect 269297 540907 269363 540910
rect 269481 540907 269547 540910
rect 299657 540970 299723 540973
rect 299841 540970 299907 540973
rect 299657 540968 299907 540970
rect 299657 540912 299662 540968
rect 299718 540912 299846 540968
rect 299902 540912 299907 540968
rect 299657 540910 299907 540912
rect 299657 540907 299723 540910
rect 299841 540907 299907 540910
rect 494145 540970 494211 540973
rect 494329 540970 494395 540973
rect 494145 540968 494395 540970
rect 494145 540912 494150 540968
rect 494206 540912 494334 540968
rect 494390 540912 494395 540968
rect 494145 540910 494395 540912
rect 494145 540907 494211 540910
rect 494329 540907 494395 540910
rect -800 538658 400 538748
rect 3417 538658 3483 538661
rect -800 538656 3483 538658
rect -800 538600 3422 538656
rect 3478 538600 3483 538656
rect -800 538598 3483 538600
rect -800 538508 400 538598
rect 3417 538595 3483 538598
rect 580257 533898 580323 533901
rect 583600 533898 584800 533988
rect 580257 533896 584800 533898
rect 580257 533840 580262 533896
rect 580318 533840 584800 533896
rect 580257 533838 584800 533840
rect 580257 533835 580323 533838
rect 583600 533748 584800 533838
rect 266997 531314 267063 531317
rect 267181 531314 267247 531317
rect 266997 531312 267247 531314
rect 266997 531256 267002 531312
rect 267058 531256 267186 531312
rect 267242 531256 267247 531312
rect 266997 531254 267247 531256
rect 266997 531251 267063 531254
rect 267181 531251 267247 531254
rect 293309 531314 293375 531317
rect 293493 531314 293559 531317
rect 293309 531312 293559 531314
rect 293309 531256 293314 531312
rect 293370 531256 293498 531312
rect 293554 531256 293559 531312
rect 293309 531254 293559 531256
rect 293309 531251 293375 531254
rect 293493 531251 293559 531254
rect -800 524092 400 524332
rect 196801 523018 196867 523021
rect 209681 523018 209747 523021
rect 196801 523016 209747 523018
rect 196801 522960 196806 523016
rect 196862 522960 209686 523016
rect 209742 522960 209747 523016
rect 196801 522958 209747 522960
rect 196801 522955 196867 522958
rect 209681 522955 209747 522958
rect 222009 523018 222075 523021
rect 359774 523018 359780 523020
rect 222009 523016 359780 523018
rect 222009 522960 222014 523016
rect 222070 522960 359780 523016
rect 222009 522958 359780 522960
rect 222009 522955 222075 522958
rect 359774 522956 359780 522958
rect 359844 522956 359850 523020
rect 201953 522882 202019 522885
rect 359590 522882 359596 522884
rect 201953 522880 359596 522882
rect 201953 522824 201958 522880
rect 202014 522824 359596 522880
rect 201953 522822 359596 522824
rect 201953 522819 202019 522822
rect 359590 522820 359596 522822
rect 359660 522820 359666 522884
rect 184841 522746 184907 522749
rect 190637 522746 190703 522749
rect 184841 522744 190703 522746
rect 184841 522688 184846 522744
rect 184902 522688 190642 522744
rect 190698 522688 190703 522744
rect 184841 522686 190703 522688
rect 184841 522683 184907 522686
rect 190637 522683 190703 522686
rect 209681 522746 209747 522749
rect 359406 522746 359412 522748
rect 209681 522744 359412 522746
rect 209681 522688 209686 522744
rect 209742 522688 359412 522744
rect 209681 522686 359412 522688
rect 209681 522683 209747 522686
rect 359406 522684 359412 522686
rect 359476 522684 359482 522748
rect 174537 522610 174603 522613
rect 370497 522610 370563 522613
rect 174537 522608 370563 522610
rect 174537 522552 174542 522608
rect 174598 522552 370502 522608
rect 370558 522552 370563 522608
rect 174537 522550 370563 522552
rect 174537 522547 174603 522550
rect 370497 522547 370563 522550
rect 28257 522474 28323 522477
rect 353477 522474 353543 522477
rect 28257 522472 353543 522474
rect 28257 522416 28262 522472
rect 28318 522416 353482 522472
rect 353538 522416 353543 522472
rect 28257 522414 353543 522416
rect 28257 522411 28323 522414
rect 353477 522411 353543 522414
rect 4889 522338 4955 522341
rect 356789 522338 356855 522341
rect 4889 522336 356855 522338
rect 4889 522280 4894 522336
rect 4950 522280 356794 522336
rect 356850 522280 356855 522336
rect 4889 522278 356855 522280
rect 4889 522275 4955 522278
rect 356789 522275 356855 522278
rect 190637 522202 190703 522205
rect 311801 522202 311867 522205
rect 190637 522200 311867 522202
rect 190637 522144 190642 522200
rect 190698 522144 311806 522200
rect 311862 522144 311867 522200
rect 190637 522142 311867 522144
rect 190637 522139 190703 522142
rect 311801 522139 311867 522142
rect 311985 522202 312051 522205
rect 325693 522202 325759 522205
rect 311985 522200 325759 522202
rect 311985 522144 311990 522200
rect 312046 522144 325698 522200
rect 325754 522144 325759 522200
rect 311985 522142 325759 522144
rect 311985 522139 312051 522142
rect 325693 522139 325759 522142
rect 335261 522202 335327 522205
rect 345013 522202 345079 522205
rect 335261 522200 345079 522202
rect 335261 522144 335266 522200
rect 335322 522144 345018 522200
rect 345074 522144 345079 522200
rect 335261 522142 345079 522144
rect 335261 522139 335327 522142
rect 345013 522139 345079 522142
rect 354581 522202 354647 522205
rect 580809 522202 580875 522205
rect 354581 522200 580875 522202
rect 354581 522144 354586 522200
rect 354642 522144 580814 522200
rect 580870 522144 580875 522200
rect 354581 522142 580875 522144
rect 354581 522139 354647 522142
rect 580809 522139 580875 522142
rect 181345 522066 181411 522069
rect 580625 522066 580691 522069
rect 181345 522064 580691 522066
rect 181345 522008 181350 522064
rect 181406 522008 580630 522064
rect 580686 522008 580691 522064
rect 181345 522006 580691 522008
rect 181345 522003 181411 522006
rect 580625 522003 580691 522006
rect 177941 521930 178007 521933
rect 580441 521930 580507 521933
rect 177941 521928 580507 521930
rect 177941 521872 177946 521928
rect 178002 521872 580446 521928
rect 580502 521872 580507 521928
rect 583600 521916 584800 522156
rect 177941 521870 580507 521872
rect 177941 521867 178007 521870
rect 580441 521867 580507 521870
rect 176193 521794 176259 521797
rect 580257 521794 580323 521797
rect 176193 521792 580323 521794
rect 176193 521736 176198 521792
rect 176254 521736 580262 521792
rect 580318 521736 580323 521792
rect 176193 521734 580323 521736
rect 176193 521731 176259 521734
rect 580257 521731 580323 521734
rect 191649 520298 191715 520301
rect 366214 520298 366220 520300
rect 191649 520296 366220 520298
rect 191649 520240 191654 520296
rect 191710 520240 366220 520296
rect 191649 520238 366220 520240
rect 191649 520235 191715 520238
rect 366214 520236 366220 520238
rect 366284 520236 366290 520300
rect 309358 519420 309364 519484
rect 309428 519482 309434 519484
rect 313222 519482 313228 519484
rect 309428 519422 313228 519482
rect 309428 519420 309434 519422
rect 313222 519420 313228 519422
rect 313292 519420 313298 519484
rect 172881 519346 172947 519349
rect 193121 519348 193187 519349
rect 173382 519346 173388 519348
rect 172881 519344 173388 519346
rect 172881 519288 172886 519344
rect 172942 519288 173388 519344
rect 172881 519286 173388 519288
rect 172881 519283 172947 519286
rect 173382 519284 173388 519286
rect 173452 519284 173458 519348
rect 193070 519346 193076 519348
rect 193030 519286 193076 519346
rect 193140 519344 193187 519348
rect 193182 519288 193187 519344
rect 193070 519284 193076 519286
rect 193140 519284 193187 519288
rect 193121 519283 193187 519284
rect 195053 519348 195119 519349
rect 198365 519348 198431 519349
rect 199929 519348 199995 519349
rect 195053 519344 195100 519348
rect 195164 519346 195170 519348
rect 195053 519288 195058 519344
rect 195053 519284 195100 519288
rect 195164 519286 195210 519346
rect 198365 519344 198412 519348
rect 198476 519346 198482 519348
rect 199878 519346 199884 519348
rect 198365 519288 198370 519344
rect 195164 519284 195170 519286
rect 198365 519284 198412 519288
rect 198476 519286 198522 519346
rect 199838 519286 199884 519346
rect 199948 519344 199995 519348
rect 199990 519288 199995 519344
rect 198476 519284 198482 519286
rect 199878 519284 199884 519286
rect 199948 519284 199995 519288
rect 195053 519283 195119 519284
rect 198365 519283 198431 519284
rect 199929 519283 199995 519284
rect 205173 519348 205239 519349
rect 210325 519348 210391 519349
rect 205173 519344 205220 519348
rect 205284 519346 205290 519348
rect 205173 519288 205178 519344
rect 205173 519284 205220 519288
rect 205284 519286 205330 519346
rect 210325 519344 210372 519348
rect 210436 519346 210442 519348
rect 225781 519346 225847 519349
rect 210325 519288 210330 519344
rect 205284 519284 205290 519286
rect 210325 519284 210372 519288
rect 210436 519286 210482 519346
rect 225781 519344 225890 519346
rect 225781 519288 225786 519344
rect 225842 519288 225890 519344
rect 210436 519284 210442 519286
rect 205173 519283 205239 519284
rect 210325 519283 210391 519284
rect 225781 519283 225890 519288
rect 234286 519284 234292 519348
rect 234356 519346 234362 519348
rect 236494 519346 236500 519348
rect 234356 519286 236500 519346
rect 234356 519284 234362 519286
rect 236494 519284 236500 519286
rect 236564 519284 236570 519348
rect 280102 519284 280108 519348
rect 280172 519346 280178 519348
rect 284886 519346 284892 519348
rect 280172 519286 284892 519346
rect 280172 519284 280178 519286
rect 284886 519284 284892 519286
rect 284956 519284 284962 519348
rect 312670 519284 312676 519348
rect 312740 519346 312746 519348
rect 315757 519346 315823 519349
rect 341609 519346 341675 519349
rect 312740 519344 315823 519346
rect 312740 519288 315762 519344
rect 315818 519288 315823 519344
rect 312740 519286 315823 519288
rect 312740 519284 312746 519286
rect 315757 519283 315823 519286
rect 341566 519344 341675 519346
rect 341566 519288 341614 519344
rect 341670 519288 341675 519344
rect 341566 519283 341675 519288
rect 358997 519348 359063 519349
rect 358997 519344 359044 519348
rect 359108 519346 359114 519348
rect 358997 519288 359002 519344
rect 358997 519284 359044 519288
rect 359108 519286 359154 519346
rect 359108 519284 359114 519286
rect 361614 519284 361620 519348
rect 361684 519346 361690 519348
rect 361941 519346 362007 519349
rect 361684 519344 362007 519346
rect 361684 519288 361946 519344
rect 362002 519288 362007 519344
rect 361684 519286 362007 519288
rect 361684 519284 361690 519286
rect 358997 519283 359063 519284
rect 361941 519283 362007 519286
rect 362902 519284 362908 519348
rect 362972 519346 362978 519348
rect 363597 519346 363663 519349
rect 362972 519344 363663 519346
rect 362972 519288 363602 519344
rect 363658 519288 363663 519344
rect 362972 519286 363663 519288
rect 362972 519284 362978 519286
rect 363597 519283 363663 519286
rect 225830 519074 225890 519283
rect 234470 519148 234476 519212
rect 234540 519210 234546 519212
rect 236678 519210 236684 519212
rect 234540 519150 236684 519210
rect 234540 519148 234546 519150
rect 236678 519148 236684 519150
rect 236748 519148 236754 519212
rect 241462 519148 241468 519212
rect 241532 519210 241538 519212
rect 246430 519210 246436 519212
rect 241532 519150 246436 519210
rect 241532 519148 241538 519150
rect 246430 519148 246436 519150
rect 246500 519148 246506 519212
rect 263174 519148 263180 519212
rect 263244 519210 263250 519212
rect 265566 519210 265572 519212
rect 263244 519150 265572 519210
rect 263244 519148 263250 519150
rect 265566 519148 265572 519150
rect 265636 519148 265642 519212
rect 294454 519148 294460 519212
rect 294524 519210 294530 519212
rect 299238 519210 299244 519212
rect 294524 519150 299244 519210
rect 294524 519148 294530 519150
rect 299238 519148 299244 519150
rect 299308 519148 299314 519212
rect 313222 519148 313228 519212
rect 313292 519210 313298 519212
rect 322790 519210 322796 519212
rect 313292 519150 322796 519210
rect 313292 519148 313298 519150
rect 322790 519148 322796 519150
rect 322860 519148 322866 519212
rect 236862 519074 236868 519076
rect 225830 519014 236868 519074
rect 236862 519012 236868 519014
rect 236932 519012 236938 519076
rect 263358 519012 263364 519076
rect 263428 519074 263434 519076
rect 263428 519014 265082 519074
rect 263428 519012 263434 519014
rect 243494 518878 244474 518938
rect 3601 518802 3667 518805
rect 241462 518802 241468 518804
rect 3601 518800 241468 518802
rect 3601 518744 3606 518800
rect 3662 518744 241468 518800
rect 3601 518742 241468 518744
rect 3601 518739 3667 518742
rect 241462 518740 241468 518742
rect 241532 518740 241538 518804
rect 210366 518604 210372 518668
rect 210436 518666 210442 518668
rect 234470 518666 234476 518668
rect 210436 518606 234476 518666
rect 210436 518604 210442 518606
rect 234470 518604 234476 518606
rect 234540 518604 234546 518668
rect 234846 518606 235274 518666
rect 182214 518468 182220 518532
rect 182284 518530 182290 518532
rect 182284 518470 191666 518530
rect 182284 518468 182290 518470
rect 37181 517986 37247 517989
rect 57881 517986 57947 517989
rect 77201 517986 77267 517989
rect 96521 517986 96587 517989
rect 115841 517986 115907 517989
rect 135161 517986 135227 517989
rect 154481 517986 154547 517989
rect 166993 517986 167059 517989
rect 176510 517986 176516 517988
rect 37181 517984 41522 517986
rect 37181 517928 37186 517984
rect 37242 517928 41522 517984
rect 37181 517926 41522 517928
rect 37181 517923 37247 517926
rect 41462 517850 41522 517926
rect 57881 517984 60842 517986
rect 57881 517928 57886 517984
rect 57942 517928 60842 517984
rect 57881 517926 60842 517928
rect 57881 517923 57947 517926
rect 50981 517850 51047 517853
rect 41462 517848 51047 517850
rect 41462 517792 50986 517848
rect 51042 517792 51047 517848
rect 41462 517790 51047 517792
rect 60782 517850 60842 517926
rect 77201 517984 80162 517986
rect 77201 517928 77206 517984
rect 77262 517928 80162 517984
rect 77201 517926 80162 517928
rect 77201 517923 77267 517926
rect 70301 517850 70367 517853
rect 60782 517848 70367 517850
rect 60782 517792 70306 517848
rect 70362 517792 70367 517848
rect 60782 517790 70367 517792
rect 80102 517850 80162 517926
rect 96521 517984 99482 517986
rect 96521 517928 96526 517984
rect 96582 517928 99482 517984
rect 96521 517926 99482 517928
rect 96521 517923 96587 517926
rect 89621 517850 89687 517853
rect 80102 517848 89687 517850
rect 80102 517792 89626 517848
rect 89682 517792 89687 517848
rect 80102 517790 89687 517792
rect 99422 517850 99482 517926
rect 115841 517984 118802 517986
rect 115841 517928 115846 517984
rect 115902 517928 118802 517984
rect 115841 517926 118802 517928
rect 115841 517923 115907 517926
rect 108941 517850 109007 517853
rect 99422 517848 109007 517850
rect 99422 517792 108946 517848
rect 109002 517792 109007 517848
rect 99422 517790 109007 517792
rect 118742 517850 118802 517926
rect 135161 517984 138122 517986
rect 135161 517928 135166 517984
rect 135222 517928 138122 517984
rect 135161 517926 138122 517928
rect 135161 517923 135227 517926
rect 128261 517850 128327 517853
rect 118742 517848 128327 517850
rect 118742 517792 128266 517848
rect 128322 517792 128327 517848
rect 118742 517790 128327 517792
rect 138062 517850 138122 517926
rect 154481 517984 157442 517986
rect 154481 517928 154486 517984
rect 154542 517928 157442 517984
rect 154481 517926 157442 517928
rect 154481 517923 154547 517926
rect 147581 517850 147647 517853
rect 138062 517848 147647 517850
rect 138062 517792 147586 517848
rect 147642 517792 147647 517848
rect 138062 517790 147647 517792
rect 157382 517850 157442 517926
rect 166993 517984 176516 517986
rect 166993 517928 166998 517984
rect 167054 517928 176516 517984
rect 166993 517926 176516 517928
rect 166993 517923 167059 517926
rect 176510 517924 176516 517926
rect 176580 517924 176586 517988
rect 176694 517924 176700 517988
rect 176764 517986 176770 517988
rect 176764 517926 182098 517986
rect 176764 517924 176770 517926
rect 166901 517850 166967 517853
rect 157382 517848 166967 517850
rect 157382 517792 166906 517848
rect 166962 517792 166967 517848
rect 157382 517790 166967 517792
rect 182038 517850 182098 517926
rect 182214 517924 182220 517988
rect 182284 517924 182290 517988
rect 182222 517850 182282 517924
rect 182038 517790 182282 517850
rect 191606 517850 191666 518470
rect 199878 518468 199884 518532
rect 199948 518530 199954 518532
rect 234846 518530 234906 518606
rect 199948 518470 234906 518530
rect 235214 518530 235274 518606
rect 236862 518604 236868 518668
rect 236932 518666 236938 518668
rect 243494 518666 243554 518878
rect 236932 518606 243554 518666
rect 236932 518604 236938 518606
rect 243854 518604 243860 518668
rect 243924 518666 243930 518668
rect 244222 518666 244228 518668
rect 243924 518606 244228 518666
rect 243924 518604 243930 518606
rect 244222 518604 244228 518606
rect 244292 518604 244298 518668
rect 244414 518666 244474 518878
rect 253606 518876 253612 518940
rect 253676 518938 253682 518940
rect 253676 518878 264898 518938
rect 253676 518876 253682 518878
rect 246430 518740 246436 518804
rect 246500 518802 246506 518804
rect 263358 518802 263364 518804
rect 246500 518742 263364 518802
rect 246500 518740 246506 518742
rect 263358 518740 263364 518742
rect 263428 518740 263434 518804
rect 253606 518666 253612 518668
rect 244414 518606 253612 518666
rect 253606 518604 253612 518606
rect 253676 518604 253682 518668
rect 253790 518604 253796 518668
rect 253860 518666 253866 518668
rect 263174 518666 263180 518668
rect 253860 518606 263180 518666
rect 253860 518604 253866 518606
rect 263174 518604 263180 518606
rect 263244 518604 263250 518668
rect 264838 518666 264898 518878
rect 265022 518802 265082 519014
rect 272926 519012 272932 519076
rect 272996 519074 273002 519076
rect 280102 519074 280108 519076
rect 272996 519014 280108 519074
rect 272996 519012 273002 519014
rect 280102 519012 280108 519014
rect 280172 519012 280178 519076
rect 294270 518876 294276 518940
rect 294340 518938 294346 518940
rect 298870 518938 298876 518940
rect 294340 518878 298876 518938
rect 294340 518876 294346 518878
rect 298870 518876 298876 518878
rect 298940 518876 298946 518940
rect 301638 518878 302066 518938
rect 301638 518802 301698 518878
rect 265022 518742 283298 518802
rect 272926 518666 272932 518668
rect 264838 518606 272932 518666
rect 272926 518604 272932 518606
rect 272996 518604 273002 518668
rect 273110 518604 273116 518668
rect 273180 518666 273186 518668
rect 283046 518666 283052 518668
rect 273180 518606 283052 518666
rect 273180 518604 273186 518606
rect 283046 518604 283052 518606
rect 283116 518604 283122 518668
rect 283238 518666 283298 518742
rect 283606 518742 301698 518802
rect 302006 518802 302066 518878
rect 302734 518876 302740 518940
rect 302804 518938 302810 518940
rect 312670 518938 312676 518940
rect 302804 518878 312676 518938
rect 302804 518876 302810 518878
rect 312670 518876 312676 518878
rect 312740 518876 312746 518940
rect 302006 518742 318074 518802
rect 283606 518666 283666 518742
rect 283238 518606 283666 518666
rect 284886 518604 284892 518668
rect 284956 518666 284962 518668
rect 294270 518666 294276 518668
rect 284956 518606 294276 518666
rect 284956 518604 284962 518606
rect 294270 518604 294276 518606
rect 294340 518604 294346 518668
rect 294638 518604 294644 518668
rect 294708 518666 294714 518668
rect 298686 518666 298692 518668
rect 294708 518606 298692 518666
rect 294708 518604 294714 518606
rect 298686 518604 298692 518606
rect 298756 518604 298762 518668
rect 298870 518604 298876 518668
rect 298940 518666 298946 518668
rect 301814 518666 301820 518668
rect 298940 518606 301820 518666
rect 298940 518604 298946 518606
rect 301814 518604 301820 518606
rect 301884 518604 301890 518668
rect 301998 518604 302004 518668
rect 302068 518666 302074 518668
rect 309174 518666 309180 518668
rect 302068 518606 309180 518666
rect 302068 518604 302074 518606
rect 309174 518604 309180 518606
rect 309244 518604 309250 518668
rect 318014 518666 318074 518742
rect 321686 518740 321692 518804
rect 321756 518802 321762 518804
rect 335302 518802 335308 518804
rect 321756 518742 335308 518802
rect 321756 518740 321762 518742
rect 335302 518740 335308 518742
rect 335372 518740 335378 518804
rect 335494 518742 335922 518802
rect 321502 518666 321508 518668
rect 318014 518606 321508 518666
rect 321502 518604 321508 518606
rect 321572 518604 321578 518668
rect 322790 518604 322796 518668
rect 322860 518666 322866 518668
rect 335494 518666 335554 518742
rect 322860 518606 335554 518666
rect 335862 518666 335922 518742
rect 336406 518740 336412 518804
rect 336476 518802 336482 518804
rect 341566 518802 341626 519283
rect 367318 518876 367324 518940
rect 367388 518938 367394 518940
rect 372061 518938 372127 518941
rect 367388 518936 372127 518938
rect 367388 518880 372066 518936
rect 372122 518880 372127 518936
rect 367388 518878 372127 518880
rect 367388 518876 367394 518878
rect 372061 518875 372127 518878
rect 336476 518742 341626 518802
rect 375281 518802 375347 518805
rect 379421 518802 379487 518805
rect 375281 518800 379487 518802
rect 375281 518744 375286 518800
rect 375342 518744 379426 518800
rect 379482 518744 379487 518800
rect 375281 518742 379487 518744
rect 336476 518740 336482 518742
rect 375281 518739 375347 518742
rect 379421 518739 379487 518742
rect 370313 518666 370379 518669
rect 335862 518664 370379 518666
rect 335862 518608 370318 518664
rect 370374 518608 370379 518664
rect 335862 518606 370379 518608
rect 322860 518604 322866 518606
rect 370313 518603 370379 518606
rect 379605 518666 379671 518669
rect 386413 518666 386479 518669
rect 379605 518664 386479 518666
rect 379605 518608 379610 518664
rect 379666 518608 386418 518664
rect 386474 518608 386479 518664
rect 379605 518606 386479 518608
rect 379605 518603 379671 518606
rect 386413 518603 386479 518606
rect 399293 518666 399359 518669
rect 405733 518666 405799 518669
rect 399293 518664 405799 518666
rect 399293 518608 399298 518664
rect 399354 518608 405738 518664
rect 405794 518608 405799 518664
rect 399293 518606 405799 518608
rect 399293 518603 399359 518606
rect 405733 518603 405799 518606
rect 418061 518666 418127 518669
rect 425053 518666 425119 518669
rect 418061 518664 425119 518666
rect 418061 518608 418066 518664
rect 418122 518608 425058 518664
rect 425114 518608 425119 518664
rect 418061 518606 425119 518608
rect 418061 518603 418127 518606
rect 425053 518603 425119 518606
rect 437381 518666 437447 518669
rect 444373 518666 444439 518669
rect 437381 518664 444439 518666
rect 437381 518608 437386 518664
rect 437442 518608 444378 518664
rect 444434 518608 444439 518664
rect 437381 518606 444439 518608
rect 437381 518603 437447 518606
rect 444373 518603 444439 518606
rect 456701 518666 456767 518669
rect 463693 518666 463759 518669
rect 456701 518664 463759 518666
rect 456701 518608 456706 518664
rect 456762 518608 463698 518664
rect 463754 518608 463759 518664
rect 456701 518606 463759 518608
rect 456701 518603 456767 518606
rect 463693 518603 463759 518606
rect 476021 518666 476087 518669
rect 483013 518666 483079 518669
rect 476021 518664 483079 518666
rect 476021 518608 476026 518664
rect 476082 518608 483018 518664
rect 483074 518608 483079 518664
rect 476021 518606 483079 518608
rect 476021 518603 476087 518606
rect 483013 518603 483079 518606
rect 495341 518666 495407 518669
rect 502333 518666 502399 518669
rect 495341 518664 502399 518666
rect 495341 518608 495346 518664
rect 495402 518608 502338 518664
rect 502394 518608 502399 518664
rect 495341 518606 502399 518608
rect 495341 518603 495407 518606
rect 502333 518603 502399 518606
rect 514661 518666 514727 518669
rect 553393 518666 553459 518669
rect 514661 518664 553459 518666
rect 514661 518608 514666 518664
rect 514722 518608 553398 518664
rect 553454 518608 553459 518664
rect 514661 518606 553459 518608
rect 514661 518603 514727 518606
rect 553393 518603 553459 518606
rect 562961 518666 563027 518669
rect 580073 518666 580139 518669
rect 562961 518664 580139 518666
rect 562961 518608 562966 518664
rect 563022 518608 580078 518664
rect 580134 518608 580139 518664
rect 562961 518606 580139 518608
rect 562961 518603 563027 518606
rect 580073 518603 580139 518606
rect 579797 518530 579863 518533
rect 235214 518528 579863 518530
rect 235214 518472 579802 518528
rect 579858 518472 579863 518528
rect 235214 518470 579863 518472
rect 199948 518468 199954 518470
rect 579797 518467 579863 518470
rect 198406 518332 198412 518396
rect 198476 518394 198482 518396
rect 234286 518394 234292 518396
rect 198476 518334 234292 518394
rect 198476 518332 198482 518334
rect 234286 518332 234292 518334
rect 234356 518332 234362 518396
rect 234654 518332 234660 518396
rect 234724 518394 234730 518396
rect 236310 518394 236316 518396
rect 234724 518334 236316 518394
rect 234724 518332 234730 518334
rect 236310 518332 236316 518334
rect 236380 518332 236386 518396
rect 236494 518332 236500 518396
rect 236564 518394 236570 518396
rect 367318 518394 367324 518396
rect 236564 518334 367324 518394
rect 236564 518332 236570 518334
rect 367318 518332 367324 518334
rect 367388 518332 367394 518396
rect 371877 518394 371943 518397
rect 579613 518394 579679 518397
rect 371877 518392 579679 518394
rect 371877 518336 371882 518392
rect 371938 518336 579618 518392
rect 579674 518336 579679 518392
rect 371877 518334 579679 518336
rect 371877 518331 371943 518334
rect 579613 518331 579679 518334
rect 195094 518196 195100 518260
rect 195164 518258 195170 518260
rect 294454 518258 294460 518260
rect 195164 518198 294460 518258
rect 195164 518196 195170 518198
rect 294454 518196 294460 518198
rect 294524 518196 294530 518260
rect 299054 518258 299060 518260
rect 295198 518198 299060 518258
rect 193070 518060 193076 518124
rect 193140 518122 193146 518124
rect 234654 518122 234660 518124
rect 193140 518062 234660 518122
rect 193140 518060 193146 518062
rect 234654 518060 234660 518062
rect 234724 518060 234730 518124
rect 236310 518060 236316 518124
rect 236380 518122 236386 518124
rect 295198 518122 295258 518198
rect 299054 518196 299060 518198
rect 299124 518196 299130 518260
rect 299238 518196 299244 518260
rect 299308 518258 299314 518260
rect 580165 518258 580231 518261
rect 299308 518256 580231 518258
rect 299308 518200 580170 518256
rect 580226 518200 580231 518256
rect 299308 518198 580231 518200
rect 299308 518196 299314 518198
rect 580165 518195 580231 518198
rect 236380 518062 295258 518122
rect 236380 518060 236386 518062
rect 299238 518060 299244 518124
rect 299308 518122 299314 518124
rect 367134 518122 367140 518124
rect 299308 518062 367140 518122
rect 299308 518060 299314 518062
rect 367134 518060 367140 518062
rect 367204 518060 367210 518124
rect 367318 518060 367324 518124
rect 367388 518122 367394 518124
rect 371877 518122 371943 518125
rect 367388 518120 371943 518122
rect 367388 518064 371882 518120
rect 371938 518064 371943 518120
rect 367388 518062 371943 518064
rect 367388 518060 367394 518062
rect 371877 518059 371943 518062
rect 372061 518122 372127 518125
rect 579705 518122 579771 518125
rect 372061 518120 579771 518122
rect 372061 518064 372066 518120
rect 372122 518064 579710 518120
rect 579766 518064 579771 518120
rect 372061 518062 579771 518064
rect 372061 518059 372127 518062
rect 579705 518059 579771 518062
rect 196014 517924 196020 517988
rect 196084 517986 196090 517988
rect 210366 517986 210372 517988
rect 196084 517926 210372 517986
rect 196084 517924 196090 517926
rect 210366 517924 210372 517926
rect 210436 517924 210442 517988
rect 219198 517924 219204 517988
rect 219268 517986 219274 517988
rect 234470 517986 234476 517988
rect 219268 517926 234476 517986
rect 219268 517924 219274 517926
rect 234470 517924 234476 517926
rect 234540 517924 234546 517988
rect 236678 517924 236684 517988
rect 236748 517986 236754 517988
rect 243302 517986 243308 517988
rect 236748 517926 243308 517986
rect 236748 517924 236754 517926
rect 243302 517924 243308 517926
rect 243372 517924 243378 517988
rect 243670 517924 243676 517988
rect 243740 517986 243746 517988
rect 244222 517986 244228 517988
rect 243740 517926 244228 517986
rect 243740 517924 243746 517926
rect 244222 517924 244228 517926
rect 244292 517924 244298 517988
rect 244406 517924 244412 517988
rect 244476 517986 244482 517988
rect 253790 517986 253796 517988
rect 244476 517926 253796 517986
rect 244476 517924 244482 517926
rect 253790 517924 253796 517926
rect 253860 517924 253866 517988
rect 254158 517924 254164 517988
rect 254228 517986 254234 517988
rect 264462 517986 264468 517988
rect 254228 517926 264468 517986
rect 254228 517924 254234 517926
rect 264462 517924 264468 517926
rect 264532 517924 264538 517988
rect 265566 517924 265572 517988
rect 265636 517986 265642 517988
rect 273110 517986 273116 517988
rect 265636 517926 273116 517986
rect 265636 517924 265642 517926
rect 273110 517924 273116 517926
rect 273180 517924 273186 517988
rect 273478 517924 273484 517988
rect 273548 517986 273554 517988
rect 282862 517986 282868 517988
rect 273548 517926 282868 517986
rect 273548 517924 273554 517926
rect 282862 517924 282868 517926
rect 282932 517924 282938 517988
rect 283046 517924 283052 517988
rect 283116 517986 283122 517988
rect 294638 517986 294644 517988
rect 283116 517926 294644 517986
rect 283116 517924 283122 517926
rect 294638 517924 294644 517926
rect 294708 517924 294714 517988
rect 298870 517924 298876 517988
rect 298940 517986 298946 517988
rect 301998 517986 302004 517988
rect 298940 517926 302004 517986
rect 298940 517924 298946 517926
rect 301998 517924 302004 517926
rect 302068 517924 302074 517988
rect 302182 517924 302188 517988
rect 302252 517986 302258 517988
rect 371141 517986 371207 517989
rect 302252 517984 371207 517986
rect 302252 517928 371146 517984
rect 371202 517928 371207 517984
rect 302252 517926 371207 517928
rect 302252 517924 302258 517926
rect 371141 517923 371207 517926
rect 405825 517986 405891 517989
rect 418061 517986 418127 517989
rect 405825 517984 418127 517986
rect 405825 517928 405830 517984
rect 405886 517928 418066 517984
rect 418122 517928 418127 517984
rect 405825 517926 418127 517928
rect 405825 517923 405891 517926
rect 418061 517923 418127 517926
rect 425145 517986 425211 517989
rect 437381 517986 437447 517989
rect 425145 517984 437447 517986
rect 425145 517928 425150 517984
rect 425206 517928 437386 517984
rect 437442 517928 437447 517984
rect 425145 517926 437447 517928
rect 425145 517923 425211 517926
rect 437381 517923 437447 517926
rect 444465 517986 444531 517989
rect 456701 517986 456767 517989
rect 444465 517984 456767 517986
rect 444465 517928 444470 517984
rect 444526 517928 456706 517984
rect 456762 517928 456767 517984
rect 444465 517926 456767 517928
rect 444465 517923 444531 517926
rect 456701 517923 456767 517926
rect 463785 517986 463851 517989
rect 476021 517986 476087 517989
rect 463785 517984 476087 517986
rect 463785 517928 463790 517984
rect 463846 517928 476026 517984
rect 476082 517928 476087 517984
rect 463785 517926 476087 517928
rect 463785 517923 463851 517926
rect 476021 517923 476087 517926
rect 483105 517986 483171 517989
rect 495341 517986 495407 517989
rect 483105 517984 495407 517986
rect 483105 517928 483110 517984
rect 483166 517928 495346 517984
rect 495402 517928 495407 517984
rect 483105 517926 495407 517928
rect 483105 517923 483171 517926
rect 495341 517923 495407 517926
rect 502425 517986 502491 517989
rect 514661 517986 514727 517989
rect 502425 517984 514727 517986
rect 502425 517928 502430 517984
rect 502486 517928 514666 517984
rect 514722 517928 514727 517984
rect 502425 517926 514727 517928
rect 502425 517923 502491 517926
rect 514661 517923 514727 517926
rect 553393 517986 553459 517989
rect 562961 517986 563027 517989
rect 553393 517984 563027 517986
rect 553393 517928 553398 517984
rect 553454 517928 562966 517984
rect 563022 517928 563027 517984
rect 553393 517926 563027 517928
rect 553393 517923 553459 517926
rect 562961 517923 563027 517926
rect 195830 517850 195836 517852
rect 191606 517790 195836 517850
rect 50981 517787 51047 517790
rect 70301 517787 70367 517790
rect 89621 517787 89687 517790
rect 108941 517787 109007 517790
rect 128261 517787 128327 517790
rect 147581 517787 147647 517790
rect 166901 517787 166967 517790
rect 195830 517788 195836 517790
rect 195900 517788 195906 517852
rect 205214 517788 205220 517852
rect 205284 517850 205290 517852
rect 298502 517850 298508 517852
rect 205284 517790 298508 517850
rect 205284 517788 205290 517790
rect 298502 517788 298508 517790
rect 298572 517788 298578 517852
rect 298870 517788 298876 517852
rect 298940 517850 298946 517852
rect 367318 517850 367324 517852
rect 298940 517790 367324 517850
rect 298940 517788 298946 517790
rect 367318 517788 367324 517790
rect 367388 517788 367394 517852
rect 386413 517850 386479 517853
rect 399293 517850 399359 517853
rect 386413 517848 399359 517850
rect 386413 517792 386418 517848
rect 386474 517792 399298 517848
rect 399354 517792 399359 517848
rect 386413 517790 399359 517792
rect 386413 517787 386479 517790
rect 399293 517787 399359 517790
rect 12525 517714 12591 517717
rect 22001 517714 22067 517717
rect 12525 517712 22067 517714
rect 12525 517656 12530 517712
rect 12586 517656 22006 517712
rect 22062 517656 22067 517712
rect 12525 517654 22067 517656
rect 12525 517651 12591 517654
rect 22001 517651 22067 517654
rect 367318 517652 367324 517716
rect 367388 517714 367394 517716
rect 368974 517714 368980 517716
rect 367388 517654 368980 517714
rect 367388 517652 367394 517654
rect 368974 517652 368980 517654
rect 369044 517652 369050 517716
rect 6269 517578 6335 517581
rect 12341 517578 12407 517581
rect 6269 517576 12407 517578
rect 6269 517520 6274 517576
rect 6330 517520 12346 517576
rect 12402 517520 12407 517576
rect 6269 517518 12407 517520
rect 6269 517515 6335 517518
rect 12341 517515 12407 517518
rect 22185 517578 22251 517581
rect 27613 517578 27679 517581
rect 22185 517576 27679 517578
rect 22185 517520 22190 517576
rect 22246 517520 27618 517576
rect 27674 517520 27679 517576
rect 22185 517518 27679 517520
rect 22185 517515 22251 517518
rect 27613 517515 27679 517518
rect 579981 510370 580047 510373
rect 583600 510370 584800 510460
rect 579981 510368 584800 510370
rect 579981 510312 579986 510368
rect 580042 510312 584800 510368
rect 579981 510310 584800 510312
rect 579981 510307 580047 510310
rect 583600 510220 584800 510310
rect -800 509962 400 510052
rect 2957 509962 3023 509965
rect -800 509960 3023 509962
rect -800 509904 2962 509960
rect 3018 509904 3023 509960
rect -800 509902 3023 509904
rect -800 509812 400 509902
rect 2957 509899 3023 509902
rect 579889 498674 579955 498677
rect 583600 498674 584800 498764
rect 579889 498672 584800 498674
rect 579889 498616 579894 498672
rect 579950 498616 584800 498672
rect 579889 498614 584800 498616
rect 579889 498611 579955 498614
rect 583600 498524 584800 498614
rect -800 495546 400 495636
rect 2773 495546 2839 495549
rect -800 495544 2839 495546
rect -800 495488 2778 495544
rect 2834 495488 2839 495544
rect -800 495486 2839 495488
rect -800 495396 400 495486
rect 2773 495483 2839 495486
rect 576853 486978 576919 486981
rect 583385 486978 583451 486981
rect 576853 486976 583451 486978
rect 576853 486920 576858 486976
rect 576914 486920 583390 486976
rect 583446 486920 583451 486976
rect 576853 486918 583451 486920
rect 576853 486915 576919 486918
rect 583385 486915 583451 486918
rect 583385 486842 583451 486845
rect 583600 486842 584800 486932
rect 583385 486840 584800 486842
rect 583385 486784 583390 486840
rect 583446 486784 584800 486840
rect 583385 486782 584800 486784
rect 583385 486779 583451 486782
rect 583600 486692 584800 486782
rect 367134 486372 367140 486436
rect 367204 486434 367210 486436
rect 371877 486434 371943 486437
rect 367204 486432 371943 486434
rect 367204 486376 371882 486432
rect 371938 486376 371943 486432
rect 367204 486374 371943 486376
rect 367204 486372 367210 486374
rect 371877 486371 371943 486374
rect 384982 486236 384988 486300
rect 385052 486298 385058 486300
rect 394601 486298 394667 486301
rect 385052 486296 394667 486298
rect 385052 486240 394606 486296
rect 394662 486240 394667 486296
rect 385052 486238 394667 486240
rect 385052 486236 385058 486238
rect 394601 486235 394667 486238
rect 367134 486162 367140 486164
rect 360150 486102 367140 486162
rect 359774 485828 359780 485892
rect 359844 485890 359850 485892
rect 360150 485890 360210 486102
rect 367134 486100 367140 486102
rect 367204 486100 367210 486164
rect 405641 486162 405707 486165
rect 405641 486160 412650 486162
rect 405641 486104 405646 486160
rect 405702 486104 412650 486160
rect 405641 486102 412650 486104
rect 405641 486099 405707 486102
rect 379605 486026 379671 486029
rect 384982 486026 384988 486028
rect 379605 486024 384988 486026
rect 379605 485968 379610 486024
rect 379666 485968 384988 486024
rect 379605 485966 384988 485968
rect 379605 485963 379671 485966
rect 384982 485964 384988 485966
rect 385052 485964 385058 486028
rect 398741 486026 398807 486029
rect 396030 486024 398807 486026
rect 396030 485968 398746 486024
rect 398802 485968 398807 486024
rect 396030 485966 398807 485968
rect 412590 486026 412650 486102
rect 422342 486102 431970 486162
rect 412590 485966 422218 486026
rect 359844 485830 360210 485890
rect 371877 485890 371943 485893
rect 379421 485890 379487 485893
rect 371877 485888 379487 485890
rect 371877 485832 371882 485888
rect 371938 485832 379426 485888
rect 379482 485832 379487 485888
rect 371877 485830 379487 485832
rect 359844 485828 359850 485830
rect 371877 485827 371943 485830
rect 379421 485827 379487 485830
rect 394601 485890 394667 485893
rect 396030 485890 396090 485966
rect 398741 485963 398807 485966
rect 394601 485888 396090 485890
rect 394601 485832 394606 485888
rect 394662 485832 396090 485888
rect 394601 485830 396090 485832
rect 422158 485890 422218 485966
rect 422342 485890 422402 486102
rect 431910 486026 431970 486102
rect 441662 486102 451290 486162
rect 431910 485966 441538 486026
rect 422158 485830 422402 485890
rect 441478 485890 441538 485966
rect 441662 485890 441722 486102
rect 451230 486026 451290 486102
rect 460982 486102 470610 486162
rect 451230 485966 460858 486026
rect 441478 485830 441722 485890
rect 460798 485890 460858 485966
rect 460982 485890 461042 486102
rect 470550 486026 470610 486102
rect 480302 486102 489930 486162
rect 470550 485966 480178 486026
rect 460798 485830 461042 485890
rect 480118 485890 480178 485966
rect 480302 485890 480362 486102
rect 489870 486026 489930 486102
rect 499622 486102 509250 486162
rect 489870 485966 499498 486026
rect 480118 485830 480362 485890
rect 499438 485890 499498 485966
rect 499622 485890 499682 486102
rect 509190 486026 509250 486102
rect 518942 486102 528570 486162
rect 509190 485966 518818 486026
rect 499438 485830 499682 485890
rect 518758 485890 518818 485966
rect 518942 485890 519002 486102
rect 528510 486026 528570 486102
rect 538262 486102 547890 486162
rect 528510 485966 538138 486026
rect 518758 485830 519002 485890
rect 538078 485890 538138 485966
rect 538262 485890 538322 486102
rect 547830 486026 547890 486102
rect 557582 486102 567210 486162
rect 547830 485966 557458 486026
rect 538078 485830 538322 485890
rect 557398 485890 557458 485966
rect 557582 485890 557642 486102
rect 567150 486026 567210 486102
rect 567150 485966 576778 486026
rect 557398 485830 557642 485890
rect 576718 485890 576778 485966
rect 576853 485890 576919 485893
rect 576718 485888 576919 485890
rect 576718 485832 576858 485888
rect 576914 485832 576919 485888
rect 576718 485830 576919 485832
rect 394601 485827 394667 485830
rect 576853 485827 576919 485830
rect -800 481130 400 481220
rect 3049 481130 3115 481133
rect -800 481128 3115 481130
rect -800 481072 3054 481128
rect 3110 481072 3115 481128
rect -800 481070 3115 481072
rect -800 480980 400 481070
rect 3049 481067 3115 481070
rect 583600 474996 584800 475236
rect -800 466700 400 466940
rect 579889 463450 579955 463453
rect 583600 463450 584800 463540
rect 579889 463448 584800 463450
rect 579889 463392 579894 463448
rect 579950 463392 584800 463448
rect 579889 463390 584800 463392
rect 579889 463387 579955 463390
rect 583600 463300 584800 463390
rect -800 452434 400 452524
rect 3049 452434 3115 452437
rect -800 452432 3115 452434
rect -800 452376 3054 452432
rect 3110 452376 3115 452432
rect -800 452374 3115 452376
rect -800 452284 400 452374
rect 3049 452371 3115 452374
rect 579889 451754 579955 451757
rect 583600 451754 584800 451844
rect 579889 451752 584800 451754
rect 579889 451696 579894 451752
rect 579950 451696 584800 451752
rect 579889 451694 584800 451696
rect 579889 451691 579955 451694
rect 583600 451604 584800 451694
rect 579889 439922 579955 439925
rect 583600 439922 584800 440012
rect 579889 439920 584800 439922
rect 579889 439864 579894 439920
rect 579950 439864 584800 439920
rect 579889 439862 584800 439864
rect 579889 439859 579955 439862
rect 583600 439772 584800 439862
rect -800 438018 400 438108
rect 3141 438018 3207 438021
rect -800 438016 3207 438018
rect -800 437960 3146 438016
rect 3202 437960 3207 438016
rect -800 437958 3207 437960
rect -800 437868 400 437958
rect 3141 437955 3207 437958
rect 583600 428076 584800 428316
rect -800 423738 400 423828
rect 3141 423738 3207 423741
rect -800 423736 3207 423738
rect -800 423680 3146 423736
rect 3202 423680 3207 423736
rect -800 423678 3207 423680
rect -800 423588 400 423678
rect 3141 423675 3207 423678
rect 579889 416530 579955 416533
rect 583600 416530 584800 416620
rect 579889 416528 584800 416530
rect 579889 416472 579894 416528
rect 579950 416472 584800 416528
rect 579889 416470 584800 416472
rect 579889 416467 579955 416470
rect 583600 416380 584800 416470
rect -800 409172 400 409412
rect 579889 404834 579955 404837
rect 583600 404834 584800 404924
rect 579889 404832 584800 404834
rect 579889 404776 579894 404832
rect 579950 404776 584800 404832
rect 579889 404774 584800 404776
rect 579889 404771 579955 404774
rect 583600 404684 584800 404774
rect -800 395042 400 395132
rect 3233 395042 3299 395045
rect -800 395040 3299 395042
rect -800 394984 3238 395040
rect 3294 394984 3299 395040
rect -800 394982 3299 394984
rect -800 394892 400 394982
rect 3233 394979 3299 394982
rect 579889 393002 579955 393005
rect 583600 393002 584800 393092
rect 579889 393000 584800 393002
rect 579889 392944 579894 393000
rect 579950 392944 584800 393000
rect 579889 392942 584800 392944
rect 579889 392939 579955 392942
rect 583600 392852 584800 392942
rect 583600 381156 584800 381396
rect -800 380626 400 380716
rect 2773 380626 2839 380629
rect -800 380624 2839 380626
rect -800 380568 2778 380624
rect 2834 380568 2839 380624
rect -800 380566 2839 380568
rect -800 380476 400 380566
rect 2773 380563 2839 380566
rect 579889 369610 579955 369613
rect 583600 369610 584800 369700
rect 579889 369608 584800 369610
rect 579889 369552 579894 369608
rect 579950 369552 584800 369608
rect 579889 369550 584800 369552
rect 579889 369547 579955 369550
rect 583600 369460 584800 369550
rect -800 366210 400 366300
rect 2773 366210 2839 366213
rect -800 366208 2839 366210
rect -800 366152 2778 366208
rect 2834 366152 2839 366208
rect -800 366150 2839 366152
rect -800 366060 400 366150
rect 2773 366147 2839 366150
rect 580073 357914 580139 357917
rect 583600 357914 584800 358004
rect 580073 357912 584800 357914
rect 580073 357856 580078 357912
rect 580134 357856 584800 357912
rect 580073 357854 584800 357856
rect 580073 357851 580139 357854
rect 583600 357764 584800 357854
rect -800 351780 400 352020
rect 580073 346082 580139 346085
rect 583600 346082 584800 346172
rect 580073 346080 584800 346082
rect 580073 346024 580078 346080
rect 580134 346024 584800 346080
rect 580073 346022 584800 346024
rect 580073 346019 580139 346022
rect 583600 345932 584800 346022
rect -800 337514 400 337604
rect 3325 337514 3391 337517
rect -800 337512 3391 337514
rect -800 337456 3330 337512
rect 3386 337456 3391 337512
rect -800 337454 3391 337456
rect -800 337364 400 337454
rect 3325 337451 3391 337454
rect 583600 334236 584800 334476
rect -800 323098 400 323188
rect 3141 323098 3207 323101
rect -800 323096 3207 323098
rect -800 323040 3146 323096
rect 3202 323040 3207 323096
rect -800 323038 3207 323040
rect -800 322948 400 323038
rect 3141 323035 3207 323038
rect 580073 322690 580139 322693
rect 583600 322690 584800 322780
rect 580073 322688 584800 322690
rect 580073 322632 580078 322688
rect 580134 322632 584800 322688
rect 580073 322630 584800 322632
rect 580073 322627 580139 322630
rect 583600 322540 584800 322630
rect 368974 310796 368980 310860
rect 369044 310858 369050 310860
rect 583385 310858 583451 310861
rect 583600 310858 584800 310948
rect 369044 310798 374010 310858
rect 369044 310796 369050 310798
rect 373950 310722 374010 310798
rect 383702 310798 393330 310858
rect 373950 310662 383578 310722
rect 383518 310586 383578 310662
rect 383702 310586 383762 310798
rect 393270 310722 393330 310798
rect 403022 310798 412650 310858
rect 393270 310662 402898 310722
rect 383518 310526 383762 310586
rect 402838 310586 402898 310662
rect 403022 310586 403082 310798
rect 412590 310722 412650 310798
rect 422342 310798 431970 310858
rect 412590 310662 422218 310722
rect 402838 310526 403082 310586
rect 422158 310586 422218 310662
rect 422342 310586 422402 310798
rect 431910 310722 431970 310798
rect 441662 310798 451290 310858
rect 431910 310662 441538 310722
rect 422158 310526 422402 310586
rect 441478 310586 441538 310662
rect 441662 310586 441722 310798
rect 451230 310722 451290 310798
rect 460982 310798 470610 310858
rect 451230 310662 460858 310722
rect 441478 310526 441722 310586
rect 460798 310586 460858 310662
rect 460982 310586 461042 310798
rect 470550 310722 470610 310798
rect 480302 310798 489930 310858
rect 470550 310662 480178 310722
rect 460798 310526 461042 310586
rect 480118 310586 480178 310662
rect 480302 310586 480362 310798
rect 489870 310722 489930 310798
rect 499622 310798 509250 310858
rect 489870 310662 499498 310722
rect 480118 310526 480362 310586
rect 499438 310586 499498 310662
rect 499622 310586 499682 310798
rect 509190 310722 509250 310798
rect 518942 310798 528570 310858
rect 509190 310662 518818 310722
rect 499438 310526 499682 310586
rect 518758 310586 518818 310662
rect 518942 310586 519002 310798
rect 528510 310722 528570 310798
rect 538262 310798 547890 310858
rect 528510 310662 538138 310722
rect 518758 310526 519002 310586
rect 538078 310586 538138 310662
rect 538262 310586 538322 310798
rect 547830 310722 547890 310798
rect 557582 310798 567210 310858
rect 547830 310662 557458 310722
rect 538078 310526 538322 310586
rect 557398 310586 557458 310662
rect 557582 310586 557642 310798
rect 567150 310722 567210 310798
rect 583385 310856 584800 310858
rect 583385 310800 583390 310856
rect 583446 310800 584800 310856
rect 583385 310798 584800 310800
rect 583385 310795 583451 310798
rect 583385 310722 583451 310725
rect 567150 310662 576778 310722
rect 557398 310526 557642 310586
rect 576718 310586 576778 310662
rect 576902 310720 583451 310722
rect 576902 310664 583390 310720
rect 583446 310664 583451 310720
rect 583600 310708 584800 310798
rect 576902 310662 583451 310664
rect 576902 310586 576962 310662
rect 583385 310659 583451 310662
rect 576718 310526 576962 310586
rect -800 308818 400 308908
rect 4061 308818 4127 308821
rect -800 308816 4127 308818
rect -800 308760 4066 308816
rect 4122 308760 4127 308816
rect -800 308758 4127 308760
rect -800 308668 400 308758
rect 4061 308755 4127 308758
rect 576853 299298 576919 299301
rect 583385 299298 583451 299301
rect 576853 299296 583451 299298
rect 576853 299240 576858 299296
rect 576914 299240 583390 299296
rect 583446 299240 583451 299296
rect 576853 299238 583451 299240
rect 576853 299235 576919 299238
rect 583385 299235 583451 299238
rect 583385 299162 583451 299165
rect 583600 299162 584800 299252
rect 583385 299160 584800 299162
rect 583385 299104 583390 299160
rect 583446 299104 584800 299160
rect 583385 299102 584800 299104
rect 583385 299099 583451 299102
rect 583600 299012 584800 299102
rect 364382 298422 374010 298482
rect 359590 298148 359596 298212
rect 359660 298210 359666 298212
rect 364382 298210 364442 298422
rect 373950 298346 374010 298422
rect 383702 298422 393330 298482
rect 373950 298286 383578 298346
rect 359660 298150 364442 298210
rect 383518 298210 383578 298286
rect 383702 298210 383762 298422
rect 393270 298346 393330 298422
rect 403022 298422 412650 298482
rect 393270 298286 402898 298346
rect 383518 298150 383762 298210
rect 402838 298210 402898 298286
rect 403022 298210 403082 298422
rect 412590 298346 412650 298422
rect 422342 298422 431970 298482
rect 412590 298286 422218 298346
rect 402838 298150 403082 298210
rect 422158 298210 422218 298286
rect 422342 298210 422402 298422
rect 431910 298346 431970 298422
rect 441662 298422 451290 298482
rect 431910 298286 441538 298346
rect 422158 298150 422402 298210
rect 441478 298210 441538 298286
rect 441662 298210 441722 298422
rect 451230 298346 451290 298422
rect 460982 298422 470610 298482
rect 451230 298286 460858 298346
rect 441478 298150 441722 298210
rect 460798 298210 460858 298286
rect 460982 298210 461042 298422
rect 470550 298346 470610 298422
rect 480302 298422 489930 298482
rect 470550 298286 480178 298346
rect 460798 298150 461042 298210
rect 480118 298210 480178 298286
rect 480302 298210 480362 298422
rect 489870 298346 489930 298422
rect 499622 298422 509250 298482
rect 489870 298286 499498 298346
rect 480118 298150 480362 298210
rect 499438 298210 499498 298286
rect 499622 298210 499682 298422
rect 509190 298346 509250 298422
rect 518942 298422 528570 298482
rect 509190 298286 518818 298346
rect 499438 298150 499682 298210
rect 518758 298210 518818 298286
rect 518942 298210 519002 298422
rect 528510 298346 528570 298422
rect 538262 298422 547890 298482
rect 528510 298286 538138 298346
rect 518758 298150 519002 298210
rect 538078 298210 538138 298286
rect 538262 298210 538322 298422
rect 547830 298346 547890 298422
rect 557582 298422 567210 298482
rect 547830 298286 557458 298346
rect 538078 298150 538322 298210
rect 557398 298210 557458 298286
rect 557582 298210 557642 298422
rect 567150 298346 567210 298422
rect 567150 298286 576778 298346
rect 557398 298150 557642 298210
rect 576718 298210 576778 298286
rect 576853 298210 576919 298213
rect 576718 298208 576919 298210
rect 576718 298152 576858 298208
rect 576914 298152 576919 298208
rect 576718 298150 576919 298152
rect 359660 298148 359666 298150
rect 576853 298147 576919 298150
rect -800 294402 400 294492
rect 3969 294402 4035 294405
rect -800 294400 4035 294402
rect -800 294344 3974 294400
rect 4030 294344 4035 294400
rect -800 294342 4035 294344
rect -800 294252 400 294342
rect 3969 294339 4035 294342
rect 583600 287316 584800 287556
rect -800 280122 400 280212
rect 3325 280122 3391 280125
rect -800 280120 3391 280122
rect -800 280064 3330 280120
rect 3386 280064 3391 280120
rect -800 280062 3391 280064
rect -800 279972 400 280062
rect 3325 280059 3391 280062
rect 579613 275770 579679 275773
rect 583600 275770 584800 275860
rect 579613 275768 584800 275770
rect 579613 275712 579618 275768
rect 579674 275712 584800 275768
rect 579613 275710 584800 275712
rect 579613 275707 579679 275710
rect 583600 275620 584800 275710
rect -800 265706 400 265796
rect 2773 265706 2839 265709
rect -800 265704 2839 265706
rect -800 265648 2778 265704
rect 2834 265648 2839 265704
rect -800 265646 2839 265648
rect -800 265556 400 265646
rect 2773 265643 2839 265646
rect 579797 263938 579863 263941
rect 583600 263938 584800 264028
rect 579797 263936 584800 263938
rect 579797 263880 579802 263936
rect 579858 263880 584800 263936
rect 579797 263878 584800 263880
rect 579797 263875 579863 263878
rect 583600 263788 584800 263878
rect 576853 252378 576919 252381
rect 583385 252378 583451 252381
rect 576853 252376 583451 252378
rect 576853 252320 576858 252376
rect 576914 252320 583390 252376
rect 583446 252320 583451 252376
rect 576853 252318 583451 252320
rect 576853 252315 576919 252318
rect 583385 252315 583451 252318
rect 583385 252242 583451 252245
rect 583600 252242 584800 252332
rect 583385 252240 584800 252242
rect 583385 252184 583390 252240
rect 583446 252184 584800 252240
rect 583385 252182 584800 252184
rect 583385 252179 583451 252182
rect 583600 252092 584800 252182
rect 364382 251502 374010 251562
rect -800 251290 400 251380
rect 3877 251290 3943 251293
rect -800 251288 3943 251290
rect -800 251232 3882 251288
rect 3938 251232 3943 251288
rect -800 251230 3943 251232
rect -800 251140 400 251230
rect 3877 251227 3943 251230
rect 359406 251228 359412 251292
rect 359476 251290 359482 251292
rect 364382 251290 364442 251502
rect 373950 251426 374010 251502
rect 383702 251502 393330 251562
rect 373950 251366 383578 251426
rect 359476 251230 364442 251290
rect 383518 251290 383578 251366
rect 383702 251290 383762 251502
rect 393270 251426 393330 251502
rect 403022 251502 412650 251562
rect 393270 251366 402898 251426
rect 383518 251230 383762 251290
rect 402838 251290 402898 251366
rect 403022 251290 403082 251502
rect 412590 251426 412650 251502
rect 422342 251502 431970 251562
rect 412590 251366 422218 251426
rect 402838 251230 403082 251290
rect 422158 251290 422218 251366
rect 422342 251290 422402 251502
rect 431910 251426 431970 251502
rect 441662 251502 451290 251562
rect 431910 251366 441538 251426
rect 422158 251230 422402 251290
rect 441478 251290 441538 251366
rect 441662 251290 441722 251502
rect 451230 251426 451290 251502
rect 460982 251502 470610 251562
rect 451230 251366 460858 251426
rect 441478 251230 441722 251290
rect 460798 251290 460858 251366
rect 460982 251290 461042 251502
rect 470550 251426 470610 251502
rect 480302 251502 489930 251562
rect 470550 251366 480178 251426
rect 460798 251230 461042 251290
rect 480118 251290 480178 251366
rect 480302 251290 480362 251502
rect 489870 251426 489930 251502
rect 499622 251502 509250 251562
rect 489870 251366 499498 251426
rect 480118 251230 480362 251290
rect 499438 251290 499498 251366
rect 499622 251290 499682 251502
rect 509190 251426 509250 251502
rect 518942 251502 528570 251562
rect 509190 251366 518818 251426
rect 499438 251230 499682 251290
rect 518758 251290 518818 251366
rect 518942 251290 519002 251502
rect 528510 251426 528570 251502
rect 538262 251502 547890 251562
rect 528510 251366 538138 251426
rect 518758 251230 519002 251290
rect 538078 251290 538138 251366
rect 538262 251290 538322 251502
rect 547830 251426 547890 251502
rect 557582 251502 567210 251562
rect 547830 251366 557458 251426
rect 538078 251230 538322 251290
rect 557398 251290 557458 251366
rect 557582 251290 557642 251502
rect 567150 251426 567210 251502
rect 567150 251366 576778 251426
rect 557398 251230 557642 251290
rect 576718 251290 576778 251366
rect 576853 251290 576919 251293
rect 576718 251288 576919 251290
rect 576718 251232 576858 251288
rect 576914 251232 576919 251288
rect 576718 251230 576919 251232
rect 359476 251228 359482 251230
rect 576853 251227 576919 251230
rect 583600 240396 584800 240636
rect -800 237010 400 237100
rect 3325 237010 3391 237013
rect -800 237008 3391 237010
rect -800 236952 3330 237008
rect 3386 236952 3391 237008
rect -800 236950 3391 236952
rect -800 236860 400 236950
rect 3325 236947 3391 236950
rect 579981 228850 580047 228853
rect 583600 228850 584800 228940
rect 579981 228848 584800 228850
rect 579981 228792 579986 228848
rect 580042 228792 584800 228848
rect 579981 228790 584800 228792
rect 579981 228787 580047 228790
rect 583600 228700 584800 228790
rect -800 222594 400 222684
rect 3785 222594 3851 222597
rect -800 222592 3851 222594
rect -800 222536 3790 222592
rect 3846 222536 3851 222592
rect -800 222534 3851 222536
rect -800 222444 400 222534
rect 3785 222531 3851 222534
rect 275461 219602 275527 219605
rect 275461 219600 275938 219602
rect 275461 219544 275466 219600
rect 275522 219544 275938 219600
rect 275461 219542 275938 219544
rect 275461 219539 275527 219542
rect 275878 219469 275938 219542
rect 275829 219464 275938 219469
rect 275829 219408 275834 219464
rect 275890 219408 275938 219464
rect 275829 219406 275938 219408
rect 275829 219403 275895 219406
rect 275921 217972 275987 217973
rect 275870 217970 275876 217972
rect 275830 217910 275876 217970
rect 275940 217968 275987 217972
rect 275982 217912 275987 217968
rect 275870 217908 275876 217910
rect 275940 217908 275987 217912
rect 275921 217907 275987 217908
rect 331305 217834 331371 217837
rect 340781 217834 340847 217837
rect 331305 217832 340847 217834
rect 331305 217776 331310 217832
rect 331366 217776 340786 217832
rect 340842 217776 340847 217832
rect 331305 217774 340847 217776
rect 331305 217771 331371 217774
rect 340781 217771 340847 217774
rect 275921 217700 275987 217701
rect 275870 217698 275876 217700
rect 275830 217638 275876 217698
rect 275940 217696 275987 217700
rect 275982 217640 275987 217696
rect 275870 217636 275876 217638
rect 275940 217636 275987 217640
rect 275921 217635 275987 217636
rect 10317 217290 10383 217293
rect 172237 217290 172303 217293
rect 10317 217288 172303 217290
rect 10317 217232 10322 217288
rect 10378 217232 172242 217288
rect 172298 217232 172303 217288
rect 10317 217230 172303 217232
rect 10317 217227 10383 217230
rect 172237 217227 172303 217230
rect 331765 217290 331831 217293
rect 470593 217290 470659 217293
rect 331765 217288 470659 217290
rect 331765 217232 331770 217288
rect 331826 217232 470598 217288
rect 470654 217232 470659 217288
rect 331765 217230 470659 217232
rect 331765 217227 331831 217230
rect 470593 217227 470659 217230
rect 580165 217018 580231 217021
rect 583600 217018 584800 217108
rect 580165 217016 584800 217018
rect 580165 216960 580170 217016
rect 580226 216960 584800 217016
rect 580165 216958 584800 216960
rect 580165 216955 580231 216958
rect 583600 216868 584800 216958
rect 212349 212666 212415 212669
rect 212030 212664 212415 212666
rect 212030 212608 212354 212664
rect 212410 212608 212415 212664
rect 212030 212606 212415 212608
rect 211889 212564 211955 212567
rect 212030 212564 212090 212606
rect 212349 212603 212415 212606
rect 211889 212562 212090 212564
rect 173249 212530 173315 212533
rect 173433 212530 173499 212533
rect 173249 212528 173499 212530
rect 173249 212472 173254 212528
rect 173310 212472 173438 212528
rect 173494 212472 173499 212528
rect 211889 212506 211894 212562
rect 211950 212506 212090 212562
rect 211889 212504 212090 212506
rect 212165 212530 212231 212533
rect 212349 212530 212415 212533
rect 212165 212528 212415 212530
rect 211889 212501 211955 212504
rect 173249 212470 173499 212472
rect 173249 212467 173315 212470
rect 173433 212467 173499 212470
rect 212165 212472 212170 212528
rect 212226 212472 212354 212528
rect 212410 212472 212415 212528
rect 212165 212470 212415 212472
rect 212165 212467 212231 212470
rect 212349 212467 212415 212470
rect 229369 212530 229435 212533
rect 229553 212530 229619 212533
rect 229369 212528 229619 212530
rect 229369 212472 229374 212528
rect 229430 212472 229558 212528
rect 229614 212472 229619 212528
rect 229369 212470 229619 212472
rect 229369 212467 229435 212470
rect 229553 212467 229619 212470
rect 232037 212530 232103 212533
rect 232313 212530 232379 212533
rect 232037 212528 232379 212530
rect 232037 212472 232042 212528
rect 232098 212472 232318 212528
rect 232374 212472 232379 212528
rect 232037 212470 232379 212472
rect 232037 212467 232103 212470
rect 232313 212467 232379 212470
rect 289169 212530 289235 212533
rect 289353 212530 289419 212533
rect 289169 212528 289419 212530
rect 289169 212472 289174 212528
rect 289230 212472 289358 212528
rect 289414 212472 289419 212528
rect 289169 212470 289419 212472
rect 289169 212467 289235 212470
rect 289353 212467 289419 212470
rect 352833 212530 352899 212533
rect 353017 212530 353083 212533
rect 352833 212528 353083 212530
rect 352833 212472 352838 212528
rect 352894 212472 353022 212528
rect 353078 212472 353083 212528
rect 352833 212470 353083 212472
rect 352833 212467 352899 212470
rect 353017 212467 353083 212470
rect 217041 211170 217107 211173
rect 217961 211170 218027 211173
rect 217041 211168 218027 211170
rect 217041 211112 217046 211168
rect 217102 211112 217966 211168
rect 218022 211112 218027 211168
rect 217041 211110 218027 211112
rect 217041 211107 217107 211110
rect 217961 211107 218027 211110
rect 282453 211170 282519 211173
rect 282637 211170 282703 211173
rect 282453 211168 282703 211170
rect 282453 211112 282458 211168
rect 282514 211112 282642 211168
rect 282698 211112 282703 211168
rect 282453 211110 282703 211112
rect 282453 211107 282519 211110
rect 282637 211107 282703 211110
rect -800 208178 400 208268
rect 3693 208178 3759 208181
rect -800 208176 3759 208178
rect -800 208120 3698 208176
rect 3754 208120 3759 208176
rect -800 208118 3759 208120
rect -800 208028 400 208118
rect 3693 208115 3759 208118
rect 576853 205458 576919 205461
rect 583385 205458 583451 205461
rect 576853 205456 583451 205458
rect 576853 205400 576858 205456
rect 576914 205400 583390 205456
rect 583446 205400 583451 205456
rect 576853 205398 583451 205400
rect 576853 205395 576919 205398
rect 583385 205395 583451 205398
rect 583385 205322 583451 205325
rect 583600 205322 584800 205412
rect 583385 205320 584800 205322
rect 583385 205264 583390 205320
rect 583446 205264 584800 205320
rect 583385 205262 584800 205264
rect 583385 205259 583451 205262
rect 583600 205172 584800 205262
rect 366214 204580 366220 204644
rect 366284 204642 366290 204644
rect 366284 204582 374010 204642
rect 366284 204580 366290 204582
rect 373950 204506 374010 204582
rect 383702 204582 393330 204642
rect 373950 204446 383578 204506
rect 383518 204370 383578 204446
rect 383702 204370 383762 204582
rect 393270 204506 393330 204582
rect 403022 204582 412650 204642
rect 393270 204446 402898 204506
rect 383518 204310 383762 204370
rect 402838 204370 402898 204446
rect 403022 204370 403082 204582
rect 412590 204506 412650 204582
rect 422342 204582 431970 204642
rect 412590 204446 422218 204506
rect 402838 204310 403082 204370
rect 422158 204370 422218 204446
rect 422342 204370 422402 204582
rect 431910 204506 431970 204582
rect 441662 204582 451290 204642
rect 431910 204446 441538 204506
rect 422158 204310 422402 204370
rect 441478 204370 441538 204446
rect 441662 204370 441722 204582
rect 451230 204506 451290 204582
rect 460982 204582 470610 204642
rect 451230 204446 460858 204506
rect 441478 204310 441722 204370
rect 460798 204370 460858 204446
rect 460982 204370 461042 204582
rect 470550 204506 470610 204582
rect 480302 204582 489930 204642
rect 470550 204446 480178 204506
rect 460798 204310 461042 204370
rect 480118 204370 480178 204446
rect 480302 204370 480362 204582
rect 489870 204506 489930 204582
rect 499622 204582 509250 204642
rect 489870 204446 499498 204506
rect 480118 204310 480362 204370
rect 499438 204370 499498 204446
rect 499622 204370 499682 204582
rect 509190 204506 509250 204582
rect 518942 204582 528570 204642
rect 509190 204446 518818 204506
rect 499438 204310 499682 204370
rect 518758 204370 518818 204446
rect 518942 204370 519002 204582
rect 528510 204506 528570 204582
rect 538262 204582 547890 204642
rect 528510 204446 538138 204506
rect 518758 204310 519002 204370
rect 538078 204370 538138 204446
rect 538262 204370 538322 204582
rect 547830 204506 547890 204582
rect 557582 204582 567210 204642
rect 547830 204446 557458 204506
rect 538078 204310 538322 204370
rect 557398 204370 557458 204446
rect 557582 204370 557642 204582
rect 567150 204506 567210 204582
rect 567150 204446 576778 204506
rect 557398 204310 557642 204370
rect 576718 204370 576778 204446
rect 576853 204370 576919 204373
rect 576718 204368 576919 204370
rect 576718 204312 576858 204368
rect 576914 204312 576919 204368
rect 576718 204310 576919 204312
rect 576853 204307 576919 204310
rect 216673 202874 216739 202877
rect 216949 202874 217015 202877
rect 216673 202872 217015 202874
rect 216673 202816 216678 202872
rect 216734 202816 216954 202872
rect 217010 202816 217015 202872
rect 216673 202814 217015 202816
rect 216673 202811 216739 202814
rect 216949 202811 217015 202814
rect 286501 202874 286567 202877
rect 286685 202874 286751 202877
rect 286501 202872 286751 202874
rect 286501 202816 286506 202872
rect 286562 202816 286690 202872
rect 286746 202816 286751 202872
rect 286501 202814 286751 202816
rect 286501 202811 286567 202814
rect 286685 202811 286751 202814
rect 289261 202874 289327 202877
rect 289445 202874 289511 202877
rect 289261 202872 289511 202874
rect 289261 202816 289266 202872
rect 289322 202816 289450 202872
rect 289506 202816 289511 202872
rect 289261 202814 289511 202816
rect 289261 202811 289327 202814
rect 289445 202811 289511 202814
rect 276933 201514 276999 201517
rect 277209 201514 277275 201517
rect 276933 201512 277275 201514
rect 276933 201456 276938 201512
rect 276994 201456 277214 201512
rect 277270 201456 277275 201512
rect 276933 201454 277275 201456
rect 276933 201451 276999 201454
rect 277209 201451 277275 201454
rect 283833 201514 283899 201517
rect 284017 201514 284083 201517
rect 283833 201512 284083 201514
rect 283833 201456 283838 201512
rect 283894 201456 284022 201512
rect 284078 201456 284083 201512
rect 283833 201454 284083 201456
rect 283833 201451 283899 201454
rect 284017 201451 284083 201454
rect 341793 201514 341859 201517
rect 341977 201514 342043 201517
rect 341793 201512 342043 201514
rect 341793 201456 341798 201512
rect 341854 201456 341982 201512
rect 342038 201456 342043 201512
rect 341793 201454 342043 201456
rect 341793 201451 341859 201454
rect 341977 201451 342043 201454
rect 354121 201514 354187 201517
rect 354397 201514 354463 201517
rect 354121 201512 354463 201514
rect 354121 201456 354126 201512
rect 354182 201456 354402 201512
rect 354458 201456 354463 201512
rect 354121 201454 354463 201456
rect 354121 201451 354187 201454
rect 354397 201451 354463 201454
rect 355409 201514 355475 201517
rect 355685 201514 355751 201517
rect 355409 201512 355751 201514
rect 355409 201456 355414 201512
rect 355470 201456 355690 201512
rect 355746 201456 355751 201512
rect 355409 201454 355751 201456
rect 355409 201451 355475 201454
rect 355685 201451 355751 201454
rect 225137 200154 225203 200157
rect 225321 200154 225387 200157
rect 225137 200152 225387 200154
rect 225137 200096 225142 200152
rect 225198 200096 225326 200152
rect 225382 200096 225387 200152
rect 225137 200094 225387 200096
rect 225137 200091 225203 200094
rect 225321 200091 225387 200094
rect -800 193898 400 193988
rect 3141 193898 3207 193901
rect -800 193896 3207 193898
rect -800 193840 3146 193896
rect 3202 193840 3207 193896
rect -800 193838 3207 193840
rect -800 193748 400 193838
rect 3141 193835 3207 193838
rect 583600 193476 584800 193716
rect 219709 193218 219775 193221
rect 219985 193218 220051 193221
rect 219709 193216 220051 193218
rect 219709 193160 219714 193216
rect 219770 193160 219990 193216
rect 220046 193160 220051 193216
rect 219709 193158 220051 193160
rect 219709 193155 219775 193158
rect 219985 193155 220051 193158
rect 232037 193218 232103 193221
rect 232221 193218 232287 193221
rect 232037 193216 232287 193218
rect 232037 193160 232042 193216
rect 232098 193160 232226 193216
rect 232282 193160 232287 193216
rect 232037 193158 232287 193160
rect 232037 193155 232103 193158
rect 232221 193155 232287 193158
rect 289261 193218 289327 193221
rect 289445 193218 289511 193221
rect 289261 193216 289511 193218
rect 289261 193160 289266 193216
rect 289322 193160 289450 193216
rect 289506 193160 289511 193216
rect 289261 193158 289511 193160
rect 289261 193155 289327 193158
rect 289445 193155 289511 193158
rect 291653 193218 291719 193221
rect 291837 193218 291903 193221
rect 291653 193216 291903 193218
rect 291653 193160 291658 193216
rect 291714 193160 291842 193216
rect 291898 193160 291903 193216
rect 291653 193158 291903 193160
rect 291653 193155 291719 193158
rect 291837 193155 291903 193158
rect 343173 193218 343239 193221
rect 343357 193218 343423 193221
rect 343173 193216 343423 193218
rect 343173 193160 343178 193216
rect 343234 193160 343362 193216
rect 343418 193160 343423 193216
rect 343173 193158 343423 193160
rect 343173 193155 343239 193158
rect 343357 193155 343423 193158
rect 344369 193218 344435 193221
rect 344645 193218 344711 193221
rect 344369 193216 344711 193218
rect 344369 193160 344374 193216
rect 344430 193160 344650 193216
rect 344706 193160 344711 193216
rect 344369 193158 344711 193160
rect 344369 193155 344435 193158
rect 344645 193155 344711 193158
rect 354213 193218 354279 193221
rect 354397 193218 354463 193221
rect 354213 193216 354463 193218
rect 354213 193160 354218 193216
rect 354274 193160 354402 193216
rect 354458 193160 354463 193216
rect 354213 193158 354463 193160
rect 354213 193155 354279 193158
rect 354397 193155 354463 193158
rect 355409 193218 355475 193221
rect 355685 193218 355751 193221
rect 355409 193216 355751 193218
rect 355409 193160 355414 193216
rect 355470 193160 355690 193216
rect 355746 193160 355751 193216
rect 355409 193158 355751 193160
rect 355409 193155 355475 193158
rect 355685 193155 355751 193158
rect 285213 191994 285279 191997
rect 285213 191992 285322 191994
rect 285213 191936 285218 191992
rect 285274 191936 285322 191992
rect 285213 191931 285322 191936
rect 285262 191861 285322 191931
rect 184013 191858 184079 191861
rect 184289 191858 184355 191861
rect 184013 191856 184355 191858
rect 184013 191800 184018 191856
rect 184074 191800 184294 191856
rect 184350 191800 184355 191856
rect 184013 191798 184355 191800
rect 184013 191795 184079 191798
rect 184289 191795 184355 191798
rect 266537 191858 266603 191861
rect 266721 191858 266787 191861
rect 266537 191856 266787 191858
rect 266537 191800 266542 191856
rect 266598 191800 266726 191856
rect 266782 191800 266787 191856
rect 266537 191798 266787 191800
rect 285262 191856 285371 191861
rect 285262 191800 285310 191856
rect 285366 191800 285371 191856
rect 285262 191798 285371 191800
rect 266537 191795 266603 191798
rect 266721 191795 266787 191798
rect 285305 191795 285371 191798
rect 230841 190498 230907 190501
rect 231025 190498 231091 190501
rect 230841 190496 231091 190498
rect 230841 190440 230846 190496
rect 230902 190440 231030 190496
rect 231086 190440 231091 190496
rect 230841 190438 231091 190440
rect 230841 190435 230907 190438
rect 231025 190435 231091 190438
rect 216673 183562 216739 183565
rect 216949 183562 217015 183565
rect 216673 183560 217015 183562
rect 216673 183504 216678 183560
rect 216734 183504 216954 183560
rect 217010 183504 217015 183560
rect 216673 183502 217015 183504
rect 216673 183499 216739 183502
rect 216949 183499 217015 183502
rect 235073 183562 235139 183565
rect 235349 183562 235415 183565
rect 235073 183560 235415 183562
rect 235073 183504 235078 183560
rect 235134 183504 235354 183560
rect 235410 183504 235415 183560
rect 235073 183502 235415 183504
rect 235073 183499 235139 183502
rect 235349 183499 235415 183502
rect 282729 183562 282795 183565
rect 282913 183562 282979 183565
rect 286593 183562 286659 183565
rect 282729 183560 282979 183562
rect 282729 183504 282734 183560
rect 282790 183504 282918 183560
rect 282974 183504 282979 183560
rect 282729 183502 282979 183504
rect 282729 183499 282795 183502
rect 282913 183499 282979 183502
rect 286550 183560 286659 183562
rect 286550 183504 286598 183560
rect 286654 183504 286659 183560
rect 286550 183499 286659 183504
rect 289261 183562 289327 183565
rect 289445 183562 289511 183565
rect 289261 183560 289511 183562
rect 289261 183504 289266 183560
rect 289322 183504 289450 183560
rect 289506 183504 289511 183560
rect 289261 183502 289511 183504
rect 289261 183499 289327 183502
rect 289445 183499 289511 183502
rect 286550 183429 286610 183499
rect 286501 183424 286610 183429
rect 286501 183368 286506 183424
rect 286562 183368 286610 183424
rect 286501 183366 286610 183368
rect 286501 183363 286567 183366
rect 229277 182202 229343 182205
rect 229553 182202 229619 182205
rect 229277 182200 229619 182202
rect 229277 182144 229282 182200
rect 229338 182144 229558 182200
rect 229614 182144 229619 182200
rect 229277 182142 229619 182144
rect 229277 182139 229343 182142
rect 229553 182139 229619 182142
rect 283833 182202 283899 182205
rect 284017 182202 284083 182205
rect 283833 182200 284083 182202
rect 283833 182144 283838 182200
rect 283894 182144 284022 182200
rect 284078 182144 284083 182200
rect 283833 182142 284083 182144
rect 283833 182139 283899 182142
rect 284017 182139 284083 182142
rect 342989 182202 343055 182205
rect 343173 182202 343239 182205
rect 342989 182200 343239 182202
rect 342989 182144 342994 182200
rect 343050 182144 343178 182200
rect 343234 182144 343239 182200
rect 342989 182142 343239 182144
rect 342989 182139 343055 182142
rect 343173 182139 343239 182142
rect 580901 181930 580967 181933
rect 583600 181930 584800 182020
rect 580901 181928 584800 181930
rect 580901 181872 580906 181928
rect 580962 181872 584800 181928
rect 580901 181870 584800 181872
rect 580901 181867 580967 181870
rect 583600 181780 584800 181870
rect 225229 180842 225295 180845
rect 225505 180842 225571 180845
rect 225229 180840 225571 180842
rect 225229 180784 225234 180840
rect 225290 180784 225510 180840
rect 225566 180784 225571 180840
rect 225229 180782 225571 180784
rect 225229 180779 225295 180782
rect 225505 180779 225571 180782
rect -800 179482 400 179572
rect 3601 179482 3667 179485
rect -800 179480 3667 179482
rect -800 179424 3606 179480
rect 3662 179424 3667 179480
rect -800 179422 3667 179424
rect -800 179332 400 179422
rect 3601 179419 3667 179422
rect 328085 174042 328151 174045
rect 328269 174042 328335 174045
rect 328085 174040 328335 174042
rect 328085 173984 328090 174040
rect 328146 173984 328274 174040
rect 328330 173984 328335 174040
rect 328085 173982 328335 173984
rect 328085 173979 328151 173982
rect 328269 173979 328335 173982
rect 317045 173906 317111 173909
rect 317229 173906 317295 173909
rect 317045 173904 317295 173906
rect 317045 173848 317050 173904
rect 317106 173848 317234 173904
rect 317290 173848 317295 173904
rect 317045 173846 317295 173848
rect 317045 173843 317111 173846
rect 317229 173843 317295 173846
rect 272977 172682 273043 172685
rect 272934 172680 273043 172682
rect 272934 172624 272982 172680
rect 273038 172624 273043 172680
rect 272934 172619 273043 172624
rect 261109 172546 261175 172549
rect 261293 172546 261359 172549
rect 261109 172544 261359 172546
rect 261109 172488 261114 172544
rect 261170 172488 261298 172544
rect 261354 172488 261359 172544
rect 261109 172486 261359 172488
rect 272934 172546 272994 172619
rect 273069 172546 273135 172549
rect 272934 172544 273135 172546
rect 272934 172488 273074 172544
rect 273130 172488 273135 172544
rect 272934 172486 273135 172488
rect 261109 172483 261175 172486
rect 261293 172483 261359 172486
rect 273069 172483 273135 172486
rect 343173 172546 343239 172549
rect 343357 172546 343423 172549
rect 343173 172544 343423 172546
rect 343173 172488 343178 172544
rect 343234 172488 343362 172544
rect 343418 172488 343423 172544
rect 343173 172486 343423 172488
rect 343173 172483 343239 172486
rect 343357 172483 343423 172486
rect 344461 172546 344527 172549
rect 344645 172546 344711 172549
rect 344461 172544 344711 172546
rect 344461 172488 344466 172544
rect 344522 172488 344650 172544
rect 344706 172488 344711 172544
rect 344461 172486 344711 172488
rect 344461 172483 344527 172486
rect 344645 172483 344711 172486
rect 360929 172546 360995 172549
rect 361113 172546 361179 172549
rect 360929 172544 361179 172546
rect 360929 172488 360934 172544
rect 360990 172488 361118 172544
rect 361174 172488 361179 172544
rect 360929 172486 361179 172488
rect 360929 172483 360995 172486
rect 361113 172483 361179 172486
rect 580165 170098 580231 170101
rect 583600 170098 584800 170188
rect 580165 170096 584800 170098
rect 580165 170040 580170 170096
rect 580226 170040 584800 170096
rect 580165 170038 584800 170040
rect 580165 170035 580231 170038
rect 583600 169948 584800 170038
rect -800 165066 400 165156
rect 2773 165066 2839 165069
rect -800 165064 2839 165066
rect -800 165008 2778 165064
rect 2834 165008 2839 165064
rect -800 165006 2839 165008
rect -800 164916 400 165006
rect 2773 165003 2839 165006
rect 235165 164386 235231 164389
rect 235030 164384 235231 164386
rect 235030 164328 235170 164384
rect 235226 164328 235231 164384
rect 235030 164326 235231 164328
rect 235030 164253 235090 164326
rect 235165 164323 235231 164326
rect 235030 164248 235139 164253
rect 235030 164192 235078 164248
rect 235134 164192 235139 164248
rect 235030 164190 235139 164192
rect 235073 164187 235139 164190
rect 282637 164250 282703 164253
rect 282821 164250 282887 164253
rect 282637 164248 282887 164250
rect 282637 164192 282642 164248
rect 282698 164192 282826 164248
rect 282882 164192 282887 164248
rect 282637 164190 282887 164192
rect 282637 164187 282703 164190
rect 282821 164187 282887 164190
rect 327993 164250 328059 164253
rect 328177 164250 328243 164253
rect 327993 164248 328243 164250
rect 327993 164192 327998 164248
rect 328054 164192 328182 164248
rect 328238 164192 328243 164248
rect 327993 164190 328243 164192
rect 327993 164187 328059 164190
rect 328177 164187 328243 164190
rect 329281 164250 329347 164253
rect 329465 164250 329531 164253
rect 329281 164248 329531 164250
rect 329281 164192 329286 164248
rect 329342 164192 329470 164248
rect 329526 164192 329531 164248
rect 329281 164190 329531 164192
rect 329281 164187 329347 164190
rect 329465 164187 329531 164190
rect 277025 162890 277091 162893
rect 283833 162890 283899 162893
rect 284017 162890 284083 162893
rect 277025 162888 277226 162890
rect 277025 162832 277030 162888
rect 277086 162832 277226 162888
rect 277025 162830 277226 162832
rect 277025 162827 277091 162830
rect 277166 162756 277226 162830
rect 283833 162888 284083 162890
rect 283833 162832 283838 162888
rect 283894 162832 284022 162888
rect 284078 162832 284083 162888
rect 283833 162830 284083 162832
rect 283833 162827 283899 162830
rect 284017 162827 284083 162830
rect 345473 162890 345539 162893
rect 345657 162890 345723 162893
rect 345473 162888 345723 162890
rect 345473 162832 345478 162888
rect 345534 162832 345662 162888
rect 345718 162832 345723 162888
rect 345473 162830 345723 162832
rect 345473 162827 345539 162830
rect 345657 162827 345723 162830
rect 277158 162692 277164 162756
rect 277228 162692 277234 162756
rect 343265 160304 343331 160309
rect 343265 160248 343270 160304
rect 343326 160248 343331 160304
rect 343265 160243 343331 160248
rect 343268 160173 343328 160243
rect 343265 160168 343331 160173
rect 343265 160112 343270 160168
rect 343326 160112 343331 160168
rect 343265 160107 343331 160112
rect 580717 158402 580783 158405
rect 583600 158402 584800 158492
rect 580717 158400 584800 158402
rect 580717 158344 580722 158400
rect 580778 158344 584800 158400
rect 580717 158342 584800 158344
rect 580717 158339 580783 158342
rect 583600 158252 584800 158342
rect 191097 154730 191163 154733
rect 191054 154728 191163 154730
rect 191054 154672 191102 154728
rect 191158 154672 191163 154728
rect 191054 154667 191163 154672
rect 194961 154730 195027 154733
rect 200389 154730 200455 154733
rect 201861 154730 201927 154733
rect 194961 154728 195162 154730
rect 194961 154672 194966 154728
rect 195022 154672 195162 154728
rect 194961 154670 195162 154672
rect 194961 154667 195027 154670
rect 191054 154597 191114 154667
rect 171409 154594 171475 154597
rect 171593 154594 171659 154597
rect 171409 154592 171659 154594
rect 171409 154536 171414 154592
rect 171470 154536 171598 154592
rect 171654 154536 171659 154592
rect 171409 154534 171659 154536
rect 171409 154531 171475 154534
rect 171593 154531 171659 154534
rect 173065 154594 173131 154597
rect 173249 154594 173315 154597
rect 173065 154592 173315 154594
rect 173065 154536 173070 154592
rect 173126 154536 173254 154592
rect 173310 154536 173315 154592
rect 173065 154534 173315 154536
rect 191054 154592 191163 154597
rect 191054 154536 191102 154592
rect 191158 154536 191163 154592
rect 191054 154534 191163 154536
rect 173065 154531 173131 154534
rect 173249 154531 173315 154534
rect 191097 154531 191163 154534
rect 194961 154594 195027 154597
rect 195102 154594 195162 154670
rect 194961 154592 195162 154594
rect 194961 154536 194966 154592
rect 195022 154536 195162 154592
rect 194961 154534 195162 154536
rect 200254 154728 200455 154730
rect 200254 154672 200394 154728
rect 200450 154672 200455 154728
rect 200254 154670 200455 154672
rect 200254 154594 200314 154670
rect 200389 154667 200455 154670
rect 201726 154728 201927 154730
rect 201726 154672 201866 154728
rect 201922 154672 201927 154728
rect 201726 154670 201927 154672
rect 200389 154594 200455 154597
rect 200254 154592 200455 154594
rect 200254 154536 200394 154592
rect 200450 154536 200455 154592
rect 200254 154534 200455 154536
rect 201726 154594 201786 154670
rect 201861 154667 201927 154670
rect 201861 154594 201927 154597
rect 201726 154592 201927 154594
rect 201726 154536 201866 154592
rect 201922 154536 201927 154592
rect 201726 154534 201927 154536
rect 194961 154531 195027 154534
rect 200389 154531 200455 154534
rect 201861 154531 201927 154534
rect 230933 154594 230999 154597
rect 231209 154594 231275 154597
rect 230933 154592 231275 154594
rect 230933 154536 230938 154592
rect 230994 154536 231214 154592
rect 231270 154536 231275 154592
rect 230933 154534 231275 154536
rect 230933 154531 230999 154534
rect 231209 154531 231275 154534
rect 262305 154594 262371 154597
rect 262581 154594 262647 154597
rect 262305 154592 262647 154594
rect 262305 154536 262310 154592
rect 262366 154536 262586 154592
rect 262642 154536 262647 154592
rect 262305 154534 262647 154536
rect 262305 154531 262371 154534
rect 262581 154531 262647 154534
rect 277117 153236 277183 153237
rect 277117 153234 277164 153236
rect 277072 153232 277164 153234
rect 277072 153176 277122 153232
rect 277072 153174 277164 153176
rect 277117 153172 277164 153174
rect 277228 153172 277234 153236
rect 289261 153234 289327 153237
rect 289445 153234 289511 153237
rect 289261 153232 289511 153234
rect 289261 153176 289266 153232
rect 289322 153176 289450 153232
rect 289506 153176 289511 153232
rect 289261 153174 289511 153176
rect 277117 153171 277183 153172
rect 289261 153171 289327 153174
rect 289445 153171 289511 153174
rect -800 150786 400 150876
rect 3325 150786 3391 150789
rect -800 150784 3391 150786
rect -800 150728 3330 150784
rect 3386 150728 3391 150784
rect -800 150726 3391 150728
rect -800 150636 400 150726
rect 3325 150723 3391 150726
rect 318517 147796 318583 147797
rect 329557 147796 329623 147797
rect 318517 147792 318564 147796
rect 318628 147794 318634 147796
rect 318517 147736 318522 147792
rect 318517 147732 318564 147736
rect 318628 147734 318674 147794
rect 329557 147792 329604 147796
rect 329668 147794 329674 147796
rect 329557 147736 329562 147792
rect 318628 147732 318634 147734
rect 329557 147732 329604 147736
rect 329668 147734 329714 147794
rect 329668 147732 329674 147734
rect 318517 147731 318583 147732
rect 329557 147731 329623 147732
rect 583600 146556 584800 146796
rect 329557 144940 329623 144941
rect 329557 144936 329604 144940
rect 329668 144938 329674 144940
rect 355501 144938 355567 144941
rect 355685 144938 355751 144941
rect 329557 144880 329562 144936
rect 329557 144876 329604 144880
rect 329668 144878 329714 144938
rect 355501 144936 355751 144938
rect 355501 144880 355506 144936
rect 355562 144880 355690 144936
rect 355746 144880 355751 144936
rect 355501 144878 355751 144880
rect 329668 144876 329674 144878
rect 329557 144875 329623 144876
rect 355501 144875 355567 144878
rect 355685 144875 355751 144878
rect 194961 143580 195027 143581
rect 194910 143578 194916 143580
rect 194870 143518 194916 143578
rect 194980 143576 195027 143580
rect 195022 143520 195027 143576
rect 194910 143516 194916 143518
rect 194980 143516 195027 143520
rect 194961 143515 195027 143516
rect 231761 143578 231827 143581
rect 232037 143578 232103 143581
rect 231761 143576 232103 143578
rect 231761 143520 231766 143576
rect 231822 143520 232042 143576
rect 232098 143520 232103 143576
rect 231761 143518 232103 143520
rect 231761 143515 231827 143518
rect 232037 143515 232103 143518
rect 277025 143578 277091 143581
rect 277209 143578 277275 143581
rect 277025 143576 277275 143578
rect 277025 143520 277030 143576
rect 277086 143520 277214 143576
rect 277270 143520 277275 143576
rect 277025 143518 277275 143520
rect 277025 143515 277091 143518
rect 277209 143515 277275 143518
rect 318517 143580 318583 143581
rect 318517 143576 318564 143580
rect 318628 143578 318634 143580
rect 318517 143520 318522 143576
rect 318517 143516 318564 143520
rect 318628 143518 318674 143578
rect 318628 143516 318634 143518
rect 318517 143515 318583 143516
rect 194961 142220 195027 142221
rect 194910 142156 194916 142220
rect 194980 142218 195027 142220
rect 194980 142216 195072 142218
rect 195022 142160 195072 142216
rect 194980 142158 195072 142160
rect 194980 142156 195027 142158
rect 194961 142155 195027 142156
rect 225321 140722 225387 140725
rect 225505 140722 225571 140725
rect 225321 140720 225571 140722
rect 225321 140664 225326 140720
rect 225382 140664 225510 140720
rect 225566 140664 225571 140720
rect 225321 140662 225571 140664
rect 225321 140659 225387 140662
rect 225505 140659 225571 140662
rect 228265 139362 228331 139365
rect 228449 139362 228515 139365
rect 228265 139360 228515 139362
rect 228265 139304 228270 139360
rect 228326 139304 228454 139360
rect 228510 139304 228515 139360
rect 228265 139302 228515 139304
rect 228265 139299 228331 139302
rect 228449 139299 228515 139302
rect 234981 138002 235047 138005
rect 235257 138002 235323 138005
rect 234981 138000 235323 138002
rect 234981 137944 234986 138000
rect 235042 137944 235262 138000
rect 235318 137944 235323 138000
rect 234981 137942 235323 137944
rect 234981 137939 235047 137942
rect 235257 137939 235323 137942
rect -800 136370 400 136460
rect 2773 136370 2839 136373
rect -800 136368 2839 136370
rect -800 136312 2778 136368
rect 2834 136312 2839 136368
rect -800 136310 2839 136312
rect -800 136220 400 136310
rect 2773 136307 2839 136310
rect 200389 135418 200455 135421
rect 201861 135418 201927 135421
rect 200389 135416 200498 135418
rect 200389 135360 200394 135416
rect 200450 135360 200498 135416
rect 200389 135355 200498 135360
rect 201861 135416 201970 135418
rect 201861 135360 201866 135416
rect 201922 135360 201970 135416
rect 201861 135355 201970 135360
rect 200438 135285 200498 135355
rect 201910 135285 201970 135355
rect 171409 135282 171475 135285
rect 171593 135282 171659 135285
rect 171409 135280 171659 135282
rect 171409 135224 171414 135280
rect 171470 135224 171598 135280
rect 171654 135224 171659 135280
rect 171409 135222 171659 135224
rect 171409 135219 171475 135222
rect 171593 135219 171659 135222
rect 173065 135282 173131 135285
rect 173249 135282 173315 135285
rect 173065 135280 173315 135282
rect 173065 135224 173070 135280
rect 173126 135224 173254 135280
rect 173310 135224 173315 135280
rect 173065 135222 173315 135224
rect 173065 135219 173131 135222
rect 173249 135219 173315 135222
rect 200389 135280 200498 135285
rect 200389 135224 200394 135280
rect 200450 135224 200498 135280
rect 200389 135222 200498 135224
rect 201861 135280 201970 135285
rect 201861 135224 201866 135280
rect 201922 135224 201970 135280
rect 201861 135222 201970 135224
rect 262305 135282 262371 135285
rect 262581 135282 262647 135285
rect 262305 135280 262647 135282
rect 262305 135224 262310 135280
rect 262366 135224 262586 135280
rect 262642 135224 262647 135280
rect 262305 135222 262647 135224
rect 200389 135219 200455 135222
rect 201861 135219 201927 135222
rect 262305 135219 262371 135222
rect 262581 135219 262647 135222
rect 580533 134874 580599 134877
rect 583600 134874 584800 134964
rect 580533 134872 584800 134874
rect 580533 134816 580538 134872
rect 580594 134816 584800 134872
rect 580533 134814 584800 134816
rect 580533 134811 580599 134814
rect 583600 134724 584800 134814
rect 291837 134058 291903 134061
rect 291837 134056 291946 134058
rect 291837 134000 291842 134056
rect 291898 134000 291946 134056
rect 291837 133995 291946 134000
rect 291886 133925 291946 133995
rect 219801 133922 219867 133925
rect 219985 133922 220051 133925
rect 219801 133920 220051 133922
rect 219801 133864 219806 133920
rect 219862 133864 219990 133920
rect 220046 133864 220051 133920
rect 219801 133862 220051 133864
rect 219801 133859 219867 133862
rect 219985 133859 220051 133862
rect 224033 133922 224099 133925
rect 224217 133922 224283 133925
rect 224033 133920 224283 133922
rect 224033 133864 224038 133920
rect 224094 133864 224222 133920
rect 224278 133864 224283 133920
rect 224033 133862 224283 133864
rect 291886 133920 291995 133925
rect 291886 133864 291934 133920
rect 291990 133864 291995 133920
rect 291886 133862 291995 133864
rect 224033 133859 224099 133862
rect 224217 133859 224283 133862
rect 291929 133859 291995 133862
rect 345657 132562 345723 132565
rect 345841 132562 345907 132565
rect 345657 132560 345907 132562
rect 345657 132504 345662 132560
rect 345718 132504 345846 132560
rect 345902 132504 345907 132560
rect 345657 132502 345907 132504
rect 345657 132499 345723 132502
rect 345841 132499 345907 132502
rect 329557 128484 329623 128485
rect 329557 128480 329604 128484
rect 329668 128482 329674 128484
rect 329557 128424 329562 128480
rect 329557 128420 329604 128424
rect 329668 128422 329714 128482
rect 329668 128420 329674 128422
rect 329557 128419 329623 128420
rect 229369 125762 229435 125765
rect 235165 125762 235231 125765
rect 229326 125760 229435 125762
rect 229326 125704 229374 125760
rect 229430 125704 229435 125760
rect 229326 125699 229435 125704
rect 235030 125760 235231 125762
rect 235030 125704 235170 125760
rect 235226 125704 235231 125760
rect 235030 125702 235231 125704
rect 229326 125629 229386 125699
rect 229277 125624 229386 125629
rect 229277 125568 229282 125624
rect 229338 125568 229386 125624
rect 229277 125566 229386 125568
rect 235030 125629 235090 125702
rect 235165 125699 235231 125702
rect 235030 125624 235139 125629
rect 235030 125568 235078 125624
rect 235134 125568 235139 125624
rect 235030 125566 235139 125568
rect 229277 125563 229343 125566
rect 235073 125563 235139 125566
rect 329557 125628 329623 125629
rect 329557 125624 329604 125628
rect 329668 125626 329674 125628
rect 329557 125568 329562 125624
rect 329557 125564 329604 125568
rect 329668 125566 329714 125626
rect 329668 125564 329674 125566
rect 329557 125563 329623 125564
rect 284293 124266 284359 124269
rect 284020 124264 284359 124266
rect 284020 124208 284298 124264
rect 284354 124208 284359 124264
rect 284020 124206 284359 124208
rect 284020 123996 284080 124206
rect 284293 124203 284359 124206
rect 291745 124266 291811 124269
rect 291929 124266 291995 124269
rect 291745 124264 291995 124266
rect 291745 124208 291750 124264
rect 291806 124208 291934 124264
rect 291990 124208 291995 124264
rect 291745 124206 291995 124208
rect 291745 124203 291811 124206
rect 291929 124203 291995 124206
rect 283966 123932 283972 123996
rect 284036 123934 284080 123996
rect 284036 123932 284042 123934
rect 580809 123178 580875 123181
rect 583600 123178 584800 123268
rect 580809 123176 584800 123178
rect 580809 123120 580814 123176
rect 580870 123120 584800 123176
rect 580809 123118 584800 123120
rect 580809 123115 580875 123118
rect 583600 123028 584800 123118
rect 362309 122906 362375 122909
rect 362585 122906 362651 122909
rect 362309 122904 362651 122906
rect 362309 122848 362314 122904
rect 362370 122848 362590 122904
rect 362646 122848 362651 122904
rect 362309 122846 362651 122848
rect 362309 122843 362375 122846
rect 362585 122843 362651 122846
rect -800 122090 400 122180
rect 2773 122090 2839 122093
rect -800 122088 2839 122090
rect -800 122032 2778 122088
rect 2834 122032 2839 122088
rect -800 122030 2839 122032
rect -800 121940 400 122030
rect 2773 122027 2839 122030
rect 189441 116106 189507 116109
rect 189398 116104 189507 116106
rect 189398 116048 189446 116104
rect 189502 116048 189507 116104
rect 189398 116043 189507 116048
rect 189398 115973 189458 116043
rect 189349 115968 189458 115973
rect 189349 115912 189354 115968
rect 189410 115912 189458 115968
rect 189349 115910 189458 115912
rect 262305 115970 262371 115973
rect 262581 115970 262647 115973
rect 262305 115968 262647 115970
rect 262305 115912 262310 115968
rect 262366 115912 262586 115968
rect 262642 115912 262647 115968
rect 262305 115910 262647 115912
rect 189349 115907 189415 115910
rect 262305 115907 262371 115910
rect 262581 115907 262647 115910
rect 580625 111482 580691 111485
rect 583600 111482 584800 111572
rect 580625 111480 584800 111482
rect 580625 111424 580630 111480
rect 580686 111424 584800 111480
rect 580625 111422 584800 111424
rect 580625 111419 580691 111422
rect 583600 111332 584800 111422
rect 329557 109172 329623 109173
rect 329557 109168 329604 109172
rect 329668 109170 329674 109172
rect 329557 109112 329562 109168
rect 329557 109108 329604 109112
rect 329668 109110 329714 109170
rect 329668 109108 329674 109110
rect 329557 109107 329623 109108
rect -800 107674 400 107764
rect 3325 107674 3391 107677
rect -800 107672 3391 107674
rect -800 107616 3330 107672
rect 3386 107616 3391 107672
rect -800 107614 3391 107616
rect -800 107524 400 107614
rect 3325 107611 3391 107614
rect 191097 106450 191163 106453
rect 235165 106450 235231 106453
rect 191054 106448 191163 106450
rect 191054 106392 191102 106448
rect 191158 106392 191163 106448
rect 191054 106387 191163 106392
rect 235030 106448 235231 106450
rect 235030 106392 235170 106448
rect 235226 106392 235231 106448
rect 235030 106390 235231 106392
rect 191054 106317 191114 106387
rect 191005 106312 191114 106317
rect 191005 106256 191010 106312
rect 191066 106256 191114 106312
rect 191005 106254 191114 106256
rect 235030 106317 235090 106390
rect 235165 106387 235231 106390
rect 361205 106450 361271 106453
rect 361205 106448 361498 106450
rect 361205 106392 361210 106448
rect 361266 106392 361498 106448
rect 361205 106390 361498 106392
rect 361205 106387 361271 106390
rect 235030 106312 235139 106317
rect 284017 106316 284083 106317
rect 235030 106256 235078 106312
rect 235134 106256 235139 106312
rect 235030 106254 235139 106256
rect 191005 106251 191071 106254
rect 235073 106251 235139 106254
rect 283966 106252 283972 106316
rect 284036 106314 284083 106316
rect 286409 106314 286475 106317
rect 286593 106314 286659 106317
rect 284036 106312 284128 106314
rect 284078 106256 284128 106312
rect 284036 106254 284128 106256
rect 286409 106312 286659 106314
rect 286409 106256 286414 106312
rect 286470 106256 286598 106312
rect 286654 106256 286659 106312
rect 286409 106254 286659 106256
rect 284036 106252 284083 106254
rect 284017 106251 284083 106252
rect 286409 106251 286475 106254
rect 286593 106251 286659 106254
rect 289169 106314 289235 106317
rect 289353 106314 289419 106317
rect 289169 106312 289419 106314
rect 289169 106256 289174 106312
rect 289230 106256 289358 106312
rect 289414 106256 289419 106312
rect 289169 106254 289419 106256
rect 289169 106251 289235 106254
rect 289353 106251 289419 106254
rect 329557 106316 329623 106317
rect 329557 106312 329604 106316
rect 329668 106314 329674 106316
rect 361297 106314 361363 106317
rect 361438 106314 361498 106390
rect 329557 106256 329562 106312
rect 329557 106252 329604 106256
rect 329668 106254 329714 106314
rect 361297 106312 361498 106314
rect 361297 106256 361302 106312
rect 361358 106256 361498 106312
rect 361297 106254 361498 106256
rect 329668 106252 329674 106254
rect 329557 106251 329623 106252
rect 361297 106251 361363 106254
rect 583600 99636 584800 99876
rect 200389 96658 200455 96661
rect 200573 96658 200639 96661
rect 200389 96656 200639 96658
rect 200389 96600 200394 96656
rect 200450 96600 200578 96656
rect 200634 96600 200639 96656
rect 200389 96598 200639 96600
rect 200389 96595 200455 96598
rect 200573 96595 200639 96598
rect 201861 96658 201927 96661
rect 202045 96658 202111 96661
rect 201861 96656 202111 96658
rect 201861 96600 201866 96656
rect 201922 96600 202050 96656
rect 202106 96600 202111 96656
rect 201861 96598 202111 96600
rect 201861 96595 201927 96598
rect 202045 96595 202111 96598
rect 262305 96658 262371 96661
rect 262581 96658 262647 96661
rect 262305 96656 262647 96658
rect 262305 96600 262310 96656
rect 262366 96600 262586 96656
rect 262642 96600 262647 96656
rect 262305 96598 262647 96600
rect 262305 96595 262371 96598
rect 262581 96595 262647 96598
rect 318333 96658 318399 96661
rect 318517 96658 318583 96661
rect 318333 96656 318583 96658
rect 318333 96600 318338 96656
rect 318394 96600 318522 96656
rect 318578 96600 318583 96656
rect 318333 96598 318583 96600
rect 318333 96595 318399 96598
rect 318517 96595 318583 96598
rect 219525 93802 219591 93805
rect 219709 93802 219775 93805
rect 219525 93800 219775 93802
rect 219525 93744 219530 93800
rect 219586 93744 219714 93800
rect 219770 93744 219775 93800
rect 219525 93742 219775 93744
rect 219525 93739 219591 93742
rect 219709 93739 219775 93742
rect -800 93258 400 93348
rect 3509 93258 3575 93261
rect -800 93256 3575 93258
rect -800 93200 3514 93256
rect 3570 93200 3575 93256
rect -800 93198 3575 93200
rect -800 93108 400 93198
rect 3509 93195 3575 93198
rect 580441 87954 580507 87957
rect 583600 87954 584800 88044
rect 580441 87952 584800 87954
rect 580441 87896 580446 87952
rect 580502 87896 584800 87952
rect 580441 87894 584800 87896
rect 580441 87891 580507 87894
rect 583600 87804 584800 87894
rect 203149 87138 203215 87141
rect 203014 87136 203215 87138
rect 203014 87080 203154 87136
rect 203210 87080 203215 87136
rect 203014 87078 203215 87080
rect 203014 87005 203074 87078
rect 203149 87075 203215 87078
rect 203014 87000 203123 87005
rect 203014 86944 203062 87000
rect 203118 86944 203123 87000
rect 203014 86942 203123 86944
rect 203057 86939 203123 86942
rect 229277 87002 229343 87005
rect 229461 87002 229527 87005
rect 229277 87000 229527 87002
rect 229277 86944 229282 87000
rect 229338 86944 229466 87000
rect 229522 86944 229527 87000
rect 229277 86942 229527 86944
rect 229277 86939 229343 86942
rect 229461 86939 229527 86942
rect 235073 87002 235139 87005
rect 235349 87002 235415 87005
rect 235073 87000 235415 87002
rect 235073 86944 235078 87000
rect 235134 86944 235354 87000
rect 235410 86944 235415 87000
rect 235073 86942 235415 86944
rect 235073 86939 235139 86942
rect 235349 86939 235415 86942
rect 298921 87002 298987 87005
rect 299197 87002 299263 87005
rect 298921 87000 299263 87002
rect 298921 86944 298926 87000
rect 298982 86944 299202 87000
rect 299258 86944 299263 87000
rect 298921 86942 299263 86944
rect 298921 86939 298987 86942
rect 299197 86939 299263 86942
rect -800 78978 400 79068
rect 3417 78978 3483 78981
rect -800 78976 3483 78978
rect -800 78920 3422 78976
rect 3478 78920 3483 78976
rect -800 78918 3483 78920
rect -800 78828 400 78918
rect 3417 78915 3483 78918
rect 258165 77210 258231 77213
rect 258349 77210 258415 77213
rect 258165 77208 258415 77210
rect 258165 77152 258170 77208
rect 258226 77152 258354 77208
rect 258410 77152 258415 77208
rect 258165 77150 258415 77152
rect 258165 77147 258231 77150
rect 258349 77147 258415 77150
rect 580349 76258 580415 76261
rect 583600 76258 584800 76348
rect 580349 76256 584800 76258
rect 580349 76200 580354 76256
rect 580410 76200 584800 76256
rect 580349 76198 584800 76200
rect 580349 76195 580415 76198
rect 583600 76108 584800 76198
rect 260925 67690 260991 67693
rect 261109 67690 261175 67693
rect 260925 67688 261175 67690
rect 260925 67632 260930 67688
rect 260986 67632 261114 67688
rect 261170 67632 261175 67688
rect 260925 67630 261175 67632
rect 260925 67627 260991 67630
rect 261109 67627 261175 67630
rect 316861 67554 316927 67557
rect 317045 67554 317111 67557
rect 318333 67554 318399 67557
rect 316861 67552 317111 67554
rect 316861 67496 316866 67552
rect 316922 67496 317050 67552
rect 317106 67496 317111 67552
rect 316861 67494 317111 67496
rect 316861 67491 316927 67494
rect 317045 67491 317111 67494
rect 318198 67552 318399 67554
rect 318198 67496 318338 67552
rect 318394 67496 318399 67552
rect 318198 67494 318399 67496
rect 318198 67418 318258 67494
rect 318333 67491 318399 67494
rect 318517 67418 318583 67421
rect 318198 67416 318583 67418
rect 318198 67360 318522 67416
rect 318578 67360 318583 67416
rect 318198 67358 318583 67360
rect 318517 67355 318583 67358
rect 194961 66194 195027 66197
rect 195094 66194 195100 66196
rect 194961 66192 195100 66194
rect 194961 66136 194966 66192
rect 195022 66136 195100 66192
rect 194961 66134 195100 66136
rect 194961 66131 195027 66134
rect 195094 66132 195100 66134
rect 195164 66132 195170 66196
rect 191097 65106 191163 65109
rect 343357 65106 343423 65109
rect 191054 65104 191163 65106
rect 191054 65048 191102 65104
rect 191158 65048 191163 65104
rect 191054 65043 191163 65048
rect 343222 65104 343423 65106
rect 343222 65048 343362 65104
rect 343418 65048 343423 65104
rect 343222 65046 343423 65048
rect 191054 64973 191114 65043
rect 343222 64973 343282 65046
rect 343357 65043 343423 65046
rect 191005 64968 191114 64973
rect 191005 64912 191010 64968
rect 191066 64912 191114 64968
rect 191005 64910 191114 64912
rect 343173 64968 343282 64973
rect 343173 64912 343178 64968
rect 343234 64912 343282 64968
rect 343173 64910 343282 64912
rect 191005 64907 191071 64910
rect 343173 64907 343239 64910
rect 749 64834 815 64837
rect 359038 64834 359044 64836
rect 749 64832 359044 64834
rect 749 64776 754 64832
rect 810 64776 359044 64832
rect 749 64774 359044 64776
rect 749 64771 815 64774
rect 359038 64772 359044 64774
rect 359108 64772 359114 64836
rect -800 64562 400 64652
rect 749 64562 815 64565
rect -800 64560 815 64562
rect -800 64504 754 64560
rect 810 64504 815 64560
rect -800 64502 815 64504
rect -800 64412 400 64502
rect 749 64499 815 64502
rect 580257 64562 580323 64565
rect 583600 64562 584800 64652
rect 580257 64560 584800 64562
rect 580257 64504 580262 64560
rect 580318 64504 584800 64560
rect 580257 64502 584800 64504
rect 580257 64499 580323 64502
rect 583600 64412 584800 64502
rect 178033 63474 178099 63477
rect 178309 63474 178375 63477
rect 178033 63472 178375 63474
rect 178033 63416 178038 63472
rect 178094 63416 178314 63472
rect 178370 63416 178375 63472
rect 178033 63414 178375 63416
rect 178033 63411 178099 63414
rect 178309 63411 178375 63414
rect 341701 62114 341767 62117
rect 341885 62114 341951 62117
rect 341701 62112 341951 62114
rect 341701 62056 341706 62112
rect 341762 62056 341890 62112
rect 341946 62056 341951 62112
rect 341701 62054 341951 62056
rect 341701 62051 341767 62054
rect 341885 62051 341951 62054
rect 211889 58170 211955 58173
rect 211846 58168 211955 58170
rect 211846 58112 211894 58168
rect 211950 58112 211955 58168
rect 211846 58107 211955 58112
rect 194869 57898 194935 57901
rect 195094 57898 195100 57900
rect 194869 57896 195100 57898
rect 194869 57840 194874 57896
rect 194930 57840 195100 57896
rect 194869 57838 195100 57840
rect 194869 57835 194935 57838
rect 195094 57836 195100 57838
rect 195164 57836 195170 57900
rect 211846 57898 211906 58107
rect 316861 58034 316927 58037
rect 316861 58032 317338 58034
rect 316861 57976 316866 58032
rect 316922 57976 317338 58032
rect 316861 57974 317338 57976
rect 316861 57971 316927 57974
rect 211981 57898 212047 57901
rect 211846 57896 212047 57898
rect 211846 57840 211986 57896
rect 212042 57840 212047 57896
rect 211846 57838 212047 57840
rect 211981 57835 212047 57838
rect 317045 57898 317111 57901
rect 317278 57898 317338 57974
rect 317045 57896 317338 57898
rect 317045 57840 317050 57896
rect 317106 57840 317338 57896
rect 317045 57838 317338 57840
rect 317045 57835 317111 57838
rect 191097 54090 191163 54093
rect 191097 54088 191298 54090
rect 191097 54032 191102 54088
rect 191158 54032 191298 54088
rect 191097 54030 191298 54032
rect 191097 54027 191163 54030
rect 191097 53954 191163 53957
rect 191238 53954 191298 54030
rect 191097 53952 191298 53954
rect 191097 53896 191102 53952
rect 191158 53896 191298 53952
rect 191097 53894 191298 53896
rect 191097 53891 191163 53894
rect 190913 53818 190979 53821
rect 191097 53818 191163 53821
rect 190913 53816 191163 53818
rect 190913 53760 190918 53816
rect 190974 53760 191102 53816
rect 191158 53760 191163 53816
rect 190913 53758 191163 53760
rect 190913 53755 190979 53758
rect 191097 53755 191163 53758
rect 583600 52716 584800 52956
rect 329414 51172 329420 51236
rect 329484 51234 329490 51236
rect 329557 51234 329623 51237
rect 329484 51232 329623 51234
rect 329484 51176 329562 51232
rect 329618 51176 329623 51232
rect 329484 51174 329623 51176
rect 329484 51172 329490 51174
rect 329557 51171 329623 51174
rect -800 50146 400 50236
rect 2773 50146 2839 50149
rect -800 50144 2839 50146
rect -800 50088 2778 50144
rect 2834 50088 2839 50144
rect -800 50086 2839 50088
rect -800 49996 400 50086
rect 2773 50083 2839 50086
rect 236361 48514 236427 48517
rect 236134 48512 236427 48514
rect 236134 48456 236366 48512
rect 236422 48456 236427 48512
rect 236134 48454 236427 48456
rect 236134 48378 236194 48454
rect 236361 48451 236427 48454
rect 236269 48378 236335 48381
rect 236134 48376 236335 48378
rect 236134 48320 236274 48376
rect 236330 48320 236335 48376
rect 236134 48318 236335 48320
rect 236269 48315 236335 48318
rect 327901 48378 327967 48381
rect 328085 48378 328151 48381
rect 329465 48380 329531 48381
rect 327901 48376 328151 48378
rect 327901 48320 327906 48376
rect 327962 48320 328090 48376
rect 328146 48320 328151 48376
rect 327901 48318 328151 48320
rect 327901 48315 327967 48318
rect 328085 48315 328151 48318
rect 329414 48316 329420 48380
rect 329484 48378 329531 48380
rect 329484 48376 329576 48378
rect 329526 48320 329576 48376
rect 329484 48318 329576 48320
rect 329484 48316 329531 48318
rect 329465 48315 329531 48316
rect 318425 46882 318491 46885
rect 318425 46880 318626 46882
rect 318425 46824 318430 46880
rect 318486 46824 318626 46880
rect 318425 46822 318626 46824
rect 318425 46819 318491 46822
rect 318333 46746 318399 46749
rect 318566 46746 318626 46822
rect 318333 46744 318626 46746
rect 318333 46688 318338 46744
rect 318394 46688 318626 46744
rect 318333 46686 318626 46688
rect 318333 46683 318399 46686
rect 234981 41442 235047 41445
rect 235349 41442 235415 41445
rect 234981 41440 235415 41442
rect 234981 41384 234986 41440
rect 235042 41384 235354 41440
rect 235410 41384 235415 41440
rect 234981 41382 235415 41384
rect 234981 41379 235047 41382
rect 235349 41379 235415 41382
rect 576853 41170 576919 41173
rect 583385 41170 583451 41173
rect 576853 41168 583451 41170
rect 576853 41112 576858 41168
rect 576914 41112 583390 41168
rect 583446 41112 583451 41168
rect 576853 41110 583451 41112
rect 576853 41107 576919 41110
rect 583385 41107 583451 41110
rect 583385 41034 583451 41037
rect 583600 41034 584800 41124
rect 583385 41032 584800 41034
rect 583385 40976 583390 41032
rect 583446 40976 584800 41032
rect 583385 40974 584800 40976
rect 583385 40971 583451 40974
rect 583600 40884 584800 40974
rect 327022 40564 327028 40628
rect 327092 40626 327098 40628
rect 327092 40566 336658 40626
rect 327092 40564 327098 40566
rect 336598 40492 336658 40566
rect 336774 40564 336780 40628
rect 336844 40626 336850 40628
rect 338205 40626 338271 40629
rect 336844 40624 338271 40626
rect 336844 40568 338210 40624
rect 338266 40568 338271 40624
rect 336844 40566 338271 40568
rect 336844 40564 336850 40566
rect 338205 40563 338271 40566
rect 307702 40428 307708 40492
rect 307772 40490 307778 40492
rect 307772 40430 317338 40490
rect 307772 40428 307778 40430
rect 173382 40292 173388 40356
rect 173452 40354 173458 40356
rect 289905 40354 289971 40357
rect 317278 40354 317338 40430
rect 321326 40430 322306 40490
rect 321326 40354 321386 40430
rect 173452 40294 176762 40354
rect 173452 40292 173458 40294
rect 176702 40218 176762 40294
rect 232270 40294 264346 40354
rect 220721 40218 220787 40221
rect 176702 40158 191850 40218
rect 191790 40082 191850 40158
rect 220721 40216 222026 40218
rect 220721 40160 220726 40216
rect 220782 40160 222026 40216
rect 220721 40158 222026 40160
rect 220721 40155 220787 40158
rect 221966 40116 222026 40158
rect 201861 40082 201927 40085
rect 212441 40082 212507 40085
rect 191790 40022 192034 40082
rect 191974 39946 192034 40022
rect 201861 40080 212507 40082
rect 201861 40024 201866 40080
rect 201922 40024 212446 40080
rect 212502 40024 212507 40080
rect 221966 40082 222394 40116
rect 232270 40082 232330 40294
rect 264286 40218 264346 40294
rect 289905 40352 304274 40354
rect 289905 40296 289910 40352
rect 289966 40296 304274 40352
rect 289905 40294 304274 40296
rect 317278 40294 321386 40354
rect 289905 40291 289971 40294
rect 270493 40218 270559 40221
rect 264286 40216 270559 40218
rect 264286 40160 270498 40216
rect 270554 40160 270559 40216
rect 264286 40158 270559 40160
rect 270493 40155 270559 40158
rect 275737 40218 275803 40221
rect 289813 40218 289879 40221
rect 275737 40216 289879 40218
rect 275737 40160 275742 40216
rect 275798 40160 289818 40216
rect 289874 40160 289879 40216
rect 275737 40158 289879 40160
rect 304214 40218 304274 40294
rect 307702 40218 307708 40220
rect 304214 40158 307708 40218
rect 275737 40155 275803 40158
rect 289813 40155 289879 40158
rect 307702 40156 307708 40158
rect 307772 40156 307778 40220
rect 322246 40218 322306 40430
rect 336590 40428 336596 40492
rect 336660 40428 336666 40492
rect 384982 40428 384988 40492
rect 385052 40490 385058 40492
rect 394601 40490 394667 40493
rect 385052 40488 394667 40490
rect 385052 40432 394606 40488
rect 394662 40432 394667 40488
rect 385052 40430 394667 40432
rect 385052 40428 385058 40430
rect 394601 40427 394667 40430
rect 327022 40292 327028 40356
rect 327092 40292 327098 40356
rect 367093 40354 367159 40357
rect 360150 40352 367159 40354
rect 360150 40296 367098 40352
rect 367154 40296 367159 40352
rect 360150 40294 367159 40296
rect 327030 40218 327090 40292
rect 322246 40158 327090 40218
rect 338205 40218 338271 40221
rect 338205 40216 347882 40218
rect 338205 40160 338210 40216
rect 338266 40160 347882 40216
rect 338205 40158 347882 40160
rect 338205 40155 338271 40158
rect 221966 40056 232330 40082
rect 201861 40022 212507 40024
rect 222334 40022 232330 40056
rect 347822 40082 347882 40158
rect 360150 40082 360210 40294
rect 367093 40291 367159 40294
rect 405641 40354 405707 40357
rect 405641 40352 412650 40354
rect 405641 40296 405646 40352
rect 405702 40296 412650 40352
rect 405641 40294 412650 40296
rect 405641 40291 405707 40294
rect 379605 40218 379671 40221
rect 384982 40218 384988 40220
rect 379605 40216 384988 40218
rect 379605 40160 379610 40216
rect 379666 40160 384988 40216
rect 379605 40158 384988 40160
rect 379605 40155 379671 40158
rect 384982 40156 384988 40158
rect 385052 40156 385058 40220
rect 398741 40218 398807 40221
rect 396030 40216 398807 40218
rect 396030 40160 398746 40216
rect 398802 40160 398807 40216
rect 396030 40158 398807 40160
rect 412590 40218 412650 40294
rect 422342 40294 431970 40354
rect 412590 40158 422218 40218
rect 347822 40022 360210 40082
rect 369945 40082 370011 40085
rect 379421 40082 379487 40085
rect 369945 40080 379487 40082
rect 369945 40024 369950 40080
rect 370006 40024 379426 40080
rect 379482 40024 379487 40080
rect 369945 40022 379487 40024
rect 201861 40019 201927 40022
rect 212441 40019 212507 40022
rect 369945 40019 370011 40022
rect 379421 40019 379487 40022
rect 394601 40082 394667 40085
rect 396030 40082 396090 40158
rect 398741 40155 398807 40158
rect 394601 40080 396090 40082
rect 394601 40024 394606 40080
rect 394662 40024 396090 40080
rect 394601 40022 396090 40024
rect 422158 40082 422218 40158
rect 422342 40082 422402 40294
rect 431910 40218 431970 40294
rect 441662 40294 451290 40354
rect 431910 40158 441538 40218
rect 422158 40022 422402 40082
rect 441478 40082 441538 40158
rect 441662 40082 441722 40294
rect 451230 40218 451290 40294
rect 460982 40294 470610 40354
rect 451230 40158 460858 40218
rect 441478 40022 441722 40082
rect 460798 40082 460858 40158
rect 460982 40082 461042 40294
rect 470550 40218 470610 40294
rect 480302 40294 489930 40354
rect 470550 40158 480178 40218
rect 460798 40022 461042 40082
rect 480118 40082 480178 40158
rect 480302 40082 480362 40294
rect 489870 40218 489930 40294
rect 499622 40294 509250 40354
rect 489870 40158 499498 40218
rect 480118 40022 480362 40082
rect 499438 40082 499498 40158
rect 499622 40082 499682 40294
rect 509190 40218 509250 40294
rect 518942 40294 528570 40354
rect 509190 40158 518818 40218
rect 499438 40022 499682 40082
rect 518758 40082 518818 40158
rect 518942 40082 519002 40294
rect 528510 40218 528570 40294
rect 538262 40294 547890 40354
rect 528510 40158 538138 40218
rect 518758 40022 519002 40082
rect 538078 40082 538138 40158
rect 538262 40082 538322 40294
rect 547830 40218 547890 40294
rect 557582 40294 567210 40354
rect 547830 40158 557458 40218
rect 538078 40022 538322 40082
rect 557398 40082 557458 40158
rect 557582 40082 557642 40294
rect 567150 40218 567210 40294
rect 567150 40158 576778 40218
rect 557398 40022 557642 40082
rect 576718 40082 576778 40158
rect 576853 40082 576919 40085
rect 576718 40080 576919 40082
rect 576718 40024 576858 40080
rect 576914 40024 576919 40080
rect 576718 40022 576919 40024
rect 394601 40019 394667 40022
rect 576853 40019 576919 40022
rect 201493 39946 201559 39949
rect 191974 39944 201559 39946
rect 191974 39888 201498 39944
rect 201554 39888 201559 39944
rect 191974 39886 201559 39888
rect 201493 39883 201559 39886
rect 195145 37362 195211 37365
rect 195102 37360 195211 37362
rect 195102 37304 195150 37360
rect 195206 37304 195211 37360
rect 195102 37299 195211 37304
rect 194869 37226 194935 37229
rect 195102 37226 195162 37299
rect 194869 37224 195162 37226
rect 194869 37168 194874 37224
rect 194930 37168 195162 37224
rect 194869 37166 195162 37168
rect 194869 37163 194935 37166
rect -800 35866 400 35956
rect 2773 35866 2839 35869
rect -800 35864 2839 35866
rect -800 35808 2778 35864
rect 2834 35808 2839 35864
rect -800 35806 2839 35808
rect -800 35716 400 35806
rect 2773 35803 2839 35806
rect 580257 29338 580323 29341
rect 583600 29338 584800 29428
rect 580257 29336 584800 29338
rect 580257 29280 580262 29336
rect 580318 29280 584800 29336
rect 580257 29278 584800 29280
rect 580257 29275 580323 29278
rect 268745 29202 268811 29205
rect 268745 29200 268946 29202
rect 268745 29144 268750 29200
rect 268806 29144 268946 29200
rect 583600 29188 584800 29278
rect 268745 29142 268946 29144
rect 268745 29139 268811 29142
rect 268745 29066 268811 29069
rect 268886 29066 268946 29142
rect 268745 29064 268946 29066
rect 268745 29008 268750 29064
rect 268806 29008 268946 29064
rect 268745 29006 268946 29008
rect 268745 29003 268811 29006
rect 473 21994 539 21997
rect 362902 21994 362908 21996
rect 473 21992 362908 21994
rect 473 21936 478 21992
rect 534 21936 362908 21992
rect 473 21934 362908 21936
rect 473 21931 539 21934
rect 362902 21932 362908 21934
rect 362972 21932 362978 21996
rect -800 21450 400 21540
rect 473 21450 539 21453
rect -800 21448 539 21450
rect -800 21392 478 21448
rect 534 21392 539 21448
rect -800 21390 539 21392
rect -800 21300 400 21390
rect 473 21387 539 21390
rect 289261 18048 289327 18053
rect 289261 17992 289266 18048
rect 289322 17992 289327 18048
rect 289261 17987 289327 17992
rect 289264 17917 289324 17987
rect 289261 17912 289327 17917
rect 289261 17856 289266 17912
rect 289322 17856 289327 17912
rect 289261 17851 289327 17856
rect 579613 17642 579679 17645
rect 583600 17642 584800 17732
rect 579613 17640 584800 17642
rect 579613 17584 579618 17640
rect 579674 17584 584800 17640
rect 579613 17582 584800 17584
rect 579613 17579 579679 17582
rect 583600 17492 584800 17582
rect 2957 10298 3023 10301
rect 361614 10298 361620 10300
rect 2957 10296 361620 10298
rect 2957 10240 2962 10296
rect 3018 10240 361620 10296
rect 2957 10238 361620 10240
rect 2957 10235 3023 10238
rect 361614 10236 361620 10238
rect 361684 10236 361690 10300
rect 362493 9618 362559 9621
rect 362493 9616 362602 9618
rect 362493 9560 362498 9616
rect 362554 9560 362602 9616
rect 362493 9555 362602 9560
rect 362542 9482 362602 9555
rect 363597 9482 363663 9485
rect 362542 9480 363663 9482
rect 362542 9424 363602 9480
rect 363658 9424 363663 9480
rect 362542 9422 363663 9424
rect 363597 9419 363663 9422
rect 331029 8938 331095 8941
rect 466821 8938 466887 8941
rect 331029 8936 466887 8938
rect 331029 8880 331034 8936
rect 331090 8880 466826 8936
rect 466882 8880 466887 8936
rect 331029 8878 466887 8880
rect 331029 8875 331095 8878
rect 466821 8875 466887 8878
rect 52821 7578 52887 7581
rect 187877 7578 187943 7581
rect 52821 7576 187943 7578
rect 52821 7520 52826 7576
rect 52882 7520 187882 7576
rect 187938 7520 187943 7576
rect 52821 7518 187943 7520
rect 52821 7515 52887 7518
rect 187877 7515 187943 7518
rect 369577 7578 369643 7581
rect 580993 7578 581059 7581
rect 369577 7576 581059 7578
rect 369577 7520 369582 7576
rect 369638 7520 580998 7576
rect 581054 7520 581059 7576
rect 369577 7518 581059 7520
rect 369577 7515 369643 7518
rect 580993 7515 581059 7518
rect -800 7170 400 7260
rect 2957 7170 3023 7173
rect -800 7168 3023 7170
rect -800 7112 2962 7168
rect 3018 7112 3023 7168
rect -800 7110 3023 7112
rect -800 7020 400 7110
rect 2957 7107 3023 7110
rect 21909 6218 21975 6221
rect 176837 6218 176903 6221
rect 21909 6216 176903 6218
rect 21909 6160 21914 6216
rect 21970 6160 176842 6216
rect 176898 6160 176903 6216
rect 21909 6158 176903 6160
rect 21909 6155 21975 6158
rect 176837 6155 176903 6158
rect 333789 6218 333855 6221
rect 476297 6218 476363 6221
rect 333789 6216 476363 6218
rect 333789 6160 333794 6216
rect 333850 6160 476302 6216
rect 476358 6160 476363 6216
rect 333789 6158 476363 6160
rect 333789 6155 333855 6158
rect 476297 6155 476363 6158
rect 583600 5796 584800 6036
rect 565 4858 631 4861
rect 170029 4858 170095 4861
rect 565 4856 170095 4858
rect 565 4800 570 4856
rect 626 4800 170034 4856
rect 170090 4800 170095 4856
rect 565 4798 170095 4800
rect 565 4795 631 4798
rect 170029 4795 170095 4798
rect 297909 4858 297975 4861
rect 372797 4858 372863 4861
rect 297909 4856 372863 4858
rect 297909 4800 297914 4856
rect 297970 4800 372802 4856
rect 372858 4800 372863 4856
rect 297909 4798 372863 4800
rect 297909 4795 297975 4798
rect 372797 4795 372863 4798
rect 306373 4178 306439 4181
rect 311065 4178 311131 4181
rect 306373 4176 311131 4178
rect 306373 4120 306378 4176
rect 306434 4120 311070 4176
rect 311126 4120 311131 4176
rect 306373 4118 311131 4120
rect 306373 4115 306439 4118
rect 311065 4115 311131 4118
rect 5257 3362 5323 3365
rect 171133 3362 171199 3365
rect 5257 3360 171199 3362
rect 5257 3304 5262 3360
rect 5318 3304 171138 3360
rect 171194 3304 171199 3360
rect 5257 3302 171199 3304
rect 5257 3299 5323 3302
rect 171133 3299 171199 3302
rect 284201 3362 284267 3365
rect 332409 3362 332475 3365
rect 284201 3360 332475 3362
rect 284201 3304 284206 3360
rect 284262 3304 332414 3360
rect 332470 3304 332475 3360
rect 284201 3302 332475 3304
rect 284201 3299 284267 3302
rect 332409 3299 332475 3302
rect 277209 3090 277275 3093
rect 280429 3090 280495 3093
rect 277209 3088 280495 3090
rect 277209 3032 277214 3088
rect 277270 3032 280434 3088
rect 280490 3032 280495 3088
rect 277209 3030 280495 3032
rect 277209 3027 277275 3030
rect 280429 3027 280495 3030
<< via3 >>
rect 267412 645824 267476 645828
rect 267412 645768 267462 645824
rect 267462 645768 267476 645824
rect 267412 645764 267476 645768
rect 267412 640188 267476 640252
rect 359780 522956 359844 523020
rect 359596 522820 359660 522884
rect 359412 522684 359476 522748
rect 366220 520236 366284 520300
rect 309364 519420 309428 519484
rect 313228 519420 313292 519484
rect 173388 519284 173452 519348
rect 193076 519344 193140 519348
rect 193076 519288 193126 519344
rect 193126 519288 193140 519344
rect 193076 519284 193140 519288
rect 195100 519344 195164 519348
rect 195100 519288 195114 519344
rect 195114 519288 195164 519344
rect 195100 519284 195164 519288
rect 198412 519344 198476 519348
rect 198412 519288 198426 519344
rect 198426 519288 198476 519344
rect 198412 519284 198476 519288
rect 199884 519344 199948 519348
rect 199884 519288 199934 519344
rect 199934 519288 199948 519344
rect 199884 519284 199948 519288
rect 205220 519344 205284 519348
rect 205220 519288 205234 519344
rect 205234 519288 205284 519344
rect 205220 519284 205284 519288
rect 210372 519344 210436 519348
rect 210372 519288 210386 519344
rect 210386 519288 210436 519344
rect 210372 519284 210436 519288
rect 234292 519284 234356 519348
rect 236500 519284 236564 519348
rect 280108 519284 280172 519348
rect 284892 519284 284956 519348
rect 312676 519284 312740 519348
rect 359044 519344 359108 519348
rect 359044 519288 359058 519344
rect 359058 519288 359108 519344
rect 359044 519284 359108 519288
rect 361620 519284 361684 519348
rect 362908 519284 362972 519348
rect 234476 519148 234540 519212
rect 236684 519148 236748 519212
rect 241468 519148 241532 519212
rect 246436 519148 246500 519212
rect 263180 519148 263244 519212
rect 265572 519148 265636 519212
rect 294460 519148 294524 519212
rect 299244 519148 299308 519212
rect 313228 519148 313292 519212
rect 322796 519148 322860 519212
rect 236868 519012 236932 519076
rect 263364 519012 263428 519076
rect 241468 518740 241532 518804
rect 210372 518604 210436 518668
rect 234476 518604 234540 518668
rect 182220 518468 182284 518532
rect 176516 517924 176580 517988
rect 176700 517924 176764 517988
rect 182220 517924 182284 517988
rect 199884 518468 199948 518532
rect 236868 518604 236932 518668
rect 243860 518604 243924 518668
rect 244228 518604 244292 518668
rect 253612 518876 253676 518940
rect 246436 518740 246500 518804
rect 263364 518740 263428 518804
rect 253612 518604 253676 518668
rect 253796 518604 253860 518668
rect 263180 518604 263244 518668
rect 272932 519012 272996 519076
rect 280108 519012 280172 519076
rect 294276 518876 294340 518940
rect 298876 518876 298940 518940
rect 272932 518604 272996 518668
rect 273116 518604 273180 518668
rect 283052 518604 283116 518668
rect 302740 518876 302804 518940
rect 312676 518876 312740 518940
rect 284892 518604 284956 518668
rect 294276 518604 294340 518668
rect 294644 518604 294708 518668
rect 298692 518604 298756 518668
rect 298876 518604 298940 518668
rect 301820 518604 301884 518668
rect 302004 518604 302068 518668
rect 309180 518604 309244 518668
rect 321692 518740 321756 518804
rect 335308 518740 335372 518804
rect 321508 518604 321572 518668
rect 322796 518604 322860 518668
rect 336412 518740 336476 518804
rect 367324 518876 367388 518940
rect 198412 518332 198476 518396
rect 234292 518332 234356 518396
rect 234660 518332 234724 518396
rect 236316 518332 236380 518396
rect 236500 518332 236564 518396
rect 367324 518332 367388 518396
rect 195100 518196 195164 518260
rect 294460 518196 294524 518260
rect 193076 518060 193140 518124
rect 234660 518060 234724 518124
rect 236316 518060 236380 518124
rect 299060 518196 299124 518260
rect 299244 518196 299308 518260
rect 299244 518060 299308 518124
rect 367140 518060 367204 518124
rect 367324 518060 367388 518124
rect 196020 517924 196084 517988
rect 210372 517924 210436 517988
rect 219204 517924 219268 517988
rect 234476 517924 234540 517988
rect 236684 517924 236748 517988
rect 243308 517924 243372 517988
rect 243676 517924 243740 517988
rect 244228 517924 244292 517988
rect 244412 517924 244476 517988
rect 253796 517924 253860 517988
rect 254164 517924 254228 517988
rect 264468 517924 264532 517988
rect 265572 517924 265636 517988
rect 273116 517924 273180 517988
rect 273484 517924 273548 517988
rect 282868 517924 282932 517988
rect 283052 517924 283116 517988
rect 294644 517924 294708 517988
rect 298876 517924 298940 517988
rect 302004 517924 302068 517988
rect 302188 517924 302252 517988
rect 195836 517788 195900 517852
rect 205220 517788 205284 517852
rect 298508 517788 298572 517852
rect 298876 517788 298940 517852
rect 367324 517788 367388 517852
rect 367324 517652 367388 517716
rect 368980 517652 369044 517716
rect 367140 486372 367204 486436
rect 384988 486236 385052 486300
rect 359780 485828 359844 485892
rect 367140 486100 367204 486164
rect 384988 485964 385052 486028
rect 368980 310796 369044 310860
rect 359596 298148 359660 298212
rect 359412 251228 359476 251292
rect 275876 217968 275940 217972
rect 275876 217912 275926 217968
rect 275926 217912 275940 217968
rect 275876 217908 275940 217912
rect 275876 217696 275940 217700
rect 275876 217640 275926 217696
rect 275926 217640 275940 217696
rect 275876 217636 275940 217640
rect 366220 204580 366284 204644
rect 277164 162692 277228 162756
rect 277164 153232 277228 153236
rect 277164 153176 277178 153232
rect 277178 153176 277228 153232
rect 277164 153172 277228 153176
rect 318564 147792 318628 147796
rect 318564 147736 318578 147792
rect 318578 147736 318628 147792
rect 318564 147732 318628 147736
rect 329604 147792 329668 147796
rect 329604 147736 329618 147792
rect 329618 147736 329668 147792
rect 329604 147732 329668 147736
rect 329604 144936 329668 144940
rect 329604 144880 329618 144936
rect 329618 144880 329668 144936
rect 329604 144876 329668 144880
rect 194916 143576 194980 143580
rect 194916 143520 194966 143576
rect 194966 143520 194980 143576
rect 194916 143516 194980 143520
rect 318564 143576 318628 143580
rect 318564 143520 318578 143576
rect 318578 143520 318628 143576
rect 318564 143516 318628 143520
rect 194916 142216 194980 142220
rect 194916 142160 194966 142216
rect 194966 142160 194980 142216
rect 194916 142156 194980 142160
rect 329604 128480 329668 128484
rect 329604 128424 329618 128480
rect 329618 128424 329668 128480
rect 329604 128420 329668 128424
rect 329604 125624 329668 125628
rect 329604 125568 329618 125624
rect 329618 125568 329668 125624
rect 329604 125564 329668 125568
rect 283972 123932 284036 123996
rect 329604 109168 329668 109172
rect 329604 109112 329618 109168
rect 329618 109112 329668 109168
rect 329604 109108 329668 109112
rect 283972 106312 284036 106316
rect 283972 106256 284022 106312
rect 284022 106256 284036 106312
rect 283972 106252 284036 106256
rect 329604 106312 329668 106316
rect 329604 106256 329618 106312
rect 329618 106256 329668 106312
rect 329604 106252 329668 106256
rect 195100 66132 195164 66196
rect 359044 64772 359108 64836
rect 195100 57836 195164 57900
rect 329420 51172 329484 51236
rect 329420 48376 329484 48380
rect 329420 48320 329470 48376
rect 329470 48320 329484 48376
rect 329420 48316 329484 48320
rect 327028 40564 327092 40628
rect 336780 40564 336844 40628
rect 307708 40428 307772 40492
rect 173388 40292 173452 40356
rect 307708 40156 307772 40220
rect 336596 40428 336660 40492
rect 384988 40428 385052 40492
rect 327028 40292 327092 40356
rect 384988 40156 385052 40220
rect 362908 21932 362972 21996
rect 361620 10236 361684 10300
<< metal4 >>
rect -8436 711278 -7836 711300
rect -8436 711042 -8254 711278
rect -8018 711042 -7836 711278
rect -8436 710958 -7836 711042
rect -8436 710722 -8254 710958
rect -8018 710722 -7836 710958
rect -8436 679254 -7836 710722
rect -8436 679018 -8254 679254
rect -8018 679018 -7836 679254
rect -8436 678934 -7836 679018
rect -8436 678698 -8254 678934
rect -8018 678698 -7836 678934
rect -8436 643254 -7836 678698
rect -8436 643018 -8254 643254
rect -8018 643018 -7836 643254
rect -8436 642934 -7836 643018
rect -8436 642698 -8254 642934
rect -8018 642698 -7836 642934
rect -8436 607254 -7836 642698
rect -8436 607018 -8254 607254
rect -8018 607018 -7836 607254
rect -8436 606934 -7836 607018
rect -8436 606698 -8254 606934
rect -8018 606698 -7836 606934
rect -8436 571254 -7836 606698
rect -8436 571018 -8254 571254
rect -8018 571018 -7836 571254
rect -8436 570934 -7836 571018
rect -8436 570698 -8254 570934
rect -8018 570698 -7836 570934
rect -8436 535254 -7836 570698
rect -8436 535018 -8254 535254
rect -8018 535018 -7836 535254
rect -8436 534934 -7836 535018
rect -8436 534698 -8254 534934
rect -8018 534698 -7836 534934
rect -8436 499254 -7836 534698
rect -8436 499018 -8254 499254
rect -8018 499018 -7836 499254
rect -8436 498934 -7836 499018
rect -8436 498698 -8254 498934
rect -8018 498698 -7836 498934
rect -8436 463254 -7836 498698
rect -8436 463018 -8254 463254
rect -8018 463018 -7836 463254
rect -8436 462934 -7836 463018
rect -8436 462698 -8254 462934
rect -8018 462698 -7836 462934
rect -8436 427254 -7836 462698
rect -8436 427018 -8254 427254
rect -8018 427018 -7836 427254
rect -8436 426934 -7836 427018
rect -8436 426698 -8254 426934
rect -8018 426698 -7836 426934
rect -8436 391254 -7836 426698
rect -8436 391018 -8254 391254
rect -8018 391018 -7836 391254
rect -8436 390934 -7836 391018
rect -8436 390698 -8254 390934
rect -8018 390698 -7836 390934
rect -8436 355254 -7836 390698
rect -8436 355018 -8254 355254
rect -8018 355018 -7836 355254
rect -8436 354934 -7836 355018
rect -8436 354698 -8254 354934
rect -8018 354698 -7836 354934
rect -8436 319254 -7836 354698
rect -8436 319018 -8254 319254
rect -8018 319018 -7836 319254
rect -8436 318934 -7836 319018
rect -8436 318698 -8254 318934
rect -8018 318698 -7836 318934
rect -8436 283254 -7836 318698
rect -8436 283018 -8254 283254
rect -8018 283018 -7836 283254
rect -8436 282934 -7836 283018
rect -8436 282698 -8254 282934
rect -8018 282698 -7836 282934
rect -8436 247254 -7836 282698
rect -8436 247018 -8254 247254
rect -8018 247018 -7836 247254
rect -8436 246934 -7836 247018
rect -8436 246698 -8254 246934
rect -8018 246698 -7836 246934
rect -8436 211254 -7836 246698
rect -8436 211018 -8254 211254
rect -8018 211018 -7836 211254
rect -8436 210934 -7836 211018
rect -8436 210698 -8254 210934
rect -8018 210698 -7836 210934
rect -8436 175254 -7836 210698
rect -8436 175018 -8254 175254
rect -8018 175018 -7836 175254
rect -8436 174934 -7836 175018
rect -8436 174698 -8254 174934
rect -8018 174698 -7836 174934
rect -8436 139254 -7836 174698
rect -8436 139018 -8254 139254
rect -8018 139018 -7836 139254
rect -8436 138934 -7836 139018
rect -8436 138698 -8254 138934
rect -8018 138698 -7836 138934
rect -8436 103254 -7836 138698
rect -8436 103018 -8254 103254
rect -8018 103018 -7836 103254
rect -8436 102934 -7836 103018
rect -8436 102698 -8254 102934
rect -8018 102698 -7836 102934
rect -8436 67254 -7836 102698
rect -8436 67018 -8254 67254
rect -8018 67018 -7836 67254
rect -8436 66934 -7836 67018
rect -8436 66698 -8254 66934
rect -8018 66698 -7836 66934
rect -8436 31254 -7836 66698
rect -8436 31018 -8254 31254
rect -8018 31018 -7836 31254
rect -8436 30934 -7836 31018
rect -8436 30698 -8254 30934
rect -8018 30698 -7836 30934
rect -8436 -6786 -7836 30698
rect -7516 710358 -6916 710380
rect -7516 710122 -7334 710358
rect -7098 710122 -6916 710358
rect -7516 710038 -6916 710122
rect -7516 709802 -7334 710038
rect -7098 709802 -6916 710038
rect -7516 697254 -6916 709802
rect 11604 710358 12204 711300
rect 11604 710122 11786 710358
rect 12022 710122 12204 710358
rect 11604 710038 12204 710122
rect 11604 709802 11786 710038
rect 12022 709802 12204 710038
rect -7516 697018 -7334 697254
rect -7098 697018 -6916 697254
rect -7516 696934 -6916 697018
rect -7516 696698 -7334 696934
rect -7098 696698 -6916 696934
rect -7516 661254 -6916 696698
rect -7516 661018 -7334 661254
rect -7098 661018 -6916 661254
rect -7516 660934 -6916 661018
rect -7516 660698 -7334 660934
rect -7098 660698 -6916 660934
rect -7516 625254 -6916 660698
rect -7516 625018 -7334 625254
rect -7098 625018 -6916 625254
rect -7516 624934 -6916 625018
rect -7516 624698 -7334 624934
rect -7098 624698 -6916 624934
rect -7516 589254 -6916 624698
rect -7516 589018 -7334 589254
rect -7098 589018 -6916 589254
rect -7516 588934 -6916 589018
rect -7516 588698 -7334 588934
rect -7098 588698 -6916 588934
rect -7516 553254 -6916 588698
rect -7516 553018 -7334 553254
rect -7098 553018 -6916 553254
rect -7516 552934 -6916 553018
rect -7516 552698 -7334 552934
rect -7098 552698 -6916 552934
rect -7516 517254 -6916 552698
rect -7516 517018 -7334 517254
rect -7098 517018 -6916 517254
rect -7516 516934 -6916 517018
rect -7516 516698 -7334 516934
rect -7098 516698 -6916 516934
rect -7516 481254 -6916 516698
rect -7516 481018 -7334 481254
rect -7098 481018 -6916 481254
rect -7516 480934 -6916 481018
rect -7516 480698 -7334 480934
rect -7098 480698 -6916 480934
rect -7516 445254 -6916 480698
rect -7516 445018 -7334 445254
rect -7098 445018 -6916 445254
rect -7516 444934 -6916 445018
rect -7516 444698 -7334 444934
rect -7098 444698 -6916 444934
rect -7516 409254 -6916 444698
rect -7516 409018 -7334 409254
rect -7098 409018 -6916 409254
rect -7516 408934 -6916 409018
rect -7516 408698 -7334 408934
rect -7098 408698 -6916 408934
rect -7516 373254 -6916 408698
rect -7516 373018 -7334 373254
rect -7098 373018 -6916 373254
rect -7516 372934 -6916 373018
rect -7516 372698 -7334 372934
rect -7098 372698 -6916 372934
rect -7516 337254 -6916 372698
rect -7516 337018 -7334 337254
rect -7098 337018 -6916 337254
rect -7516 336934 -6916 337018
rect -7516 336698 -7334 336934
rect -7098 336698 -6916 336934
rect -7516 301254 -6916 336698
rect -7516 301018 -7334 301254
rect -7098 301018 -6916 301254
rect -7516 300934 -6916 301018
rect -7516 300698 -7334 300934
rect -7098 300698 -6916 300934
rect -7516 265254 -6916 300698
rect -7516 265018 -7334 265254
rect -7098 265018 -6916 265254
rect -7516 264934 -6916 265018
rect -7516 264698 -7334 264934
rect -7098 264698 -6916 264934
rect -7516 229254 -6916 264698
rect -7516 229018 -7334 229254
rect -7098 229018 -6916 229254
rect -7516 228934 -6916 229018
rect -7516 228698 -7334 228934
rect -7098 228698 -6916 228934
rect -7516 193254 -6916 228698
rect -7516 193018 -7334 193254
rect -7098 193018 -6916 193254
rect -7516 192934 -6916 193018
rect -7516 192698 -7334 192934
rect -7098 192698 -6916 192934
rect -7516 157254 -6916 192698
rect -7516 157018 -7334 157254
rect -7098 157018 -6916 157254
rect -7516 156934 -6916 157018
rect -7516 156698 -7334 156934
rect -7098 156698 -6916 156934
rect -7516 121254 -6916 156698
rect -7516 121018 -7334 121254
rect -7098 121018 -6916 121254
rect -7516 120934 -6916 121018
rect -7516 120698 -7334 120934
rect -7098 120698 -6916 120934
rect -7516 85254 -6916 120698
rect -7516 85018 -7334 85254
rect -7098 85018 -6916 85254
rect -7516 84934 -6916 85018
rect -7516 84698 -7334 84934
rect -7098 84698 -6916 84934
rect -7516 49254 -6916 84698
rect -7516 49018 -7334 49254
rect -7098 49018 -6916 49254
rect -7516 48934 -6916 49018
rect -7516 48698 -7334 48934
rect -7098 48698 -6916 48934
rect -7516 13254 -6916 48698
rect -7516 13018 -7334 13254
rect -7098 13018 -6916 13254
rect -7516 12934 -6916 13018
rect -7516 12698 -7334 12934
rect -7098 12698 -6916 12934
rect -7516 -5866 -6916 12698
rect -6596 709438 -5996 709460
rect -6596 709202 -6414 709438
rect -6178 709202 -5996 709438
rect -6596 709118 -5996 709202
rect -6596 708882 -6414 709118
rect -6178 708882 -5996 709118
rect -6596 675654 -5996 708882
rect -6596 675418 -6414 675654
rect -6178 675418 -5996 675654
rect -6596 675334 -5996 675418
rect -6596 675098 -6414 675334
rect -6178 675098 -5996 675334
rect -6596 639654 -5996 675098
rect -6596 639418 -6414 639654
rect -6178 639418 -5996 639654
rect -6596 639334 -5996 639418
rect -6596 639098 -6414 639334
rect -6178 639098 -5996 639334
rect -6596 603654 -5996 639098
rect -6596 603418 -6414 603654
rect -6178 603418 -5996 603654
rect -6596 603334 -5996 603418
rect -6596 603098 -6414 603334
rect -6178 603098 -5996 603334
rect -6596 567654 -5996 603098
rect -6596 567418 -6414 567654
rect -6178 567418 -5996 567654
rect -6596 567334 -5996 567418
rect -6596 567098 -6414 567334
rect -6178 567098 -5996 567334
rect -6596 531654 -5996 567098
rect -6596 531418 -6414 531654
rect -6178 531418 -5996 531654
rect -6596 531334 -5996 531418
rect -6596 531098 -6414 531334
rect -6178 531098 -5996 531334
rect -6596 495654 -5996 531098
rect -6596 495418 -6414 495654
rect -6178 495418 -5996 495654
rect -6596 495334 -5996 495418
rect -6596 495098 -6414 495334
rect -6178 495098 -5996 495334
rect -6596 459654 -5996 495098
rect -6596 459418 -6414 459654
rect -6178 459418 -5996 459654
rect -6596 459334 -5996 459418
rect -6596 459098 -6414 459334
rect -6178 459098 -5996 459334
rect -6596 423654 -5996 459098
rect -6596 423418 -6414 423654
rect -6178 423418 -5996 423654
rect -6596 423334 -5996 423418
rect -6596 423098 -6414 423334
rect -6178 423098 -5996 423334
rect -6596 387654 -5996 423098
rect -6596 387418 -6414 387654
rect -6178 387418 -5996 387654
rect -6596 387334 -5996 387418
rect -6596 387098 -6414 387334
rect -6178 387098 -5996 387334
rect -6596 351654 -5996 387098
rect -6596 351418 -6414 351654
rect -6178 351418 -5996 351654
rect -6596 351334 -5996 351418
rect -6596 351098 -6414 351334
rect -6178 351098 -5996 351334
rect -6596 315654 -5996 351098
rect -6596 315418 -6414 315654
rect -6178 315418 -5996 315654
rect -6596 315334 -5996 315418
rect -6596 315098 -6414 315334
rect -6178 315098 -5996 315334
rect -6596 279654 -5996 315098
rect -6596 279418 -6414 279654
rect -6178 279418 -5996 279654
rect -6596 279334 -5996 279418
rect -6596 279098 -6414 279334
rect -6178 279098 -5996 279334
rect -6596 243654 -5996 279098
rect -6596 243418 -6414 243654
rect -6178 243418 -5996 243654
rect -6596 243334 -5996 243418
rect -6596 243098 -6414 243334
rect -6178 243098 -5996 243334
rect -6596 207654 -5996 243098
rect -6596 207418 -6414 207654
rect -6178 207418 -5996 207654
rect -6596 207334 -5996 207418
rect -6596 207098 -6414 207334
rect -6178 207098 -5996 207334
rect -6596 171654 -5996 207098
rect -6596 171418 -6414 171654
rect -6178 171418 -5996 171654
rect -6596 171334 -5996 171418
rect -6596 171098 -6414 171334
rect -6178 171098 -5996 171334
rect -6596 135654 -5996 171098
rect -6596 135418 -6414 135654
rect -6178 135418 -5996 135654
rect -6596 135334 -5996 135418
rect -6596 135098 -6414 135334
rect -6178 135098 -5996 135334
rect -6596 99654 -5996 135098
rect -6596 99418 -6414 99654
rect -6178 99418 -5996 99654
rect -6596 99334 -5996 99418
rect -6596 99098 -6414 99334
rect -6178 99098 -5996 99334
rect -6596 63654 -5996 99098
rect -6596 63418 -6414 63654
rect -6178 63418 -5996 63654
rect -6596 63334 -5996 63418
rect -6596 63098 -6414 63334
rect -6178 63098 -5996 63334
rect -6596 27654 -5996 63098
rect -6596 27418 -6414 27654
rect -6178 27418 -5996 27654
rect -6596 27334 -5996 27418
rect -6596 27098 -6414 27334
rect -6178 27098 -5996 27334
rect -6596 -4946 -5996 27098
rect -5676 708518 -5076 708540
rect -5676 708282 -5494 708518
rect -5258 708282 -5076 708518
rect -5676 708198 -5076 708282
rect -5676 707962 -5494 708198
rect -5258 707962 -5076 708198
rect -5676 693654 -5076 707962
rect 8004 708518 8604 709460
rect 8004 708282 8186 708518
rect 8422 708282 8604 708518
rect 8004 708198 8604 708282
rect 8004 707962 8186 708198
rect 8422 707962 8604 708198
rect -5676 693418 -5494 693654
rect -5258 693418 -5076 693654
rect -5676 693334 -5076 693418
rect -5676 693098 -5494 693334
rect -5258 693098 -5076 693334
rect -5676 657654 -5076 693098
rect -5676 657418 -5494 657654
rect -5258 657418 -5076 657654
rect -5676 657334 -5076 657418
rect -5676 657098 -5494 657334
rect -5258 657098 -5076 657334
rect -5676 621654 -5076 657098
rect -5676 621418 -5494 621654
rect -5258 621418 -5076 621654
rect -5676 621334 -5076 621418
rect -5676 621098 -5494 621334
rect -5258 621098 -5076 621334
rect -5676 585654 -5076 621098
rect -5676 585418 -5494 585654
rect -5258 585418 -5076 585654
rect -5676 585334 -5076 585418
rect -5676 585098 -5494 585334
rect -5258 585098 -5076 585334
rect -5676 549654 -5076 585098
rect -5676 549418 -5494 549654
rect -5258 549418 -5076 549654
rect -5676 549334 -5076 549418
rect -5676 549098 -5494 549334
rect -5258 549098 -5076 549334
rect -5676 513654 -5076 549098
rect -5676 513418 -5494 513654
rect -5258 513418 -5076 513654
rect -5676 513334 -5076 513418
rect -5676 513098 -5494 513334
rect -5258 513098 -5076 513334
rect -5676 477654 -5076 513098
rect -5676 477418 -5494 477654
rect -5258 477418 -5076 477654
rect -5676 477334 -5076 477418
rect -5676 477098 -5494 477334
rect -5258 477098 -5076 477334
rect -5676 441654 -5076 477098
rect -5676 441418 -5494 441654
rect -5258 441418 -5076 441654
rect -5676 441334 -5076 441418
rect -5676 441098 -5494 441334
rect -5258 441098 -5076 441334
rect -5676 405654 -5076 441098
rect -5676 405418 -5494 405654
rect -5258 405418 -5076 405654
rect -5676 405334 -5076 405418
rect -5676 405098 -5494 405334
rect -5258 405098 -5076 405334
rect -5676 369654 -5076 405098
rect -5676 369418 -5494 369654
rect -5258 369418 -5076 369654
rect -5676 369334 -5076 369418
rect -5676 369098 -5494 369334
rect -5258 369098 -5076 369334
rect -5676 333654 -5076 369098
rect -5676 333418 -5494 333654
rect -5258 333418 -5076 333654
rect -5676 333334 -5076 333418
rect -5676 333098 -5494 333334
rect -5258 333098 -5076 333334
rect -5676 297654 -5076 333098
rect -5676 297418 -5494 297654
rect -5258 297418 -5076 297654
rect -5676 297334 -5076 297418
rect -5676 297098 -5494 297334
rect -5258 297098 -5076 297334
rect -5676 261654 -5076 297098
rect -5676 261418 -5494 261654
rect -5258 261418 -5076 261654
rect -5676 261334 -5076 261418
rect -5676 261098 -5494 261334
rect -5258 261098 -5076 261334
rect -5676 225654 -5076 261098
rect -5676 225418 -5494 225654
rect -5258 225418 -5076 225654
rect -5676 225334 -5076 225418
rect -5676 225098 -5494 225334
rect -5258 225098 -5076 225334
rect -5676 189654 -5076 225098
rect -5676 189418 -5494 189654
rect -5258 189418 -5076 189654
rect -5676 189334 -5076 189418
rect -5676 189098 -5494 189334
rect -5258 189098 -5076 189334
rect -5676 153654 -5076 189098
rect -5676 153418 -5494 153654
rect -5258 153418 -5076 153654
rect -5676 153334 -5076 153418
rect -5676 153098 -5494 153334
rect -5258 153098 -5076 153334
rect -5676 117654 -5076 153098
rect -5676 117418 -5494 117654
rect -5258 117418 -5076 117654
rect -5676 117334 -5076 117418
rect -5676 117098 -5494 117334
rect -5258 117098 -5076 117334
rect -5676 81654 -5076 117098
rect -5676 81418 -5494 81654
rect -5258 81418 -5076 81654
rect -5676 81334 -5076 81418
rect -5676 81098 -5494 81334
rect -5258 81098 -5076 81334
rect -5676 45654 -5076 81098
rect -5676 45418 -5494 45654
rect -5258 45418 -5076 45654
rect -5676 45334 -5076 45418
rect -5676 45098 -5494 45334
rect -5258 45098 -5076 45334
rect -5676 9654 -5076 45098
rect -5676 9418 -5494 9654
rect -5258 9418 -5076 9654
rect -5676 9334 -5076 9418
rect -5676 9098 -5494 9334
rect -5258 9098 -5076 9334
rect -5676 -4026 -5076 9098
rect -4756 707598 -4156 707620
rect -4756 707362 -4574 707598
rect -4338 707362 -4156 707598
rect -4756 707278 -4156 707362
rect -4756 707042 -4574 707278
rect -4338 707042 -4156 707278
rect -4756 672054 -4156 707042
rect -4756 671818 -4574 672054
rect -4338 671818 -4156 672054
rect -4756 671734 -4156 671818
rect -4756 671498 -4574 671734
rect -4338 671498 -4156 671734
rect -4756 636054 -4156 671498
rect -4756 635818 -4574 636054
rect -4338 635818 -4156 636054
rect -4756 635734 -4156 635818
rect -4756 635498 -4574 635734
rect -4338 635498 -4156 635734
rect -4756 600054 -4156 635498
rect -4756 599818 -4574 600054
rect -4338 599818 -4156 600054
rect -4756 599734 -4156 599818
rect -4756 599498 -4574 599734
rect -4338 599498 -4156 599734
rect -4756 564054 -4156 599498
rect -4756 563818 -4574 564054
rect -4338 563818 -4156 564054
rect -4756 563734 -4156 563818
rect -4756 563498 -4574 563734
rect -4338 563498 -4156 563734
rect -4756 528054 -4156 563498
rect -4756 527818 -4574 528054
rect -4338 527818 -4156 528054
rect -4756 527734 -4156 527818
rect -4756 527498 -4574 527734
rect -4338 527498 -4156 527734
rect -4756 492054 -4156 527498
rect -4756 491818 -4574 492054
rect -4338 491818 -4156 492054
rect -4756 491734 -4156 491818
rect -4756 491498 -4574 491734
rect -4338 491498 -4156 491734
rect -4756 456054 -4156 491498
rect -4756 455818 -4574 456054
rect -4338 455818 -4156 456054
rect -4756 455734 -4156 455818
rect -4756 455498 -4574 455734
rect -4338 455498 -4156 455734
rect -4756 420054 -4156 455498
rect -4756 419818 -4574 420054
rect -4338 419818 -4156 420054
rect -4756 419734 -4156 419818
rect -4756 419498 -4574 419734
rect -4338 419498 -4156 419734
rect -4756 384054 -4156 419498
rect -4756 383818 -4574 384054
rect -4338 383818 -4156 384054
rect -4756 383734 -4156 383818
rect -4756 383498 -4574 383734
rect -4338 383498 -4156 383734
rect -4756 348054 -4156 383498
rect -4756 347818 -4574 348054
rect -4338 347818 -4156 348054
rect -4756 347734 -4156 347818
rect -4756 347498 -4574 347734
rect -4338 347498 -4156 347734
rect -4756 312054 -4156 347498
rect -4756 311818 -4574 312054
rect -4338 311818 -4156 312054
rect -4756 311734 -4156 311818
rect -4756 311498 -4574 311734
rect -4338 311498 -4156 311734
rect -4756 276054 -4156 311498
rect -4756 275818 -4574 276054
rect -4338 275818 -4156 276054
rect -4756 275734 -4156 275818
rect -4756 275498 -4574 275734
rect -4338 275498 -4156 275734
rect -4756 240054 -4156 275498
rect -4756 239818 -4574 240054
rect -4338 239818 -4156 240054
rect -4756 239734 -4156 239818
rect -4756 239498 -4574 239734
rect -4338 239498 -4156 239734
rect -4756 204054 -4156 239498
rect -4756 203818 -4574 204054
rect -4338 203818 -4156 204054
rect -4756 203734 -4156 203818
rect -4756 203498 -4574 203734
rect -4338 203498 -4156 203734
rect -4756 168054 -4156 203498
rect -4756 167818 -4574 168054
rect -4338 167818 -4156 168054
rect -4756 167734 -4156 167818
rect -4756 167498 -4574 167734
rect -4338 167498 -4156 167734
rect -4756 132054 -4156 167498
rect -4756 131818 -4574 132054
rect -4338 131818 -4156 132054
rect -4756 131734 -4156 131818
rect -4756 131498 -4574 131734
rect -4338 131498 -4156 131734
rect -4756 96054 -4156 131498
rect -4756 95818 -4574 96054
rect -4338 95818 -4156 96054
rect -4756 95734 -4156 95818
rect -4756 95498 -4574 95734
rect -4338 95498 -4156 95734
rect -4756 60054 -4156 95498
rect -4756 59818 -4574 60054
rect -4338 59818 -4156 60054
rect -4756 59734 -4156 59818
rect -4756 59498 -4574 59734
rect -4338 59498 -4156 59734
rect -4756 24054 -4156 59498
rect -4756 23818 -4574 24054
rect -4338 23818 -4156 24054
rect -4756 23734 -4156 23818
rect -4756 23498 -4574 23734
rect -4338 23498 -4156 23734
rect -4756 -3106 -4156 23498
rect -3836 706678 -3236 706700
rect -3836 706442 -3654 706678
rect -3418 706442 -3236 706678
rect -3836 706358 -3236 706442
rect -3836 706122 -3654 706358
rect -3418 706122 -3236 706358
rect -3836 690054 -3236 706122
rect 4404 706678 5004 707620
rect 4404 706442 4586 706678
rect 4822 706442 5004 706678
rect 4404 706358 5004 706442
rect 4404 706122 4586 706358
rect 4822 706122 5004 706358
rect -3836 689818 -3654 690054
rect -3418 689818 -3236 690054
rect -3836 689734 -3236 689818
rect -3836 689498 -3654 689734
rect -3418 689498 -3236 689734
rect -3836 654054 -3236 689498
rect -3836 653818 -3654 654054
rect -3418 653818 -3236 654054
rect -3836 653734 -3236 653818
rect -3836 653498 -3654 653734
rect -3418 653498 -3236 653734
rect -3836 618054 -3236 653498
rect -3836 617818 -3654 618054
rect -3418 617818 -3236 618054
rect -3836 617734 -3236 617818
rect -3836 617498 -3654 617734
rect -3418 617498 -3236 617734
rect -3836 582054 -3236 617498
rect -3836 581818 -3654 582054
rect -3418 581818 -3236 582054
rect -3836 581734 -3236 581818
rect -3836 581498 -3654 581734
rect -3418 581498 -3236 581734
rect -3836 546054 -3236 581498
rect -3836 545818 -3654 546054
rect -3418 545818 -3236 546054
rect -3836 545734 -3236 545818
rect -3836 545498 -3654 545734
rect -3418 545498 -3236 545734
rect -3836 510054 -3236 545498
rect -3836 509818 -3654 510054
rect -3418 509818 -3236 510054
rect -3836 509734 -3236 509818
rect -3836 509498 -3654 509734
rect -3418 509498 -3236 509734
rect -3836 474054 -3236 509498
rect -3836 473818 -3654 474054
rect -3418 473818 -3236 474054
rect -3836 473734 -3236 473818
rect -3836 473498 -3654 473734
rect -3418 473498 -3236 473734
rect -3836 438054 -3236 473498
rect -3836 437818 -3654 438054
rect -3418 437818 -3236 438054
rect -3836 437734 -3236 437818
rect -3836 437498 -3654 437734
rect -3418 437498 -3236 437734
rect -3836 402054 -3236 437498
rect -3836 401818 -3654 402054
rect -3418 401818 -3236 402054
rect -3836 401734 -3236 401818
rect -3836 401498 -3654 401734
rect -3418 401498 -3236 401734
rect -3836 366054 -3236 401498
rect -3836 365818 -3654 366054
rect -3418 365818 -3236 366054
rect -3836 365734 -3236 365818
rect -3836 365498 -3654 365734
rect -3418 365498 -3236 365734
rect -3836 330054 -3236 365498
rect -3836 329818 -3654 330054
rect -3418 329818 -3236 330054
rect -3836 329734 -3236 329818
rect -3836 329498 -3654 329734
rect -3418 329498 -3236 329734
rect -3836 294054 -3236 329498
rect -3836 293818 -3654 294054
rect -3418 293818 -3236 294054
rect -3836 293734 -3236 293818
rect -3836 293498 -3654 293734
rect -3418 293498 -3236 293734
rect -3836 258054 -3236 293498
rect -3836 257818 -3654 258054
rect -3418 257818 -3236 258054
rect -3836 257734 -3236 257818
rect -3836 257498 -3654 257734
rect -3418 257498 -3236 257734
rect -3836 222054 -3236 257498
rect -3836 221818 -3654 222054
rect -3418 221818 -3236 222054
rect -3836 221734 -3236 221818
rect -3836 221498 -3654 221734
rect -3418 221498 -3236 221734
rect -3836 186054 -3236 221498
rect -3836 185818 -3654 186054
rect -3418 185818 -3236 186054
rect -3836 185734 -3236 185818
rect -3836 185498 -3654 185734
rect -3418 185498 -3236 185734
rect -3836 150054 -3236 185498
rect -3836 149818 -3654 150054
rect -3418 149818 -3236 150054
rect -3836 149734 -3236 149818
rect -3836 149498 -3654 149734
rect -3418 149498 -3236 149734
rect -3836 114054 -3236 149498
rect -3836 113818 -3654 114054
rect -3418 113818 -3236 114054
rect -3836 113734 -3236 113818
rect -3836 113498 -3654 113734
rect -3418 113498 -3236 113734
rect -3836 78054 -3236 113498
rect -3836 77818 -3654 78054
rect -3418 77818 -3236 78054
rect -3836 77734 -3236 77818
rect -3836 77498 -3654 77734
rect -3418 77498 -3236 77734
rect -3836 42054 -3236 77498
rect -3836 41818 -3654 42054
rect -3418 41818 -3236 42054
rect -3836 41734 -3236 41818
rect -3836 41498 -3654 41734
rect -3418 41498 -3236 41734
rect -3836 6054 -3236 41498
rect -3836 5818 -3654 6054
rect -3418 5818 -3236 6054
rect -3836 5734 -3236 5818
rect -3836 5498 -3654 5734
rect -3418 5498 -3236 5734
rect -3836 -2186 -3236 5498
rect -2916 705758 -2316 705780
rect -2916 705522 -2734 705758
rect -2498 705522 -2316 705758
rect -2916 705438 -2316 705522
rect -2916 705202 -2734 705438
rect -2498 705202 -2316 705438
rect -2916 668454 -2316 705202
rect -2916 668218 -2734 668454
rect -2498 668218 -2316 668454
rect -2916 668134 -2316 668218
rect -2916 667898 -2734 668134
rect -2498 667898 -2316 668134
rect -2916 632454 -2316 667898
rect -2916 632218 -2734 632454
rect -2498 632218 -2316 632454
rect -2916 632134 -2316 632218
rect -2916 631898 -2734 632134
rect -2498 631898 -2316 632134
rect -2916 596454 -2316 631898
rect -2916 596218 -2734 596454
rect -2498 596218 -2316 596454
rect -2916 596134 -2316 596218
rect -2916 595898 -2734 596134
rect -2498 595898 -2316 596134
rect -2916 560454 -2316 595898
rect -2916 560218 -2734 560454
rect -2498 560218 -2316 560454
rect -2916 560134 -2316 560218
rect -2916 559898 -2734 560134
rect -2498 559898 -2316 560134
rect -2916 524454 -2316 559898
rect -2916 524218 -2734 524454
rect -2498 524218 -2316 524454
rect -2916 524134 -2316 524218
rect -2916 523898 -2734 524134
rect -2498 523898 -2316 524134
rect -2916 488454 -2316 523898
rect -2916 488218 -2734 488454
rect -2498 488218 -2316 488454
rect -2916 488134 -2316 488218
rect -2916 487898 -2734 488134
rect -2498 487898 -2316 488134
rect -2916 452454 -2316 487898
rect -2916 452218 -2734 452454
rect -2498 452218 -2316 452454
rect -2916 452134 -2316 452218
rect -2916 451898 -2734 452134
rect -2498 451898 -2316 452134
rect -2916 416454 -2316 451898
rect -2916 416218 -2734 416454
rect -2498 416218 -2316 416454
rect -2916 416134 -2316 416218
rect -2916 415898 -2734 416134
rect -2498 415898 -2316 416134
rect -2916 380454 -2316 415898
rect -2916 380218 -2734 380454
rect -2498 380218 -2316 380454
rect -2916 380134 -2316 380218
rect -2916 379898 -2734 380134
rect -2498 379898 -2316 380134
rect -2916 344454 -2316 379898
rect -2916 344218 -2734 344454
rect -2498 344218 -2316 344454
rect -2916 344134 -2316 344218
rect -2916 343898 -2734 344134
rect -2498 343898 -2316 344134
rect -2916 308454 -2316 343898
rect -2916 308218 -2734 308454
rect -2498 308218 -2316 308454
rect -2916 308134 -2316 308218
rect -2916 307898 -2734 308134
rect -2498 307898 -2316 308134
rect -2916 272454 -2316 307898
rect -2916 272218 -2734 272454
rect -2498 272218 -2316 272454
rect -2916 272134 -2316 272218
rect -2916 271898 -2734 272134
rect -2498 271898 -2316 272134
rect -2916 236454 -2316 271898
rect -2916 236218 -2734 236454
rect -2498 236218 -2316 236454
rect -2916 236134 -2316 236218
rect -2916 235898 -2734 236134
rect -2498 235898 -2316 236134
rect -2916 200454 -2316 235898
rect -2916 200218 -2734 200454
rect -2498 200218 -2316 200454
rect -2916 200134 -2316 200218
rect -2916 199898 -2734 200134
rect -2498 199898 -2316 200134
rect -2916 164454 -2316 199898
rect -2916 164218 -2734 164454
rect -2498 164218 -2316 164454
rect -2916 164134 -2316 164218
rect -2916 163898 -2734 164134
rect -2498 163898 -2316 164134
rect -2916 128454 -2316 163898
rect -2916 128218 -2734 128454
rect -2498 128218 -2316 128454
rect -2916 128134 -2316 128218
rect -2916 127898 -2734 128134
rect -2498 127898 -2316 128134
rect -2916 92454 -2316 127898
rect -2916 92218 -2734 92454
rect -2498 92218 -2316 92454
rect -2916 92134 -2316 92218
rect -2916 91898 -2734 92134
rect -2498 91898 -2316 92134
rect -2916 56454 -2316 91898
rect -2916 56218 -2734 56454
rect -2498 56218 -2316 56454
rect -2916 56134 -2316 56218
rect -2916 55898 -2734 56134
rect -2498 55898 -2316 56134
rect -2916 20454 -2316 55898
rect -2916 20218 -2734 20454
rect -2498 20218 -2316 20454
rect -2916 20134 -2316 20218
rect -2916 19898 -2734 20134
rect -2498 19898 -2316 20134
rect -2916 -1266 -2316 19898
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 686454 -1396 704282
rect -1996 686218 -1814 686454
rect -1578 686218 -1396 686454
rect -1996 686134 -1396 686218
rect -1996 685898 -1814 686134
rect -1578 685898 -1396 686134
rect -1996 650454 -1396 685898
rect -1996 650218 -1814 650454
rect -1578 650218 -1396 650454
rect -1996 650134 -1396 650218
rect -1996 649898 -1814 650134
rect -1578 649898 -1396 650134
rect -1996 614454 -1396 649898
rect -1996 614218 -1814 614454
rect -1578 614218 -1396 614454
rect -1996 614134 -1396 614218
rect -1996 613898 -1814 614134
rect -1578 613898 -1396 614134
rect -1996 578454 -1396 613898
rect -1996 578218 -1814 578454
rect -1578 578218 -1396 578454
rect -1996 578134 -1396 578218
rect -1996 577898 -1814 578134
rect -1578 577898 -1396 578134
rect -1996 542454 -1396 577898
rect -1996 542218 -1814 542454
rect -1578 542218 -1396 542454
rect -1996 542134 -1396 542218
rect -1996 541898 -1814 542134
rect -1578 541898 -1396 542134
rect -1996 506454 -1396 541898
rect -1996 506218 -1814 506454
rect -1578 506218 -1396 506454
rect -1996 506134 -1396 506218
rect -1996 505898 -1814 506134
rect -1578 505898 -1396 506134
rect -1996 470454 -1396 505898
rect -1996 470218 -1814 470454
rect -1578 470218 -1396 470454
rect -1996 470134 -1396 470218
rect -1996 469898 -1814 470134
rect -1578 469898 -1396 470134
rect -1996 434454 -1396 469898
rect -1996 434218 -1814 434454
rect -1578 434218 -1396 434454
rect -1996 434134 -1396 434218
rect -1996 433898 -1814 434134
rect -1578 433898 -1396 434134
rect -1996 398454 -1396 433898
rect -1996 398218 -1814 398454
rect -1578 398218 -1396 398454
rect -1996 398134 -1396 398218
rect -1996 397898 -1814 398134
rect -1578 397898 -1396 398134
rect -1996 362454 -1396 397898
rect -1996 362218 -1814 362454
rect -1578 362218 -1396 362454
rect -1996 362134 -1396 362218
rect -1996 361898 -1814 362134
rect -1578 361898 -1396 362134
rect -1996 326454 -1396 361898
rect -1996 326218 -1814 326454
rect -1578 326218 -1396 326454
rect -1996 326134 -1396 326218
rect -1996 325898 -1814 326134
rect -1578 325898 -1396 326134
rect -1996 290454 -1396 325898
rect -1996 290218 -1814 290454
rect -1578 290218 -1396 290454
rect -1996 290134 -1396 290218
rect -1996 289898 -1814 290134
rect -1578 289898 -1396 290134
rect -1996 254454 -1396 289898
rect -1996 254218 -1814 254454
rect -1578 254218 -1396 254454
rect -1996 254134 -1396 254218
rect -1996 253898 -1814 254134
rect -1578 253898 -1396 254134
rect -1996 218454 -1396 253898
rect -1996 218218 -1814 218454
rect -1578 218218 -1396 218454
rect -1996 218134 -1396 218218
rect -1996 217898 -1814 218134
rect -1578 217898 -1396 218134
rect -1996 182454 -1396 217898
rect -1996 182218 -1814 182454
rect -1578 182218 -1396 182454
rect -1996 182134 -1396 182218
rect -1996 181898 -1814 182134
rect -1578 181898 -1396 182134
rect -1996 146454 -1396 181898
rect -1996 146218 -1814 146454
rect -1578 146218 -1396 146454
rect -1996 146134 -1396 146218
rect -1996 145898 -1814 146134
rect -1578 145898 -1396 146134
rect -1996 110454 -1396 145898
rect -1996 110218 -1814 110454
rect -1578 110218 -1396 110454
rect -1996 110134 -1396 110218
rect -1996 109898 -1814 110134
rect -1578 109898 -1396 110134
rect -1996 74454 -1396 109898
rect -1996 74218 -1814 74454
rect -1578 74218 -1396 74454
rect -1996 74134 -1396 74218
rect -1996 73898 -1814 74134
rect -1578 73898 -1396 74134
rect -1996 38454 -1396 73898
rect -1996 38218 -1814 38454
rect -1578 38218 -1396 38454
rect -1996 38134 -1396 38218
rect -1996 37898 -1814 38134
rect -1578 37898 -1396 38134
rect -1996 2454 -1396 37898
rect -1996 2218 -1814 2454
rect -1578 2218 -1396 2454
rect -1996 2134 -1396 2218
rect -1996 1898 -1814 2134
rect -1578 1898 -1396 2134
rect -1996 -346 -1396 1898
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 804 704838 1404 705780
rect 804 704602 986 704838
rect 1222 704602 1404 704838
rect 804 704518 1404 704602
rect 804 704282 986 704518
rect 1222 704282 1404 704518
rect 804 686454 1404 704282
rect 804 686218 986 686454
rect 1222 686218 1404 686454
rect 804 686134 1404 686218
rect 804 685898 986 686134
rect 1222 685898 1404 686134
rect 804 650454 1404 685898
rect 804 650218 986 650454
rect 1222 650218 1404 650454
rect 804 650134 1404 650218
rect 804 649898 986 650134
rect 1222 649898 1404 650134
rect 804 614454 1404 649898
rect 804 614218 986 614454
rect 1222 614218 1404 614454
rect 804 614134 1404 614218
rect 804 613898 986 614134
rect 1222 613898 1404 614134
rect 804 578454 1404 613898
rect 804 578218 986 578454
rect 1222 578218 1404 578454
rect 804 578134 1404 578218
rect 804 577898 986 578134
rect 1222 577898 1404 578134
rect 804 542454 1404 577898
rect 804 542218 986 542454
rect 1222 542218 1404 542454
rect 804 542134 1404 542218
rect 804 541898 986 542134
rect 1222 541898 1404 542134
rect 804 506454 1404 541898
rect 804 506218 986 506454
rect 1222 506218 1404 506454
rect 804 506134 1404 506218
rect 804 505898 986 506134
rect 1222 505898 1404 506134
rect 804 470454 1404 505898
rect 804 470218 986 470454
rect 1222 470218 1404 470454
rect 804 470134 1404 470218
rect 804 469898 986 470134
rect 1222 469898 1404 470134
rect 804 434454 1404 469898
rect 804 434218 986 434454
rect 1222 434218 1404 434454
rect 804 434134 1404 434218
rect 804 433898 986 434134
rect 1222 433898 1404 434134
rect 804 398454 1404 433898
rect 804 398218 986 398454
rect 1222 398218 1404 398454
rect 804 398134 1404 398218
rect 804 397898 986 398134
rect 1222 397898 1404 398134
rect 804 362454 1404 397898
rect 804 362218 986 362454
rect 1222 362218 1404 362454
rect 804 362134 1404 362218
rect 804 361898 986 362134
rect 1222 361898 1404 362134
rect 804 326454 1404 361898
rect 804 326218 986 326454
rect 1222 326218 1404 326454
rect 804 326134 1404 326218
rect 804 325898 986 326134
rect 1222 325898 1404 326134
rect 804 290454 1404 325898
rect 804 290218 986 290454
rect 1222 290218 1404 290454
rect 804 290134 1404 290218
rect 804 289898 986 290134
rect 1222 289898 1404 290134
rect 804 254454 1404 289898
rect 804 254218 986 254454
rect 1222 254218 1404 254454
rect 804 254134 1404 254218
rect 804 253898 986 254134
rect 1222 253898 1404 254134
rect 804 218454 1404 253898
rect 804 218218 986 218454
rect 1222 218218 1404 218454
rect 804 218134 1404 218218
rect 804 217898 986 218134
rect 1222 217898 1404 218134
rect 804 182454 1404 217898
rect 804 182218 986 182454
rect 1222 182218 1404 182454
rect 804 182134 1404 182218
rect 804 181898 986 182134
rect 1222 181898 1404 182134
rect 804 146454 1404 181898
rect 804 146218 986 146454
rect 1222 146218 1404 146454
rect 804 146134 1404 146218
rect 804 145898 986 146134
rect 1222 145898 1404 146134
rect 804 110454 1404 145898
rect 804 110218 986 110454
rect 1222 110218 1404 110454
rect 804 110134 1404 110218
rect 804 109898 986 110134
rect 1222 109898 1404 110134
rect 804 74454 1404 109898
rect 804 74218 986 74454
rect 1222 74218 1404 74454
rect 804 74134 1404 74218
rect 804 73898 986 74134
rect 1222 73898 1404 74134
rect 804 38454 1404 73898
rect 804 38218 986 38454
rect 1222 38218 1404 38454
rect 804 38134 1404 38218
rect 804 37898 986 38134
rect 1222 37898 1404 38134
rect 804 2454 1404 37898
rect 804 2218 986 2454
rect 1222 2218 1404 2454
rect 804 2134 1404 2218
rect 804 1898 986 2134
rect 1222 1898 1404 2134
rect 804 -346 1404 1898
rect 804 -582 986 -346
rect 1222 -582 1404 -346
rect 804 -666 1404 -582
rect 804 -902 986 -666
rect 1222 -902 1404 -666
rect -2916 -1502 -2734 -1266
rect -2498 -1502 -2316 -1266
rect -2916 -1586 -2316 -1502
rect -2916 -1822 -2734 -1586
rect -2498 -1822 -2316 -1586
rect -2916 -1844 -2316 -1822
rect 804 -1844 1404 -902
rect 4404 690054 5004 706122
rect 4404 689818 4586 690054
rect 4822 689818 5004 690054
rect 4404 689734 5004 689818
rect 4404 689498 4586 689734
rect 4822 689498 5004 689734
rect 4404 654054 5004 689498
rect 4404 653818 4586 654054
rect 4822 653818 5004 654054
rect 4404 653734 5004 653818
rect 4404 653498 4586 653734
rect 4822 653498 5004 653734
rect 4404 618054 5004 653498
rect 4404 617818 4586 618054
rect 4822 617818 5004 618054
rect 4404 617734 5004 617818
rect 4404 617498 4586 617734
rect 4822 617498 5004 617734
rect 4404 582054 5004 617498
rect 4404 581818 4586 582054
rect 4822 581818 5004 582054
rect 4404 581734 5004 581818
rect 4404 581498 4586 581734
rect 4822 581498 5004 581734
rect 4404 546054 5004 581498
rect 4404 545818 4586 546054
rect 4822 545818 5004 546054
rect 4404 545734 5004 545818
rect 4404 545498 4586 545734
rect 4822 545498 5004 545734
rect 4404 510054 5004 545498
rect 4404 509818 4586 510054
rect 4822 509818 5004 510054
rect 4404 509734 5004 509818
rect 4404 509498 4586 509734
rect 4822 509498 5004 509734
rect 4404 474054 5004 509498
rect 4404 473818 4586 474054
rect 4822 473818 5004 474054
rect 4404 473734 5004 473818
rect 4404 473498 4586 473734
rect 4822 473498 5004 473734
rect 4404 438054 5004 473498
rect 4404 437818 4586 438054
rect 4822 437818 5004 438054
rect 4404 437734 5004 437818
rect 4404 437498 4586 437734
rect 4822 437498 5004 437734
rect 4404 402054 5004 437498
rect 4404 401818 4586 402054
rect 4822 401818 5004 402054
rect 4404 401734 5004 401818
rect 4404 401498 4586 401734
rect 4822 401498 5004 401734
rect 4404 366054 5004 401498
rect 4404 365818 4586 366054
rect 4822 365818 5004 366054
rect 4404 365734 5004 365818
rect 4404 365498 4586 365734
rect 4822 365498 5004 365734
rect 4404 330054 5004 365498
rect 4404 329818 4586 330054
rect 4822 329818 5004 330054
rect 4404 329734 5004 329818
rect 4404 329498 4586 329734
rect 4822 329498 5004 329734
rect 4404 294054 5004 329498
rect 4404 293818 4586 294054
rect 4822 293818 5004 294054
rect 4404 293734 5004 293818
rect 4404 293498 4586 293734
rect 4822 293498 5004 293734
rect 4404 258054 5004 293498
rect 4404 257818 4586 258054
rect 4822 257818 5004 258054
rect 4404 257734 5004 257818
rect 4404 257498 4586 257734
rect 4822 257498 5004 257734
rect 4404 222054 5004 257498
rect 4404 221818 4586 222054
rect 4822 221818 5004 222054
rect 4404 221734 5004 221818
rect 4404 221498 4586 221734
rect 4822 221498 5004 221734
rect 4404 186054 5004 221498
rect 4404 185818 4586 186054
rect 4822 185818 5004 186054
rect 4404 185734 5004 185818
rect 4404 185498 4586 185734
rect 4822 185498 5004 185734
rect 4404 150054 5004 185498
rect 4404 149818 4586 150054
rect 4822 149818 5004 150054
rect 4404 149734 5004 149818
rect 4404 149498 4586 149734
rect 4822 149498 5004 149734
rect 4404 114054 5004 149498
rect 4404 113818 4586 114054
rect 4822 113818 5004 114054
rect 4404 113734 5004 113818
rect 4404 113498 4586 113734
rect 4822 113498 5004 113734
rect 4404 78054 5004 113498
rect 4404 77818 4586 78054
rect 4822 77818 5004 78054
rect 4404 77734 5004 77818
rect 4404 77498 4586 77734
rect 4822 77498 5004 77734
rect 4404 42054 5004 77498
rect 4404 41818 4586 42054
rect 4822 41818 5004 42054
rect 4404 41734 5004 41818
rect 4404 41498 4586 41734
rect 4822 41498 5004 41734
rect 4404 6054 5004 41498
rect 4404 5818 4586 6054
rect 4822 5818 5004 6054
rect 4404 5734 5004 5818
rect 4404 5498 4586 5734
rect 4822 5498 5004 5734
rect -3836 -2422 -3654 -2186
rect -3418 -2422 -3236 -2186
rect -3836 -2506 -3236 -2422
rect -3836 -2742 -3654 -2506
rect -3418 -2742 -3236 -2506
rect -3836 -2764 -3236 -2742
rect 4404 -2186 5004 5498
rect 4404 -2422 4586 -2186
rect 4822 -2422 5004 -2186
rect 4404 -2506 5004 -2422
rect 4404 -2742 4586 -2506
rect 4822 -2742 5004 -2506
rect -4756 -3342 -4574 -3106
rect -4338 -3342 -4156 -3106
rect -4756 -3426 -4156 -3342
rect -4756 -3662 -4574 -3426
rect -4338 -3662 -4156 -3426
rect -4756 -3684 -4156 -3662
rect 4404 -3684 5004 -2742
rect 8004 693654 8604 707962
rect 8004 693418 8186 693654
rect 8422 693418 8604 693654
rect 8004 693334 8604 693418
rect 8004 693098 8186 693334
rect 8422 693098 8604 693334
rect 8004 657654 8604 693098
rect 8004 657418 8186 657654
rect 8422 657418 8604 657654
rect 8004 657334 8604 657418
rect 8004 657098 8186 657334
rect 8422 657098 8604 657334
rect 8004 621654 8604 657098
rect 8004 621418 8186 621654
rect 8422 621418 8604 621654
rect 8004 621334 8604 621418
rect 8004 621098 8186 621334
rect 8422 621098 8604 621334
rect 8004 585654 8604 621098
rect 8004 585418 8186 585654
rect 8422 585418 8604 585654
rect 8004 585334 8604 585418
rect 8004 585098 8186 585334
rect 8422 585098 8604 585334
rect 8004 549654 8604 585098
rect 8004 549418 8186 549654
rect 8422 549418 8604 549654
rect 8004 549334 8604 549418
rect 8004 549098 8186 549334
rect 8422 549098 8604 549334
rect 8004 513654 8604 549098
rect 8004 513418 8186 513654
rect 8422 513418 8604 513654
rect 8004 513334 8604 513418
rect 8004 513098 8186 513334
rect 8422 513098 8604 513334
rect 8004 477654 8604 513098
rect 8004 477418 8186 477654
rect 8422 477418 8604 477654
rect 8004 477334 8604 477418
rect 8004 477098 8186 477334
rect 8422 477098 8604 477334
rect 8004 441654 8604 477098
rect 8004 441418 8186 441654
rect 8422 441418 8604 441654
rect 8004 441334 8604 441418
rect 8004 441098 8186 441334
rect 8422 441098 8604 441334
rect 8004 405654 8604 441098
rect 8004 405418 8186 405654
rect 8422 405418 8604 405654
rect 8004 405334 8604 405418
rect 8004 405098 8186 405334
rect 8422 405098 8604 405334
rect 8004 369654 8604 405098
rect 8004 369418 8186 369654
rect 8422 369418 8604 369654
rect 8004 369334 8604 369418
rect 8004 369098 8186 369334
rect 8422 369098 8604 369334
rect 8004 333654 8604 369098
rect 8004 333418 8186 333654
rect 8422 333418 8604 333654
rect 8004 333334 8604 333418
rect 8004 333098 8186 333334
rect 8422 333098 8604 333334
rect 8004 297654 8604 333098
rect 8004 297418 8186 297654
rect 8422 297418 8604 297654
rect 8004 297334 8604 297418
rect 8004 297098 8186 297334
rect 8422 297098 8604 297334
rect 8004 261654 8604 297098
rect 8004 261418 8186 261654
rect 8422 261418 8604 261654
rect 8004 261334 8604 261418
rect 8004 261098 8186 261334
rect 8422 261098 8604 261334
rect 8004 225654 8604 261098
rect 8004 225418 8186 225654
rect 8422 225418 8604 225654
rect 8004 225334 8604 225418
rect 8004 225098 8186 225334
rect 8422 225098 8604 225334
rect 8004 189654 8604 225098
rect 8004 189418 8186 189654
rect 8422 189418 8604 189654
rect 8004 189334 8604 189418
rect 8004 189098 8186 189334
rect 8422 189098 8604 189334
rect 8004 153654 8604 189098
rect 8004 153418 8186 153654
rect 8422 153418 8604 153654
rect 8004 153334 8604 153418
rect 8004 153098 8186 153334
rect 8422 153098 8604 153334
rect 8004 117654 8604 153098
rect 8004 117418 8186 117654
rect 8422 117418 8604 117654
rect 8004 117334 8604 117418
rect 8004 117098 8186 117334
rect 8422 117098 8604 117334
rect 8004 81654 8604 117098
rect 8004 81418 8186 81654
rect 8422 81418 8604 81654
rect 8004 81334 8604 81418
rect 8004 81098 8186 81334
rect 8422 81098 8604 81334
rect 8004 45654 8604 81098
rect 8004 45418 8186 45654
rect 8422 45418 8604 45654
rect 8004 45334 8604 45418
rect 8004 45098 8186 45334
rect 8422 45098 8604 45334
rect 8004 9654 8604 45098
rect 8004 9418 8186 9654
rect 8422 9418 8604 9654
rect 8004 9334 8604 9418
rect 8004 9098 8186 9334
rect 8422 9098 8604 9334
rect -5676 -4262 -5494 -4026
rect -5258 -4262 -5076 -4026
rect -5676 -4346 -5076 -4262
rect -5676 -4582 -5494 -4346
rect -5258 -4582 -5076 -4346
rect -5676 -4604 -5076 -4582
rect 8004 -4026 8604 9098
rect 8004 -4262 8186 -4026
rect 8422 -4262 8604 -4026
rect 8004 -4346 8604 -4262
rect 8004 -4582 8186 -4346
rect 8422 -4582 8604 -4346
rect -6596 -5182 -6414 -4946
rect -6178 -5182 -5996 -4946
rect -6596 -5266 -5996 -5182
rect -6596 -5502 -6414 -5266
rect -6178 -5502 -5996 -5266
rect -6596 -5524 -5996 -5502
rect 8004 -5524 8604 -4582
rect 11604 697254 12204 709802
rect 29604 711278 30204 711300
rect 29604 711042 29786 711278
rect 30022 711042 30204 711278
rect 29604 710958 30204 711042
rect 29604 710722 29786 710958
rect 30022 710722 30204 710958
rect 26004 709438 26604 709460
rect 26004 709202 26186 709438
rect 26422 709202 26604 709438
rect 26004 709118 26604 709202
rect 26004 708882 26186 709118
rect 26422 708882 26604 709118
rect 22404 707598 23004 707620
rect 22404 707362 22586 707598
rect 22822 707362 23004 707598
rect 22404 707278 23004 707362
rect 22404 707042 22586 707278
rect 22822 707042 23004 707278
rect 11604 697018 11786 697254
rect 12022 697018 12204 697254
rect 11604 696934 12204 697018
rect 11604 696698 11786 696934
rect 12022 696698 12204 696934
rect 11604 661254 12204 696698
rect 11604 661018 11786 661254
rect 12022 661018 12204 661254
rect 11604 660934 12204 661018
rect 11604 660698 11786 660934
rect 12022 660698 12204 660934
rect 11604 625254 12204 660698
rect 11604 625018 11786 625254
rect 12022 625018 12204 625254
rect 11604 624934 12204 625018
rect 11604 624698 11786 624934
rect 12022 624698 12204 624934
rect 11604 589254 12204 624698
rect 11604 589018 11786 589254
rect 12022 589018 12204 589254
rect 11604 588934 12204 589018
rect 11604 588698 11786 588934
rect 12022 588698 12204 588934
rect 11604 553254 12204 588698
rect 11604 553018 11786 553254
rect 12022 553018 12204 553254
rect 11604 552934 12204 553018
rect 11604 552698 11786 552934
rect 12022 552698 12204 552934
rect 11604 517254 12204 552698
rect 11604 517018 11786 517254
rect 12022 517018 12204 517254
rect 11604 516934 12204 517018
rect 11604 516698 11786 516934
rect 12022 516698 12204 516934
rect 11604 481254 12204 516698
rect 11604 481018 11786 481254
rect 12022 481018 12204 481254
rect 11604 480934 12204 481018
rect 11604 480698 11786 480934
rect 12022 480698 12204 480934
rect 11604 445254 12204 480698
rect 11604 445018 11786 445254
rect 12022 445018 12204 445254
rect 11604 444934 12204 445018
rect 11604 444698 11786 444934
rect 12022 444698 12204 444934
rect 11604 409254 12204 444698
rect 11604 409018 11786 409254
rect 12022 409018 12204 409254
rect 11604 408934 12204 409018
rect 11604 408698 11786 408934
rect 12022 408698 12204 408934
rect 11604 373254 12204 408698
rect 11604 373018 11786 373254
rect 12022 373018 12204 373254
rect 11604 372934 12204 373018
rect 11604 372698 11786 372934
rect 12022 372698 12204 372934
rect 11604 337254 12204 372698
rect 11604 337018 11786 337254
rect 12022 337018 12204 337254
rect 11604 336934 12204 337018
rect 11604 336698 11786 336934
rect 12022 336698 12204 336934
rect 11604 301254 12204 336698
rect 11604 301018 11786 301254
rect 12022 301018 12204 301254
rect 11604 300934 12204 301018
rect 11604 300698 11786 300934
rect 12022 300698 12204 300934
rect 11604 265254 12204 300698
rect 11604 265018 11786 265254
rect 12022 265018 12204 265254
rect 11604 264934 12204 265018
rect 11604 264698 11786 264934
rect 12022 264698 12204 264934
rect 11604 229254 12204 264698
rect 11604 229018 11786 229254
rect 12022 229018 12204 229254
rect 11604 228934 12204 229018
rect 11604 228698 11786 228934
rect 12022 228698 12204 228934
rect 11604 193254 12204 228698
rect 11604 193018 11786 193254
rect 12022 193018 12204 193254
rect 11604 192934 12204 193018
rect 11604 192698 11786 192934
rect 12022 192698 12204 192934
rect 11604 157254 12204 192698
rect 11604 157018 11786 157254
rect 12022 157018 12204 157254
rect 11604 156934 12204 157018
rect 11604 156698 11786 156934
rect 12022 156698 12204 156934
rect 11604 121254 12204 156698
rect 11604 121018 11786 121254
rect 12022 121018 12204 121254
rect 11604 120934 12204 121018
rect 11604 120698 11786 120934
rect 12022 120698 12204 120934
rect 11604 85254 12204 120698
rect 11604 85018 11786 85254
rect 12022 85018 12204 85254
rect 11604 84934 12204 85018
rect 11604 84698 11786 84934
rect 12022 84698 12204 84934
rect 11604 49254 12204 84698
rect 11604 49018 11786 49254
rect 12022 49018 12204 49254
rect 11604 48934 12204 49018
rect 11604 48698 11786 48934
rect 12022 48698 12204 48934
rect 11604 13254 12204 48698
rect 11604 13018 11786 13254
rect 12022 13018 12204 13254
rect 11604 12934 12204 13018
rect 11604 12698 11786 12934
rect 12022 12698 12204 12934
rect -7516 -6102 -7334 -5866
rect -7098 -6102 -6916 -5866
rect -7516 -6186 -6916 -6102
rect -7516 -6422 -7334 -6186
rect -7098 -6422 -6916 -6186
rect -7516 -6444 -6916 -6422
rect 11604 -5866 12204 12698
rect 18804 705758 19404 705780
rect 18804 705522 18986 705758
rect 19222 705522 19404 705758
rect 18804 705438 19404 705522
rect 18804 705202 18986 705438
rect 19222 705202 19404 705438
rect 18804 668454 19404 705202
rect 18804 668218 18986 668454
rect 19222 668218 19404 668454
rect 18804 668134 19404 668218
rect 18804 667898 18986 668134
rect 19222 667898 19404 668134
rect 18804 632454 19404 667898
rect 18804 632218 18986 632454
rect 19222 632218 19404 632454
rect 18804 632134 19404 632218
rect 18804 631898 18986 632134
rect 19222 631898 19404 632134
rect 18804 596454 19404 631898
rect 18804 596218 18986 596454
rect 19222 596218 19404 596454
rect 18804 596134 19404 596218
rect 18804 595898 18986 596134
rect 19222 595898 19404 596134
rect 18804 560454 19404 595898
rect 18804 560218 18986 560454
rect 19222 560218 19404 560454
rect 18804 560134 19404 560218
rect 18804 559898 18986 560134
rect 19222 559898 19404 560134
rect 18804 524454 19404 559898
rect 18804 524218 18986 524454
rect 19222 524218 19404 524454
rect 18804 524134 19404 524218
rect 18804 523898 18986 524134
rect 19222 523898 19404 524134
rect 18804 488454 19404 523898
rect 18804 488218 18986 488454
rect 19222 488218 19404 488454
rect 18804 488134 19404 488218
rect 18804 487898 18986 488134
rect 19222 487898 19404 488134
rect 18804 452454 19404 487898
rect 18804 452218 18986 452454
rect 19222 452218 19404 452454
rect 18804 452134 19404 452218
rect 18804 451898 18986 452134
rect 19222 451898 19404 452134
rect 18804 416454 19404 451898
rect 18804 416218 18986 416454
rect 19222 416218 19404 416454
rect 18804 416134 19404 416218
rect 18804 415898 18986 416134
rect 19222 415898 19404 416134
rect 18804 380454 19404 415898
rect 18804 380218 18986 380454
rect 19222 380218 19404 380454
rect 18804 380134 19404 380218
rect 18804 379898 18986 380134
rect 19222 379898 19404 380134
rect 18804 344454 19404 379898
rect 18804 344218 18986 344454
rect 19222 344218 19404 344454
rect 18804 344134 19404 344218
rect 18804 343898 18986 344134
rect 19222 343898 19404 344134
rect 18804 308454 19404 343898
rect 18804 308218 18986 308454
rect 19222 308218 19404 308454
rect 18804 308134 19404 308218
rect 18804 307898 18986 308134
rect 19222 307898 19404 308134
rect 18804 272454 19404 307898
rect 18804 272218 18986 272454
rect 19222 272218 19404 272454
rect 18804 272134 19404 272218
rect 18804 271898 18986 272134
rect 19222 271898 19404 272134
rect 18804 236454 19404 271898
rect 18804 236218 18986 236454
rect 19222 236218 19404 236454
rect 18804 236134 19404 236218
rect 18804 235898 18986 236134
rect 19222 235898 19404 236134
rect 18804 200454 19404 235898
rect 18804 200218 18986 200454
rect 19222 200218 19404 200454
rect 18804 200134 19404 200218
rect 18804 199898 18986 200134
rect 19222 199898 19404 200134
rect 18804 164454 19404 199898
rect 18804 164218 18986 164454
rect 19222 164218 19404 164454
rect 18804 164134 19404 164218
rect 18804 163898 18986 164134
rect 19222 163898 19404 164134
rect 18804 128454 19404 163898
rect 18804 128218 18986 128454
rect 19222 128218 19404 128454
rect 18804 128134 19404 128218
rect 18804 127898 18986 128134
rect 19222 127898 19404 128134
rect 18804 92454 19404 127898
rect 18804 92218 18986 92454
rect 19222 92218 19404 92454
rect 18804 92134 19404 92218
rect 18804 91898 18986 92134
rect 19222 91898 19404 92134
rect 18804 56454 19404 91898
rect 18804 56218 18986 56454
rect 19222 56218 19404 56454
rect 18804 56134 19404 56218
rect 18804 55898 18986 56134
rect 19222 55898 19404 56134
rect 18804 20454 19404 55898
rect 18804 20218 18986 20454
rect 19222 20218 19404 20454
rect 18804 20134 19404 20218
rect 18804 19898 18986 20134
rect 19222 19898 19404 20134
rect 18804 -1266 19404 19898
rect 18804 -1502 18986 -1266
rect 19222 -1502 19404 -1266
rect 18804 -1586 19404 -1502
rect 18804 -1822 18986 -1586
rect 19222 -1822 19404 -1586
rect 18804 -1844 19404 -1822
rect 22404 672054 23004 707042
rect 22404 671818 22586 672054
rect 22822 671818 23004 672054
rect 22404 671734 23004 671818
rect 22404 671498 22586 671734
rect 22822 671498 23004 671734
rect 22404 636054 23004 671498
rect 22404 635818 22586 636054
rect 22822 635818 23004 636054
rect 22404 635734 23004 635818
rect 22404 635498 22586 635734
rect 22822 635498 23004 635734
rect 22404 600054 23004 635498
rect 22404 599818 22586 600054
rect 22822 599818 23004 600054
rect 22404 599734 23004 599818
rect 22404 599498 22586 599734
rect 22822 599498 23004 599734
rect 22404 564054 23004 599498
rect 22404 563818 22586 564054
rect 22822 563818 23004 564054
rect 22404 563734 23004 563818
rect 22404 563498 22586 563734
rect 22822 563498 23004 563734
rect 22404 528054 23004 563498
rect 22404 527818 22586 528054
rect 22822 527818 23004 528054
rect 22404 527734 23004 527818
rect 22404 527498 22586 527734
rect 22822 527498 23004 527734
rect 22404 492054 23004 527498
rect 22404 491818 22586 492054
rect 22822 491818 23004 492054
rect 22404 491734 23004 491818
rect 22404 491498 22586 491734
rect 22822 491498 23004 491734
rect 22404 456054 23004 491498
rect 22404 455818 22586 456054
rect 22822 455818 23004 456054
rect 22404 455734 23004 455818
rect 22404 455498 22586 455734
rect 22822 455498 23004 455734
rect 22404 420054 23004 455498
rect 22404 419818 22586 420054
rect 22822 419818 23004 420054
rect 22404 419734 23004 419818
rect 22404 419498 22586 419734
rect 22822 419498 23004 419734
rect 22404 384054 23004 419498
rect 22404 383818 22586 384054
rect 22822 383818 23004 384054
rect 22404 383734 23004 383818
rect 22404 383498 22586 383734
rect 22822 383498 23004 383734
rect 22404 348054 23004 383498
rect 22404 347818 22586 348054
rect 22822 347818 23004 348054
rect 22404 347734 23004 347818
rect 22404 347498 22586 347734
rect 22822 347498 23004 347734
rect 22404 312054 23004 347498
rect 22404 311818 22586 312054
rect 22822 311818 23004 312054
rect 22404 311734 23004 311818
rect 22404 311498 22586 311734
rect 22822 311498 23004 311734
rect 22404 276054 23004 311498
rect 22404 275818 22586 276054
rect 22822 275818 23004 276054
rect 22404 275734 23004 275818
rect 22404 275498 22586 275734
rect 22822 275498 23004 275734
rect 22404 240054 23004 275498
rect 22404 239818 22586 240054
rect 22822 239818 23004 240054
rect 22404 239734 23004 239818
rect 22404 239498 22586 239734
rect 22822 239498 23004 239734
rect 22404 204054 23004 239498
rect 22404 203818 22586 204054
rect 22822 203818 23004 204054
rect 22404 203734 23004 203818
rect 22404 203498 22586 203734
rect 22822 203498 23004 203734
rect 22404 168054 23004 203498
rect 22404 167818 22586 168054
rect 22822 167818 23004 168054
rect 22404 167734 23004 167818
rect 22404 167498 22586 167734
rect 22822 167498 23004 167734
rect 22404 132054 23004 167498
rect 22404 131818 22586 132054
rect 22822 131818 23004 132054
rect 22404 131734 23004 131818
rect 22404 131498 22586 131734
rect 22822 131498 23004 131734
rect 22404 96054 23004 131498
rect 22404 95818 22586 96054
rect 22822 95818 23004 96054
rect 22404 95734 23004 95818
rect 22404 95498 22586 95734
rect 22822 95498 23004 95734
rect 22404 60054 23004 95498
rect 22404 59818 22586 60054
rect 22822 59818 23004 60054
rect 22404 59734 23004 59818
rect 22404 59498 22586 59734
rect 22822 59498 23004 59734
rect 22404 24054 23004 59498
rect 22404 23818 22586 24054
rect 22822 23818 23004 24054
rect 22404 23734 23004 23818
rect 22404 23498 22586 23734
rect 22822 23498 23004 23734
rect 22404 -3106 23004 23498
rect 22404 -3342 22586 -3106
rect 22822 -3342 23004 -3106
rect 22404 -3426 23004 -3342
rect 22404 -3662 22586 -3426
rect 22822 -3662 23004 -3426
rect 22404 -3684 23004 -3662
rect 26004 675654 26604 708882
rect 26004 675418 26186 675654
rect 26422 675418 26604 675654
rect 26004 675334 26604 675418
rect 26004 675098 26186 675334
rect 26422 675098 26604 675334
rect 26004 639654 26604 675098
rect 26004 639418 26186 639654
rect 26422 639418 26604 639654
rect 26004 639334 26604 639418
rect 26004 639098 26186 639334
rect 26422 639098 26604 639334
rect 26004 603654 26604 639098
rect 26004 603418 26186 603654
rect 26422 603418 26604 603654
rect 26004 603334 26604 603418
rect 26004 603098 26186 603334
rect 26422 603098 26604 603334
rect 26004 567654 26604 603098
rect 26004 567418 26186 567654
rect 26422 567418 26604 567654
rect 26004 567334 26604 567418
rect 26004 567098 26186 567334
rect 26422 567098 26604 567334
rect 26004 531654 26604 567098
rect 26004 531418 26186 531654
rect 26422 531418 26604 531654
rect 26004 531334 26604 531418
rect 26004 531098 26186 531334
rect 26422 531098 26604 531334
rect 26004 495654 26604 531098
rect 26004 495418 26186 495654
rect 26422 495418 26604 495654
rect 26004 495334 26604 495418
rect 26004 495098 26186 495334
rect 26422 495098 26604 495334
rect 26004 459654 26604 495098
rect 26004 459418 26186 459654
rect 26422 459418 26604 459654
rect 26004 459334 26604 459418
rect 26004 459098 26186 459334
rect 26422 459098 26604 459334
rect 26004 423654 26604 459098
rect 26004 423418 26186 423654
rect 26422 423418 26604 423654
rect 26004 423334 26604 423418
rect 26004 423098 26186 423334
rect 26422 423098 26604 423334
rect 26004 387654 26604 423098
rect 26004 387418 26186 387654
rect 26422 387418 26604 387654
rect 26004 387334 26604 387418
rect 26004 387098 26186 387334
rect 26422 387098 26604 387334
rect 26004 351654 26604 387098
rect 26004 351418 26186 351654
rect 26422 351418 26604 351654
rect 26004 351334 26604 351418
rect 26004 351098 26186 351334
rect 26422 351098 26604 351334
rect 26004 315654 26604 351098
rect 26004 315418 26186 315654
rect 26422 315418 26604 315654
rect 26004 315334 26604 315418
rect 26004 315098 26186 315334
rect 26422 315098 26604 315334
rect 26004 279654 26604 315098
rect 26004 279418 26186 279654
rect 26422 279418 26604 279654
rect 26004 279334 26604 279418
rect 26004 279098 26186 279334
rect 26422 279098 26604 279334
rect 26004 243654 26604 279098
rect 26004 243418 26186 243654
rect 26422 243418 26604 243654
rect 26004 243334 26604 243418
rect 26004 243098 26186 243334
rect 26422 243098 26604 243334
rect 26004 207654 26604 243098
rect 26004 207418 26186 207654
rect 26422 207418 26604 207654
rect 26004 207334 26604 207418
rect 26004 207098 26186 207334
rect 26422 207098 26604 207334
rect 26004 171654 26604 207098
rect 26004 171418 26186 171654
rect 26422 171418 26604 171654
rect 26004 171334 26604 171418
rect 26004 171098 26186 171334
rect 26422 171098 26604 171334
rect 26004 135654 26604 171098
rect 26004 135418 26186 135654
rect 26422 135418 26604 135654
rect 26004 135334 26604 135418
rect 26004 135098 26186 135334
rect 26422 135098 26604 135334
rect 26004 99654 26604 135098
rect 26004 99418 26186 99654
rect 26422 99418 26604 99654
rect 26004 99334 26604 99418
rect 26004 99098 26186 99334
rect 26422 99098 26604 99334
rect 26004 63654 26604 99098
rect 26004 63418 26186 63654
rect 26422 63418 26604 63654
rect 26004 63334 26604 63418
rect 26004 63098 26186 63334
rect 26422 63098 26604 63334
rect 26004 27654 26604 63098
rect 26004 27418 26186 27654
rect 26422 27418 26604 27654
rect 26004 27334 26604 27418
rect 26004 27098 26186 27334
rect 26422 27098 26604 27334
rect 26004 -4946 26604 27098
rect 26004 -5182 26186 -4946
rect 26422 -5182 26604 -4946
rect 26004 -5266 26604 -5182
rect 26004 -5502 26186 -5266
rect 26422 -5502 26604 -5266
rect 26004 -5524 26604 -5502
rect 29604 679254 30204 710722
rect 47604 710358 48204 711300
rect 47604 710122 47786 710358
rect 48022 710122 48204 710358
rect 47604 710038 48204 710122
rect 47604 709802 47786 710038
rect 48022 709802 48204 710038
rect 44004 708518 44604 709460
rect 44004 708282 44186 708518
rect 44422 708282 44604 708518
rect 44004 708198 44604 708282
rect 44004 707962 44186 708198
rect 44422 707962 44604 708198
rect 40404 706678 41004 707620
rect 40404 706442 40586 706678
rect 40822 706442 41004 706678
rect 40404 706358 41004 706442
rect 40404 706122 40586 706358
rect 40822 706122 41004 706358
rect 29604 679018 29786 679254
rect 30022 679018 30204 679254
rect 29604 678934 30204 679018
rect 29604 678698 29786 678934
rect 30022 678698 30204 678934
rect 29604 643254 30204 678698
rect 29604 643018 29786 643254
rect 30022 643018 30204 643254
rect 29604 642934 30204 643018
rect 29604 642698 29786 642934
rect 30022 642698 30204 642934
rect 29604 607254 30204 642698
rect 29604 607018 29786 607254
rect 30022 607018 30204 607254
rect 29604 606934 30204 607018
rect 29604 606698 29786 606934
rect 30022 606698 30204 606934
rect 29604 571254 30204 606698
rect 29604 571018 29786 571254
rect 30022 571018 30204 571254
rect 29604 570934 30204 571018
rect 29604 570698 29786 570934
rect 30022 570698 30204 570934
rect 29604 535254 30204 570698
rect 29604 535018 29786 535254
rect 30022 535018 30204 535254
rect 29604 534934 30204 535018
rect 29604 534698 29786 534934
rect 30022 534698 30204 534934
rect 29604 499254 30204 534698
rect 29604 499018 29786 499254
rect 30022 499018 30204 499254
rect 29604 498934 30204 499018
rect 29604 498698 29786 498934
rect 30022 498698 30204 498934
rect 29604 463254 30204 498698
rect 29604 463018 29786 463254
rect 30022 463018 30204 463254
rect 29604 462934 30204 463018
rect 29604 462698 29786 462934
rect 30022 462698 30204 462934
rect 29604 427254 30204 462698
rect 29604 427018 29786 427254
rect 30022 427018 30204 427254
rect 29604 426934 30204 427018
rect 29604 426698 29786 426934
rect 30022 426698 30204 426934
rect 29604 391254 30204 426698
rect 29604 391018 29786 391254
rect 30022 391018 30204 391254
rect 29604 390934 30204 391018
rect 29604 390698 29786 390934
rect 30022 390698 30204 390934
rect 29604 355254 30204 390698
rect 29604 355018 29786 355254
rect 30022 355018 30204 355254
rect 29604 354934 30204 355018
rect 29604 354698 29786 354934
rect 30022 354698 30204 354934
rect 29604 319254 30204 354698
rect 29604 319018 29786 319254
rect 30022 319018 30204 319254
rect 29604 318934 30204 319018
rect 29604 318698 29786 318934
rect 30022 318698 30204 318934
rect 29604 283254 30204 318698
rect 29604 283018 29786 283254
rect 30022 283018 30204 283254
rect 29604 282934 30204 283018
rect 29604 282698 29786 282934
rect 30022 282698 30204 282934
rect 29604 247254 30204 282698
rect 29604 247018 29786 247254
rect 30022 247018 30204 247254
rect 29604 246934 30204 247018
rect 29604 246698 29786 246934
rect 30022 246698 30204 246934
rect 29604 211254 30204 246698
rect 29604 211018 29786 211254
rect 30022 211018 30204 211254
rect 29604 210934 30204 211018
rect 29604 210698 29786 210934
rect 30022 210698 30204 210934
rect 29604 175254 30204 210698
rect 29604 175018 29786 175254
rect 30022 175018 30204 175254
rect 29604 174934 30204 175018
rect 29604 174698 29786 174934
rect 30022 174698 30204 174934
rect 29604 139254 30204 174698
rect 29604 139018 29786 139254
rect 30022 139018 30204 139254
rect 29604 138934 30204 139018
rect 29604 138698 29786 138934
rect 30022 138698 30204 138934
rect 29604 103254 30204 138698
rect 29604 103018 29786 103254
rect 30022 103018 30204 103254
rect 29604 102934 30204 103018
rect 29604 102698 29786 102934
rect 30022 102698 30204 102934
rect 29604 67254 30204 102698
rect 29604 67018 29786 67254
rect 30022 67018 30204 67254
rect 29604 66934 30204 67018
rect 29604 66698 29786 66934
rect 30022 66698 30204 66934
rect 29604 31254 30204 66698
rect 29604 31018 29786 31254
rect 30022 31018 30204 31254
rect 29604 30934 30204 31018
rect 29604 30698 29786 30934
rect 30022 30698 30204 30934
rect 11604 -6102 11786 -5866
rect 12022 -6102 12204 -5866
rect 11604 -6186 12204 -6102
rect 11604 -6422 11786 -6186
rect 12022 -6422 12204 -6186
rect -8436 -7022 -8254 -6786
rect -8018 -7022 -7836 -6786
rect -8436 -7106 -7836 -7022
rect -8436 -7342 -8254 -7106
rect -8018 -7342 -7836 -7106
rect -8436 -7364 -7836 -7342
rect 11604 -7364 12204 -6422
rect 29604 -6786 30204 30698
rect 36804 704838 37404 705780
rect 36804 704602 36986 704838
rect 37222 704602 37404 704838
rect 36804 704518 37404 704602
rect 36804 704282 36986 704518
rect 37222 704282 37404 704518
rect 36804 686454 37404 704282
rect 36804 686218 36986 686454
rect 37222 686218 37404 686454
rect 36804 686134 37404 686218
rect 36804 685898 36986 686134
rect 37222 685898 37404 686134
rect 36804 650454 37404 685898
rect 36804 650218 36986 650454
rect 37222 650218 37404 650454
rect 36804 650134 37404 650218
rect 36804 649898 36986 650134
rect 37222 649898 37404 650134
rect 36804 614454 37404 649898
rect 36804 614218 36986 614454
rect 37222 614218 37404 614454
rect 36804 614134 37404 614218
rect 36804 613898 36986 614134
rect 37222 613898 37404 614134
rect 36804 578454 37404 613898
rect 36804 578218 36986 578454
rect 37222 578218 37404 578454
rect 36804 578134 37404 578218
rect 36804 577898 36986 578134
rect 37222 577898 37404 578134
rect 36804 542454 37404 577898
rect 36804 542218 36986 542454
rect 37222 542218 37404 542454
rect 36804 542134 37404 542218
rect 36804 541898 36986 542134
rect 37222 541898 37404 542134
rect 36804 506454 37404 541898
rect 36804 506218 36986 506454
rect 37222 506218 37404 506454
rect 36804 506134 37404 506218
rect 36804 505898 36986 506134
rect 37222 505898 37404 506134
rect 36804 470454 37404 505898
rect 36804 470218 36986 470454
rect 37222 470218 37404 470454
rect 36804 470134 37404 470218
rect 36804 469898 36986 470134
rect 37222 469898 37404 470134
rect 36804 434454 37404 469898
rect 36804 434218 36986 434454
rect 37222 434218 37404 434454
rect 36804 434134 37404 434218
rect 36804 433898 36986 434134
rect 37222 433898 37404 434134
rect 36804 398454 37404 433898
rect 36804 398218 36986 398454
rect 37222 398218 37404 398454
rect 36804 398134 37404 398218
rect 36804 397898 36986 398134
rect 37222 397898 37404 398134
rect 36804 362454 37404 397898
rect 36804 362218 36986 362454
rect 37222 362218 37404 362454
rect 36804 362134 37404 362218
rect 36804 361898 36986 362134
rect 37222 361898 37404 362134
rect 36804 326454 37404 361898
rect 36804 326218 36986 326454
rect 37222 326218 37404 326454
rect 36804 326134 37404 326218
rect 36804 325898 36986 326134
rect 37222 325898 37404 326134
rect 36804 290454 37404 325898
rect 36804 290218 36986 290454
rect 37222 290218 37404 290454
rect 36804 290134 37404 290218
rect 36804 289898 36986 290134
rect 37222 289898 37404 290134
rect 36804 254454 37404 289898
rect 36804 254218 36986 254454
rect 37222 254218 37404 254454
rect 36804 254134 37404 254218
rect 36804 253898 36986 254134
rect 37222 253898 37404 254134
rect 36804 218454 37404 253898
rect 36804 218218 36986 218454
rect 37222 218218 37404 218454
rect 36804 218134 37404 218218
rect 36804 217898 36986 218134
rect 37222 217898 37404 218134
rect 36804 182454 37404 217898
rect 36804 182218 36986 182454
rect 37222 182218 37404 182454
rect 36804 182134 37404 182218
rect 36804 181898 36986 182134
rect 37222 181898 37404 182134
rect 36804 146454 37404 181898
rect 36804 146218 36986 146454
rect 37222 146218 37404 146454
rect 36804 146134 37404 146218
rect 36804 145898 36986 146134
rect 37222 145898 37404 146134
rect 36804 110454 37404 145898
rect 36804 110218 36986 110454
rect 37222 110218 37404 110454
rect 36804 110134 37404 110218
rect 36804 109898 36986 110134
rect 37222 109898 37404 110134
rect 36804 74454 37404 109898
rect 36804 74218 36986 74454
rect 37222 74218 37404 74454
rect 36804 74134 37404 74218
rect 36804 73898 36986 74134
rect 37222 73898 37404 74134
rect 36804 38454 37404 73898
rect 36804 38218 36986 38454
rect 37222 38218 37404 38454
rect 36804 38134 37404 38218
rect 36804 37898 36986 38134
rect 37222 37898 37404 38134
rect 36804 2454 37404 37898
rect 36804 2218 36986 2454
rect 37222 2218 37404 2454
rect 36804 2134 37404 2218
rect 36804 1898 36986 2134
rect 37222 1898 37404 2134
rect 36804 -346 37404 1898
rect 36804 -582 36986 -346
rect 37222 -582 37404 -346
rect 36804 -666 37404 -582
rect 36804 -902 36986 -666
rect 37222 -902 37404 -666
rect 36804 -1844 37404 -902
rect 40404 690054 41004 706122
rect 40404 689818 40586 690054
rect 40822 689818 41004 690054
rect 40404 689734 41004 689818
rect 40404 689498 40586 689734
rect 40822 689498 41004 689734
rect 40404 654054 41004 689498
rect 40404 653818 40586 654054
rect 40822 653818 41004 654054
rect 40404 653734 41004 653818
rect 40404 653498 40586 653734
rect 40822 653498 41004 653734
rect 40404 618054 41004 653498
rect 40404 617818 40586 618054
rect 40822 617818 41004 618054
rect 40404 617734 41004 617818
rect 40404 617498 40586 617734
rect 40822 617498 41004 617734
rect 40404 582054 41004 617498
rect 40404 581818 40586 582054
rect 40822 581818 41004 582054
rect 40404 581734 41004 581818
rect 40404 581498 40586 581734
rect 40822 581498 41004 581734
rect 40404 546054 41004 581498
rect 40404 545818 40586 546054
rect 40822 545818 41004 546054
rect 40404 545734 41004 545818
rect 40404 545498 40586 545734
rect 40822 545498 41004 545734
rect 40404 510054 41004 545498
rect 40404 509818 40586 510054
rect 40822 509818 41004 510054
rect 40404 509734 41004 509818
rect 40404 509498 40586 509734
rect 40822 509498 41004 509734
rect 40404 474054 41004 509498
rect 40404 473818 40586 474054
rect 40822 473818 41004 474054
rect 40404 473734 41004 473818
rect 40404 473498 40586 473734
rect 40822 473498 41004 473734
rect 40404 438054 41004 473498
rect 40404 437818 40586 438054
rect 40822 437818 41004 438054
rect 40404 437734 41004 437818
rect 40404 437498 40586 437734
rect 40822 437498 41004 437734
rect 40404 402054 41004 437498
rect 40404 401818 40586 402054
rect 40822 401818 41004 402054
rect 40404 401734 41004 401818
rect 40404 401498 40586 401734
rect 40822 401498 41004 401734
rect 40404 366054 41004 401498
rect 40404 365818 40586 366054
rect 40822 365818 41004 366054
rect 40404 365734 41004 365818
rect 40404 365498 40586 365734
rect 40822 365498 41004 365734
rect 40404 330054 41004 365498
rect 40404 329818 40586 330054
rect 40822 329818 41004 330054
rect 40404 329734 41004 329818
rect 40404 329498 40586 329734
rect 40822 329498 41004 329734
rect 40404 294054 41004 329498
rect 40404 293818 40586 294054
rect 40822 293818 41004 294054
rect 40404 293734 41004 293818
rect 40404 293498 40586 293734
rect 40822 293498 41004 293734
rect 40404 258054 41004 293498
rect 40404 257818 40586 258054
rect 40822 257818 41004 258054
rect 40404 257734 41004 257818
rect 40404 257498 40586 257734
rect 40822 257498 41004 257734
rect 40404 222054 41004 257498
rect 40404 221818 40586 222054
rect 40822 221818 41004 222054
rect 40404 221734 41004 221818
rect 40404 221498 40586 221734
rect 40822 221498 41004 221734
rect 40404 186054 41004 221498
rect 40404 185818 40586 186054
rect 40822 185818 41004 186054
rect 40404 185734 41004 185818
rect 40404 185498 40586 185734
rect 40822 185498 41004 185734
rect 40404 150054 41004 185498
rect 40404 149818 40586 150054
rect 40822 149818 41004 150054
rect 40404 149734 41004 149818
rect 40404 149498 40586 149734
rect 40822 149498 41004 149734
rect 40404 114054 41004 149498
rect 40404 113818 40586 114054
rect 40822 113818 41004 114054
rect 40404 113734 41004 113818
rect 40404 113498 40586 113734
rect 40822 113498 41004 113734
rect 40404 78054 41004 113498
rect 40404 77818 40586 78054
rect 40822 77818 41004 78054
rect 40404 77734 41004 77818
rect 40404 77498 40586 77734
rect 40822 77498 41004 77734
rect 40404 42054 41004 77498
rect 40404 41818 40586 42054
rect 40822 41818 41004 42054
rect 40404 41734 41004 41818
rect 40404 41498 40586 41734
rect 40822 41498 41004 41734
rect 40404 6054 41004 41498
rect 40404 5818 40586 6054
rect 40822 5818 41004 6054
rect 40404 5734 41004 5818
rect 40404 5498 40586 5734
rect 40822 5498 41004 5734
rect 40404 -2186 41004 5498
rect 40404 -2422 40586 -2186
rect 40822 -2422 41004 -2186
rect 40404 -2506 41004 -2422
rect 40404 -2742 40586 -2506
rect 40822 -2742 41004 -2506
rect 40404 -3684 41004 -2742
rect 44004 693654 44604 707962
rect 44004 693418 44186 693654
rect 44422 693418 44604 693654
rect 44004 693334 44604 693418
rect 44004 693098 44186 693334
rect 44422 693098 44604 693334
rect 44004 657654 44604 693098
rect 44004 657418 44186 657654
rect 44422 657418 44604 657654
rect 44004 657334 44604 657418
rect 44004 657098 44186 657334
rect 44422 657098 44604 657334
rect 44004 621654 44604 657098
rect 44004 621418 44186 621654
rect 44422 621418 44604 621654
rect 44004 621334 44604 621418
rect 44004 621098 44186 621334
rect 44422 621098 44604 621334
rect 44004 585654 44604 621098
rect 44004 585418 44186 585654
rect 44422 585418 44604 585654
rect 44004 585334 44604 585418
rect 44004 585098 44186 585334
rect 44422 585098 44604 585334
rect 44004 549654 44604 585098
rect 44004 549418 44186 549654
rect 44422 549418 44604 549654
rect 44004 549334 44604 549418
rect 44004 549098 44186 549334
rect 44422 549098 44604 549334
rect 44004 513654 44604 549098
rect 44004 513418 44186 513654
rect 44422 513418 44604 513654
rect 44004 513334 44604 513418
rect 44004 513098 44186 513334
rect 44422 513098 44604 513334
rect 44004 477654 44604 513098
rect 44004 477418 44186 477654
rect 44422 477418 44604 477654
rect 44004 477334 44604 477418
rect 44004 477098 44186 477334
rect 44422 477098 44604 477334
rect 44004 441654 44604 477098
rect 44004 441418 44186 441654
rect 44422 441418 44604 441654
rect 44004 441334 44604 441418
rect 44004 441098 44186 441334
rect 44422 441098 44604 441334
rect 44004 405654 44604 441098
rect 44004 405418 44186 405654
rect 44422 405418 44604 405654
rect 44004 405334 44604 405418
rect 44004 405098 44186 405334
rect 44422 405098 44604 405334
rect 44004 369654 44604 405098
rect 44004 369418 44186 369654
rect 44422 369418 44604 369654
rect 44004 369334 44604 369418
rect 44004 369098 44186 369334
rect 44422 369098 44604 369334
rect 44004 333654 44604 369098
rect 44004 333418 44186 333654
rect 44422 333418 44604 333654
rect 44004 333334 44604 333418
rect 44004 333098 44186 333334
rect 44422 333098 44604 333334
rect 44004 297654 44604 333098
rect 44004 297418 44186 297654
rect 44422 297418 44604 297654
rect 44004 297334 44604 297418
rect 44004 297098 44186 297334
rect 44422 297098 44604 297334
rect 44004 261654 44604 297098
rect 44004 261418 44186 261654
rect 44422 261418 44604 261654
rect 44004 261334 44604 261418
rect 44004 261098 44186 261334
rect 44422 261098 44604 261334
rect 44004 225654 44604 261098
rect 44004 225418 44186 225654
rect 44422 225418 44604 225654
rect 44004 225334 44604 225418
rect 44004 225098 44186 225334
rect 44422 225098 44604 225334
rect 44004 189654 44604 225098
rect 44004 189418 44186 189654
rect 44422 189418 44604 189654
rect 44004 189334 44604 189418
rect 44004 189098 44186 189334
rect 44422 189098 44604 189334
rect 44004 153654 44604 189098
rect 44004 153418 44186 153654
rect 44422 153418 44604 153654
rect 44004 153334 44604 153418
rect 44004 153098 44186 153334
rect 44422 153098 44604 153334
rect 44004 117654 44604 153098
rect 44004 117418 44186 117654
rect 44422 117418 44604 117654
rect 44004 117334 44604 117418
rect 44004 117098 44186 117334
rect 44422 117098 44604 117334
rect 44004 81654 44604 117098
rect 44004 81418 44186 81654
rect 44422 81418 44604 81654
rect 44004 81334 44604 81418
rect 44004 81098 44186 81334
rect 44422 81098 44604 81334
rect 44004 45654 44604 81098
rect 44004 45418 44186 45654
rect 44422 45418 44604 45654
rect 44004 45334 44604 45418
rect 44004 45098 44186 45334
rect 44422 45098 44604 45334
rect 44004 9654 44604 45098
rect 44004 9418 44186 9654
rect 44422 9418 44604 9654
rect 44004 9334 44604 9418
rect 44004 9098 44186 9334
rect 44422 9098 44604 9334
rect 44004 -4026 44604 9098
rect 44004 -4262 44186 -4026
rect 44422 -4262 44604 -4026
rect 44004 -4346 44604 -4262
rect 44004 -4582 44186 -4346
rect 44422 -4582 44604 -4346
rect 44004 -5524 44604 -4582
rect 47604 697254 48204 709802
rect 65604 711278 66204 711300
rect 65604 711042 65786 711278
rect 66022 711042 66204 711278
rect 65604 710958 66204 711042
rect 65604 710722 65786 710958
rect 66022 710722 66204 710958
rect 62004 709438 62604 709460
rect 62004 709202 62186 709438
rect 62422 709202 62604 709438
rect 62004 709118 62604 709202
rect 62004 708882 62186 709118
rect 62422 708882 62604 709118
rect 58404 707598 59004 707620
rect 58404 707362 58586 707598
rect 58822 707362 59004 707598
rect 58404 707278 59004 707362
rect 58404 707042 58586 707278
rect 58822 707042 59004 707278
rect 47604 697018 47786 697254
rect 48022 697018 48204 697254
rect 47604 696934 48204 697018
rect 47604 696698 47786 696934
rect 48022 696698 48204 696934
rect 47604 661254 48204 696698
rect 47604 661018 47786 661254
rect 48022 661018 48204 661254
rect 47604 660934 48204 661018
rect 47604 660698 47786 660934
rect 48022 660698 48204 660934
rect 47604 625254 48204 660698
rect 47604 625018 47786 625254
rect 48022 625018 48204 625254
rect 47604 624934 48204 625018
rect 47604 624698 47786 624934
rect 48022 624698 48204 624934
rect 47604 589254 48204 624698
rect 47604 589018 47786 589254
rect 48022 589018 48204 589254
rect 47604 588934 48204 589018
rect 47604 588698 47786 588934
rect 48022 588698 48204 588934
rect 47604 553254 48204 588698
rect 47604 553018 47786 553254
rect 48022 553018 48204 553254
rect 47604 552934 48204 553018
rect 47604 552698 47786 552934
rect 48022 552698 48204 552934
rect 47604 517254 48204 552698
rect 47604 517018 47786 517254
rect 48022 517018 48204 517254
rect 47604 516934 48204 517018
rect 47604 516698 47786 516934
rect 48022 516698 48204 516934
rect 47604 481254 48204 516698
rect 47604 481018 47786 481254
rect 48022 481018 48204 481254
rect 47604 480934 48204 481018
rect 47604 480698 47786 480934
rect 48022 480698 48204 480934
rect 47604 445254 48204 480698
rect 47604 445018 47786 445254
rect 48022 445018 48204 445254
rect 47604 444934 48204 445018
rect 47604 444698 47786 444934
rect 48022 444698 48204 444934
rect 47604 409254 48204 444698
rect 47604 409018 47786 409254
rect 48022 409018 48204 409254
rect 47604 408934 48204 409018
rect 47604 408698 47786 408934
rect 48022 408698 48204 408934
rect 47604 373254 48204 408698
rect 47604 373018 47786 373254
rect 48022 373018 48204 373254
rect 47604 372934 48204 373018
rect 47604 372698 47786 372934
rect 48022 372698 48204 372934
rect 47604 337254 48204 372698
rect 47604 337018 47786 337254
rect 48022 337018 48204 337254
rect 47604 336934 48204 337018
rect 47604 336698 47786 336934
rect 48022 336698 48204 336934
rect 47604 301254 48204 336698
rect 47604 301018 47786 301254
rect 48022 301018 48204 301254
rect 47604 300934 48204 301018
rect 47604 300698 47786 300934
rect 48022 300698 48204 300934
rect 47604 265254 48204 300698
rect 47604 265018 47786 265254
rect 48022 265018 48204 265254
rect 47604 264934 48204 265018
rect 47604 264698 47786 264934
rect 48022 264698 48204 264934
rect 47604 229254 48204 264698
rect 47604 229018 47786 229254
rect 48022 229018 48204 229254
rect 47604 228934 48204 229018
rect 47604 228698 47786 228934
rect 48022 228698 48204 228934
rect 47604 193254 48204 228698
rect 47604 193018 47786 193254
rect 48022 193018 48204 193254
rect 47604 192934 48204 193018
rect 47604 192698 47786 192934
rect 48022 192698 48204 192934
rect 47604 157254 48204 192698
rect 47604 157018 47786 157254
rect 48022 157018 48204 157254
rect 47604 156934 48204 157018
rect 47604 156698 47786 156934
rect 48022 156698 48204 156934
rect 47604 121254 48204 156698
rect 47604 121018 47786 121254
rect 48022 121018 48204 121254
rect 47604 120934 48204 121018
rect 47604 120698 47786 120934
rect 48022 120698 48204 120934
rect 47604 85254 48204 120698
rect 47604 85018 47786 85254
rect 48022 85018 48204 85254
rect 47604 84934 48204 85018
rect 47604 84698 47786 84934
rect 48022 84698 48204 84934
rect 47604 49254 48204 84698
rect 47604 49018 47786 49254
rect 48022 49018 48204 49254
rect 47604 48934 48204 49018
rect 47604 48698 47786 48934
rect 48022 48698 48204 48934
rect 47604 13254 48204 48698
rect 47604 13018 47786 13254
rect 48022 13018 48204 13254
rect 47604 12934 48204 13018
rect 47604 12698 47786 12934
rect 48022 12698 48204 12934
rect 29604 -7022 29786 -6786
rect 30022 -7022 30204 -6786
rect 29604 -7106 30204 -7022
rect 29604 -7342 29786 -7106
rect 30022 -7342 30204 -7106
rect 29604 -7364 30204 -7342
rect 47604 -5866 48204 12698
rect 54804 705758 55404 705780
rect 54804 705522 54986 705758
rect 55222 705522 55404 705758
rect 54804 705438 55404 705522
rect 54804 705202 54986 705438
rect 55222 705202 55404 705438
rect 54804 668454 55404 705202
rect 54804 668218 54986 668454
rect 55222 668218 55404 668454
rect 54804 668134 55404 668218
rect 54804 667898 54986 668134
rect 55222 667898 55404 668134
rect 54804 632454 55404 667898
rect 54804 632218 54986 632454
rect 55222 632218 55404 632454
rect 54804 632134 55404 632218
rect 54804 631898 54986 632134
rect 55222 631898 55404 632134
rect 54804 596454 55404 631898
rect 54804 596218 54986 596454
rect 55222 596218 55404 596454
rect 54804 596134 55404 596218
rect 54804 595898 54986 596134
rect 55222 595898 55404 596134
rect 54804 560454 55404 595898
rect 54804 560218 54986 560454
rect 55222 560218 55404 560454
rect 54804 560134 55404 560218
rect 54804 559898 54986 560134
rect 55222 559898 55404 560134
rect 54804 524454 55404 559898
rect 54804 524218 54986 524454
rect 55222 524218 55404 524454
rect 54804 524134 55404 524218
rect 54804 523898 54986 524134
rect 55222 523898 55404 524134
rect 54804 488454 55404 523898
rect 54804 488218 54986 488454
rect 55222 488218 55404 488454
rect 54804 488134 55404 488218
rect 54804 487898 54986 488134
rect 55222 487898 55404 488134
rect 54804 452454 55404 487898
rect 54804 452218 54986 452454
rect 55222 452218 55404 452454
rect 54804 452134 55404 452218
rect 54804 451898 54986 452134
rect 55222 451898 55404 452134
rect 54804 416454 55404 451898
rect 54804 416218 54986 416454
rect 55222 416218 55404 416454
rect 54804 416134 55404 416218
rect 54804 415898 54986 416134
rect 55222 415898 55404 416134
rect 54804 380454 55404 415898
rect 54804 380218 54986 380454
rect 55222 380218 55404 380454
rect 54804 380134 55404 380218
rect 54804 379898 54986 380134
rect 55222 379898 55404 380134
rect 54804 344454 55404 379898
rect 54804 344218 54986 344454
rect 55222 344218 55404 344454
rect 54804 344134 55404 344218
rect 54804 343898 54986 344134
rect 55222 343898 55404 344134
rect 54804 308454 55404 343898
rect 54804 308218 54986 308454
rect 55222 308218 55404 308454
rect 54804 308134 55404 308218
rect 54804 307898 54986 308134
rect 55222 307898 55404 308134
rect 54804 272454 55404 307898
rect 54804 272218 54986 272454
rect 55222 272218 55404 272454
rect 54804 272134 55404 272218
rect 54804 271898 54986 272134
rect 55222 271898 55404 272134
rect 54804 236454 55404 271898
rect 54804 236218 54986 236454
rect 55222 236218 55404 236454
rect 54804 236134 55404 236218
rect 54804 235898 54986 236134
rect 55222 235898 55404 236134
rect 54804 200454 55404 235898
rect 54804 200218 54986 200454
rect 55222 200218 55404 200454
rect 54804 200134 55404 200218
rect 54804 199898 54986 200134
rect 55222 199898 55404 200134
rect 54804 164454 55404 199898
rect 54804 164218 54986 164454
rect 55222 164218 55404 164454
rect 54804 164134 55404 164218
rect 54804 163898 54986 164134
rect 55222 163898 55404 164134
rect 54804 128454 55404 163898
rect 54804 128218 54986 128454
rect 55222 128218 55404 128454
rect 54804 128134 55404 128218
rect 54804 127898 54986 128134
rect 55222 127898 55404 128134
rect 54804 92454 55404 127898
rect 54804 92218 54986 92454
rect 55222 92218 55404 92454
rect 54804 92134 55404 92218
rect 54804 91898 54986 92134
rect 55222 91898 55404 92134
rect 54804 56454 55404 91898
rect 54804 56218 54986 56454
rect 55222 56218 55404 56454
rect 54804 56134 55404 56218
rect 54804 55898 54986 56134
rect 55222 55898 55404 56134
rect 54804 20454 55404 55898
rect 54804 20218 54986 20454
rect 55222 20218 55404 20454
rect 54804 20134 55404 20218
rect 54804 19898 54986 20134
rect 55222 19898 55404 20134
rect 54804 -1266 55404 19898
rect 54804 -1502 54986 -1266
rect 55222 -1502 55404 -1266
rect 54804 -1586 55404 -1502
rect 54804 -1822 54986 -1586
rect 55222 -1822 55404 -1586
rect 54804 -1844 55404 -1822
rect 58404 672054 59004 707042
rect 58404 671818 58586 672054
rect 58822 671818 59004 672054
rect 58404 671734 59004 671818
rect 58404 671498 58586 671734
rect 58822 671498 59004 671734
rect 58404 636054 59004 671498
rect 58404 635818 58586 636054
rect 58822 635818 59004 636054
rect 58404 635734 59004 635818
rect 58404 635498 58586 635734
rect 58822 635498 59004 635734
rect 58404 600054 59004 635498
rect 58404 599818 58586 600054
rect 58822 599818 59004 600054
rect 58404 599734 59004 599818
rect 58404 599498 58586 599734
rect 58822 599498 59004 599734
rect 58404 564054 59004 599498
rect 58404 563818 58586 564054
rect 58822 563818 59004 564054
rect 58404 563734 59004 563818
rect 58404 563498 58586 563734
rect 58822 563498 59004 563734
rect 58404 528054 59004 563498
rect 58404 527818 58586 528054
rect 58822 527818 59004 528054
rect 58404 527734 59004 527818
rect 58404 527498 58586 527734
rect 58822 527498 59004 527734
rect 58404 492054 59004 527498
rect 58404 491818 58586 492054
rect 58822 491818 59004 492054
rect 58404 491734 59004 491818
rect 58404 491498 58586 491734
rect 58822 491498 59004 491734
rect 58404 456054 59004 491498
rect 58404 455818 58586 456054
rect 58822 455818 59004 456054
rect 58404 455734 59004 455818
rect 58404 455498 58586 455734
rect 58822 455498 59004 455734
rect 58404 420054 59004 455498
rect 58404 419818 58586 420054
rect 58822 419818 59004 420054
rect 58404 419734 59004 419818
rect 58404 419498 58586 419734
rect 58822 419498 59004 419734
rect 58404 384054 59004 419498
rect 58404 383818 58586 384054
rect 58822 383818 59004 384054
rect 58404 383734 59004 383818
rect 58404 383498 58586 383734
rect 58822 383498 59004 383734
rect 58404 348054 59004 383498
rect 58404 347818 58586 348054
rect 58822 347818 59004 348054
rect 58404 347734 59004 347818
rect 58404 347498 58586 347734
rect 58822 347498 59004 347734
rect 58404 312054 59004 347498
rect 58404 311818 58586 312054
rect 58822 311818 59004 312054
rect 58404 311734 59004 311818
rect 58404 311498 58586 311734
rect 58822 311498 59004 311734
rect 58404 276054 59004 311498
rect 58404 275818 58586 276054
rect 58822 275818 59004 276054
rect 58404 275734 59004 275818
rect 58404 275498 58586 275734
rect 58822 275498 59004 275734
rect 58404 240054 59004 275498
rect 58404 239818 58586 240054
rect 58822 239818 59004 240054
rect 58404 239734 59004 239818
rect 58404 239498 58586 239734
rect 58822 239498 59004 239734
rect 58404 204054 59004 239498
rect 58404 203818 58586 204054
rect 58822 203818 59004 204054
rect 58404 203734 59004 203818
rect 58404 203498 58586 203734
rect 58822 203498 59004 203734
rect 58404 168054 59004 203498
rect 58404 167818 58586 168054
rect 58822 167818 59004 168054
rect 58404 167734 59004 167818
rect 58404 167498 58586 167734
rect 58822 167498 59004 167734
rect 58404 132054 59004 167498
rect 58404 131818 58586 132054
rect 58822 131818 59004 132054
rect 58404 131734 59004 131818
rect 58404 131498 58586 131734
rect 58822 131498 59004 131734
rect 58404 96054 59004 131498
rect 58404 95818 58586 96054
rect 58822 95818 59004 96054
rect 58404 95734 59004 95818
rect 58404 95498 58586 95734
rect 58822 95498 59004 95734
rect 58404 60054 59004 95498
rect 58404 59818 58586 60054
rect 58822 59818 59004 60054
rect 58404 59734 59004 59818
rect 58404 59498 58586 59734
rect 58822 59498 59004 59734
rect 58404 24054 59004 59498
rect 58404 23818 58586 24054
rect 58822 23818 59004 24054
rect 58404 23734 59004 23818
rect 58404 23498 58586 23734
rect 58822 23498 59004 23734
rect 58404 -3106 59004 23498
rect 58404 -3342 58586 -3106
rect 58822 -3342 59004 -3106
rect 58404 -3426 59004 -3342
rect 58404 -3662 58586 -3426
rect 58822 -3662 59004 -3426
rect 58404 -3684 59004 -3662
rect 62004 675654 62604 708882
rect 62004 675418 62186 675654
rect 62422 675418 62604 675654
rect 62004 675334 62604 675418
rect 62004 675098 62186 675334
rect 62422 675098 62604 675334
rect 62004 639654 62604 675098
rect 62004 639418 62186 639654
rect 62422 639418 62604 639654
rect 62004 639334 62604 639418
rect 62004 639098 62186 639334
rect 62422 639098 62604 639334
rect 62004 603654 62604 639098
rect 62004 603418 62186 603654
rect 62422 603418 62604 603654
rect 62004 603334 62604 603418
rect 62004 603098 62186 603334
rect 62422 603098 62604 603334
rect 62004 567654 62604 603098
rect 62004 567418 62186 567654
rect 62422 567418 62604 567654
rect 62004 567334 62604 567418
rect 62004 567098 62186 567334
rect 62422 567098 62604 567334
rect 62004 531654 62604 567098
rect 62004 531418 62186 531654
rect 62422 531418 62604 531654
rect 62004 531334 62604 531418
rect 62004 531098 62186 531334
rect 62422 531098 62604 531334
rect 62004 495654 62604 531098
rect 62004 495418 62186 495654
rect 62422 495418 62604 495654
rect 62004 495334 62604 495418
rect 62004 495098 62186 495334
rect 62422 495098 62604 495334
rect 62004 459654 62604 495098
rect 62004 459418 62186 459654
rect 62422 459418 62604 459654
rect 62004 459334 62604 459418
rect 62004 459098 62186 459334
rect 62422 459098 62604 459334
rect 62004 423654 62604 459098
rect 62004 423418 62186 423654
rect 62422 423418 62604 423654
rect 62004 423334 62604 423418
rect 62004 423098 62186 423334
rect 62422 423098 62604 423334
rect 62004 387654 62604 423098
rect 62004 387418 62186 387654
rect 62422 387418 62604 387654
rect 62004 387334 62604 387418
rect 62004 387098 62186 387334
rect 62422 387098 62604 387334
rect 62004 351654 62604 387098
rect 62004 351418 62186 351654
rect 62422 351418 62604 351654
rect 62004 351334 62604 351418
rect 62004 351098 62186 351334
rect 62422 351098 62604 351334
rect 62004 315654 62604 351098
rect 62004 315418 62186 315654
rect 62422 315418 62604 315654
rect 62004 315334 62604 315418
rect 62004 315098 62186 315334
rect 62422 315098 62604 315334
rect 62004 279654 62604 315098
rect 62004 279418 62186 279654
rect 62422 279418 62604 279654
rect 62004 279334 62604 279418
rect 62004 279098 62186 279334
rect 62422 279098 62604 279334
rect 62004 243654 62604 279098
rect 62004 243418 62186 243654
rect 62422 243418 62604 243654
rect 62004 243334 62604 243418
rect 62004 243098 62186 243334
rect 62422 243098 62604 243334
rect 62004 207654 62604 243098
rect 62004 207418 62186 207654
rect 62422 207418 62604 207654
rect 62004 207334 62604 207418
rect 62004 207098 62186 207334
rect 62422 207098 62604 207334
rect 62004 171654 62604 207098
rect 62004 171418 62186 171654
rect 62422 171418 62604 171654
rect 62004 171334 62604 171418
rect 62004 171098 62186 171334
rect 62422 171098 62604 171334
rect 62004 135654 62604 171098
rect 62004 135418 62186 135654
rect 62422 135418 62604 135654
rect 62004 135334 62604 135418
rect 62004 135098 62186 135334
rect 62422 135098 62604 135334
rect 62004 99654 62604 135098
rect 62004 99418 62186 99654
rect 62422 99418 62604 99654
rect 62004 99334 62604 99418
rect 62004 99098 62186 99334
rect 62422 99098 62604 99334
rect 62004 63654 62604 99098
rect 62004 63418 62186 63654
rect 62422 63418 62604 63654
rect 62004 63334 62604 63418
rect 62004 63098 62186 63334
rect 62422 63098 62604 63334
rect 62004 27654 62604 63098
rect 62004 27418 62186 27654
rect 62422 27418 62604 27654
rect 62004 27334 62604 27418
rect 62004 27098 62186 27334
rect 62422 27098 62604 27334
rect 62004 -4946 62604 27098
rect 62004 -5182 62186 -4946
rect 62422 -5182 62604 -4946
rect 62004 -5266 62604 -5182
rect 62004 -5502 62186 -5266
rect 62422 -5502 62604 -5266
rect 62004 -5524 62604 -5502
rect 65604 679254 66204 710722
rect 83604 710358 84204 711300
rect 83604 710122 83786 710358
rect 84022 710122 84204 710358
rect 83604 710038 84204 710122
rect 83604 709802 83786 710038
rect 84022 709802 84204 710038
rect 80004 708518 80604 709460
rect 80004 708282 80186 708518
rect 80422 708282 80604 708518
rect 80004 708198 80604 708282
rect 80004 707962 80186 708198
rect 80422 707962 80604 708198
rect 76404 706678 77004 707620
rect 76404 706442 76586 706678
rect 76822 706442 77004 706678
rect 76404 706358 77004 706442
rect 76404 706122 76586 706358
rect 76822 706122 77004 706358
rect 65604 679018 65786 679254
rect 66022 679018 66204 679254
rect 65604 678934 66204 679018
rect 65604 678698 65786 678934
rect 66022 678698 66204 678934
rect 65604 643254 66204 678698
rect 65604 643018 65786 643254
rect 66022 643018 66204 643254
rect 65604 642934 66204 643018
rect 65604 642698 65786 642934
rect 66022 642698 66204 642934
rect 65604 607254 66204 642698
rect 65604 607018 65786 607254
rect 66022 607018 66204 607254
rect 65604 606934 66204 607018
rect 65604 606698 65786 606934
rect 66022 606698 66204 606934
rect 65604 571254 66204 606698
rect 65604 571018 65786 571254
rect 66022 571018 66204 571254
rect 65604 570934 66204 571018
rect 65604 570698 65786 570934
rect 66022 570698 66204 570934
rect 65604 535254 66204 570698
rect 65604 535018 65786 535254
rect 66022 535018 66204 535254
rect 65604 534934 66204 535018
rect 65604 534698 65786 534934
rect 66022 534698 66204 534934
rect 65604 499254 66204 534698
rect 65604 499018 65786 499254
rect 66022 499018 66204 499254
rect 65604 498934 66204 499018
rect 65604 498698 65786 498934
rect 66022 498698 66204 498934
rect 65604 463254 66204 498698
rect 65604 463018 65786 463254
rect 66022 463018 66204 463254
rect 65604 462934 66204 463018
rect 65604 462698 65786 462934
rect 66022 462698 66204 462934
rect 65604 427254 66204 462698
rect 65604 427018 65786 427254
rect 66022 427018 66204 427254
rect 65604 426934 66204 427018
rect 65604 426698 65786 426934
rect 66022 426698 66204 426934
rect 65604 391254 66204 426698
rect 65604 391018 65786 391254
rect 66022 391018 66204 391254
rect 65604 390934 66204 391018
rect 65604 390698 65786 390934
rect 66022 390698 66204 390934
rect 65604 355254 66204 390698
rect 65604 355018 65786 355254
rect 66022 355018 66204 355254
rect 65604 354934 66204 355018
rect 65604 354698 65786 354934
rect 66022 354698 66204 354934
rect 65604 319254 66204 354698
rect 65604 319018 65786 319254
rect 66022 319018 66204 319254
rect 65604 318934 66204 319018
rect 65604 318698 65786 318934
rect 66022 318698 66204 318934
rect 65604 283254 66204 318698
rect 65604 283018 65786 283254
rect 66022 283018 66204 283254
rect 65604 282934 66204 283018
rect 65604 282698 65786 282934
rect 66022 282698 66204 282934
rect 65604 247254 66204 282698
rect 65604 247018 65786 247254
rect 66022 247018 66204 247254
rect 65604 246934 66204 247018
rect 65604 246698 65786 246934
rect 66022 246698 66204 246934
rect 65604 211254 66204 246698
rect 65604 211018 65786 211254
rect 66022 211018 66204 211254
rect 65604 210934 66204 211018
rect 65604 210698 65786 210934
rect 66022 210698 66204 210934
rect 65604 175254 66204 210698
rect 65604 175018 65786 175254
rect 66022 175018 66204 175254
rect 65604 174934 66204 175018
rect 65604 174698 65786 174934
rect 66022 174698 66204 174934
rect 65604 139254 66204 174698
rect 65604 139018 65786 139254
rect 66022 139018 66204 139254
rect 65604 138934 66204 139018
rect 65604 138698 65786 138934
rect 66022 138698 66204 138934
rect 65604 103254 66204 138698
rect 65604 103018 65786 103254
rect 66022 103018 66204 103254
rect 65604 102934 66204 103018
rect 65604 102698 65786 102934
rect 66022 102698 66204 102934
rect 65604 67254 66204 102698
rect 65604 67018 65786 67254
rect 66022 67018 66204 67254
rect 65604 66934 66204 67018
rect 65604 66698 65786 66934
rect 66022 66698 66204 66934
rect 65604 31254 66204 66698
rect 65604 31018 65786 31254
rect 66022 31018 66204 31254
rect 65604 30934 66204 31018
rect 65604 30698 65786 30934
rect 66022 30698 66204 30934
rect 47604 -6102 47786 -5866
rect 48022 -6102 48204 -5866
rect 47604 -6186 48204 -6102
rect 47604 -6422 47786 -6186
rect 48022 -6422 48204 -6186
rect 47604 -7364 48204 -6422
rect 65604 -6786 66204 30698
rect 72804 704838 73404 705780
rect 72804 704602 72986 704838
rect 73222 704602 73404 704838
rect 72804 704518 73404 704602
rect 72804 704282 72986 704518
rect 73222 704282 73404 704518
rect 72804 686454 73404 704282
rect 72804 686218 72986 686454
rect 73222 686218 73404 686454
rect 72804 686134 73404 686218
rect 72804 685898 72986 686134
rect 73222 685898 73404 686134
rect 72804 650454 73404 685898
rect 72804 650218 72986 650454
rect 73222 650218 73404 650454
rect 72804 650134 73404 650218
rect 72804 649898 72986 650134
rect 73222 649898 73404 650134
rect 72804 614454 73404 649898
rect 72804 614218 72986 614454
rect 73222 614218 73404 614454
rect 72804 614134 73404 614218
rect 72804 613898 72986 614134
rect 73222 613898 73404 614134
rect 72804 578454 73404 613898
rect 72804 578218 72986 578454
rect 73222 578218 73404 578454
rect 72804 578134 73404 578218
rect 72804 577898 72986 578134
rect 73222 577898 73404 578134
rect 72804 542454 73404 577898
rect 72804 542218 72986 542454
rect 73222 542218 73404 542454
rect 72804 542134 73404 542218
rect 72804 541898 72986 542134
rect 73222 541898 73404 542134
rect 72804 506454 73404 541898
rect 72804 506218 72986 506454
rect 73222 506218 73404 506454
rect 72804 506134 73404 506218
rect 72804 505898 72986 506134
rect 73222 505898 73404 506134
rect 72804 470454 73404 505898
rect 72804 470218 72986 470454
rect 73222 470218 73404 470454
rect 72804 470134 73404 470218
rect 72804 469898 72986 470134
rect 73222 469898 73404 470134
rect 72804 434454 73404 469898
rect 72804 434218 72986 434454
rect 73222 434218 73404 434454
rect 72804 434134 73404 434218
rect 72804 433898 72986 434134
rect 73222 433898 73404 434134
rect 72804 398454 73404 433898
rect 72804 398218 72986 398454
rect 73222 398218 73404 398454
rect 72804 398134 73404 398218
rect 72804 397898 72986 398134
rect 73222 397898 73404 398134
rect 72804 362454 73404 397898
rect 72804 362218 72986 362454
rect 73222 362218 73404 362454
rect 72804 362134 73404 362218
rect 72804 361898 72986 362134
rect 73222 361898 73404 362134
rect 72804 326454 73404 361898
rect 72804 326218 72986 326454
rect 73222 326218 73404 326454
rect 72804 326134 73404 326218
rect 72804 325898 72986 326134
rect 73222 325898 73404 326134
rect 72804 290454 73404 325898
rect 72804 290218 72986 290454
rect 73222 290218 73404 290454
rect 72804 290134 73404 290218
rect 72804 289898 72986 290134
rect 73222 289898 73404 290134
rect 72804 254454 73404 289898
rect 72804 254218 72986 254454
rect 73222 254218 73404 254454
rect 72804 254134 73404 254218
rect 72804 253898 72986 254134
rect 73222 253898 73404 254134
rect 72804 218454 73404 253898
rect 72804 218218 72986 218454
rect 73222 218218 73404 218454
rect 72804 218134 73404 218218
rect 72804 217898 72986 218134
rect 73222 217898 73404 218134
rect 72804 182454 73404 217898
rect 72804 182218 72986 182454
rect 73222 182218 73404 182454
rect 72804 182134 73404 182218
rect 72804 181898 72986 182134
rect 73222 181898 73404 182134
rect 72804 146454 73404 181898
rect 72804 146218 72986 146454
rect 73222 146218 73404 146454
rect 72804 146134 73404 146218
rect 72804 145898 72986 146134
rect 73222 145898 73404 146134
rect 72804 110454 73404 145898
rect 72804 110218 72986 110454
rect 73222 110218 73404 110454
rect 72804 110134 73404 110218
rect 72804 109898 72986 110134
rect 73222 109898 73404 110134
rect 72804 74454 73404 109898
rect 72804 74218 72986 74454
rect 73222 74218 73404 74454
rect 72804 74134 73404 74218
rect 72804 73898 72986 74134
rect 73222 73898 73404 74134
rect 72804 38454 73404 73898
rect 72804 38218 72986 38454
rect 73222 38218 73404 38454
rect 72804 38134 73404 38218
rect 72804 37898 72986 38134
rect 73222 37898 73404 38134
rect 72804 2454 73404 37898
rect 72804 2218 72986 2454
rect 73222 2218 73404 2454
rect 72804 2134 73404 2218
rect 72804 1898 72986 2134
rect 73222 1898 73404 2134
rect 72804 -346 73404 1898
rect 72804 -582 72986 -346
rect 73222 -582 73404 -346
rect 72804 -666 73404 -582
rect 72804 -902 72986 -666
rect 73222 -902 73404 -666
rect 72804 -1844 73404 -902
rect 76404 690054 77004 706122
rect 76404 689818 76586 690054
rect 76822 689818 77004 690054
rect 76404 689734 77004 689818
rect 76404 689498 76586 689734
rect 76822 689498 77004 689734
rect 76404 654054 77004 689498
rect 76404 653818 76586 654054
rect 76822 653818 77004 654054
rect 76404 653734 77004 653818
rect 76404 653498 76586 653734
rect 76822 653498 77004 653734
rect 76404 618054 77004 653498
rect 76404 617818 76586 618054
rect 76822 617818 77004 618054
rect 76404 617734 77004 617818
rect 76404 617498 76586 617734
rect 76822 617498 77004 617734
rect 76404 582054 77004 617498
rect 76404 581818 76586 582054
rect 76822 581818 77004 582054
rect 76404 581734 77004 581818
rect 76404 581498 76586 581734
rect 76822 581498 77004 581734
rect 76404 546054 77004 581498
rect 76404 545818 76586 546054
rect 76822 545818 77004 546054
rect 76404 545734 77004 545818
rect 76404 545498 76586 545734
rect 76822 545498 77004 545734
rect 76404 510054 77004 545498
rect 76404 509818 76586 510054
rect 76822 509818 77004 510054
rect 76404 509734 77004 509818
rect 76404 509498 76586 509734
rect 76822 509498 77004 509734
rect 76404 474054 77004 509498
rect 76404 473818 76586 474054
rect 76822 473818 77004 474054
rect 76404 473734 77004 473818
rect 76404 473498 76586 473734
rect 76822 473498 77004 473734
rect 76404 438054 77004 473498
rect 76404 437818 76586 438054
rect 76822 437818 77004 438054
rect 76404 437734 77004 437818
rect 76404 437498 76586 437734
rect 76822 437498 77004 437734
rect 76404 402054 77004 437498
rect 76404 401818 76586 402054
rect 76822 401818 77004 402054
rect 76404 401734 77004 401818
rect 76404 401498 76586 401734
rect 76822 401498 77004 401734
rect 76404 366054 77004 401498
rect 76404 365818 76586 366054
rect 76822 365818 77004 366054
rect 76404 365734 77004 365818
rect 76404 365498 76586 365734
rect 76822 365498 77004 365734
rect 76404 330054 77004 365498
rect 76404 329818 76586 330054
rect 76822 329818 77004 330054
rect 76404 329734 77004 329818
rect 76404 329498 76586 329734
rect 76822 329498 77004 329734
rect 76404 294054 77004 329498
rect 76404 293818 76586 294054
rect 76822 293818 77004 294054
rect 76404 293734 77004 293818
rect 76404 293498 76586 293734
rect 76822 293498 77004 293734
rect 76404 258054 77004 293498
rect 76404 257818 76586 258054
rect 76822 257818 77004 258054
rect 76404 257734 77004 257818
rect 76404 257498 76586 257734
rect 76822 257498 77004 257734
rect 76404 222054 77004 257498
rect 76404 221818 76586 222054
rect 76822 221818 77004 222054
rect 76404 221734 77004 221818
rect 76404 221498 76586 221734
rect 76822 221498 77004 221734
rect 76404 186054 77004 221498
rect 76404 185818 76586 186054
rect 76822 185818 77004 186054
rect 76404 185734 77004 185818
rect 76404 185498 76586 185734
rect 76822 185498 77004 185734
rect 76404 150054 77004 185498
rect 76404 149818 76586 150054
rect 76822 149818 77004 150054
rect 76404 149734 77004 149818
rect 76404 149498 76586 149734
rect 76822 149498 77004 149734
rect 76404 114054 77004 149498
rect 76404 113818 76586 114054
rect 76822 113818 77004 114054
rect 76404 113734 77004 113818
rect 76404 113498 76586 113734
rect 76822 113498 77004 113734
rect 76404 78054 77004 113498
rect 76404 77818 76586 78054
rect 76822 77818 77004 78054
rect 76404 77734 77004 77818
rect 76404 77498 76586 77734
rect 76822 77498 77004 77734
rect 76404 42054 77004 77498
rect 76404 41818 76586 42054
rect 76822 41818 77004 42054
rect 76404 41734 77004 41818
rect 76404 41498 76586 41734
rect 76822 41498 77004 41734
rect 76404 6054 77004 41498
rect 76404 5818 76586 6054
rect 76822 5818 77004 6054
rect 76404 5734 77004 5818
rect 76404 5498 76586 5734
rect 76822 5498 77004 5734
rect 76404 -2186 77004 5498
rect 76404 -2422 76586 -2186
rect 76822 -2422 77004 -2186
rect 76404 -2506 77004 -2422
rect 76404 -2742 76586 -2506
rect 76822 -2742 77004 -2506
rect 76404 -3684 77004 -2742
rect 80004 693654 80604 707962
rect 80004 693418 80186 693654
rect 80422 693418 80604 693654
rect 80004 693334 80604 693418
rect 80004 693098 80186 693334
rect 80422 693098 80604 693334
rect 80004 657654 80604 693098
rect 80004 657418 80186 657654
rect 80422 657418 80604 657654
rect 80004 657334 80604 657418
rect 80004 657098 80186 657334
rect 80422 657098 80604 657334
rect 80004 621654 80604 657098
rect 80004 621418 80186 621654
rect 80422 621418 80604 621654
rect 80004 621334 80604 621418
rect 80004 621098 80186 621334
rect 80422 621098 80604 621334
rect 80004 585654 80604 621098
rect 80004 585418 80186 585654
rect 80422 585418 80604 585654
rect 80004 585334 80604 585418
rect 80004 585098 80186 585334
rect 80422 585098 80604 585334
rect 80004 549654 80604 585098
rect 80004 549418 80186 549654
rect 80422 549418 80604 549654
rect 80004 549334 80604 549418
rect 80004 549098 80186 549334
rect 80422 549098 80604 549334
rect 80004 513654 80604 549098
rect 80004 513418 80186 513654
rect 80422 513418 80604 513654
rect 80004 513334 80604 513418
rect 80004 513098 80186 513334
rect 80422 513098 80604 513334
rect 80004 477654 80604 513098
rect 80004 477418 80186 477654
rect 80422 477418 80604 477654
rect 80004 477334 80604 477418
rect 80004 477098 80186 477334
rect 80422 477098 80604 477334
rect 80004 441654 80604 477098
rect 80004 441418 80186 441654
rect 80422 441418 80604 441654
rect 80004 441334 80604 441418
rect 80004 441098 80186 441334
rect 80422 441098 80604 441334
rect 80004 405654 80604 441098
rect 80004 405418 80186 405654
rect 80422 405418 80604 405654
rect 80004 405334 80604 405418
rect 80004 405098 80186 405334
rect 80422 405098 80604 405334
rect 80004 369654 80604 405098
rect 80004 369418 80186 369654
rect 80422 369418 80604 369654
rect 80004 369334 80604 369418
rect 80004 369098 80186 369334
rect 80422 369098 80604 369334
rect 80004 333654 80604 369098
rect 80004 333418 80186 333654
rect 80422 333418 80604 333654
rect 80004 333334 80604 333418
rect 80004 333098 80186 333334
rect 80422 333098 80604 333334
rect 80004 297654 80604 333098
rect 80004 297418 80186 297654
rect 80422 297418 80604 297654
rect 80004 297334 80604 297418
rect 80004 297098 80186 297334
rect 80422 297098 80604 297334
rect 80004 261654 80604 297098
rect 80004 261418 80186 261654
rect 80422 261418 80604 261654
rect 80004 261334 80604 261418
rect 80004 261098 80186 261334
rect 80422 261098 80604 261334
rect 80004 225654 80604 261098
rect 80004 225418 80186 225654
rect 80422 225418 80604 225654
rect 80004 225334 80604 225418
rect 80004 225098 80186 225334
rect 80422 225098 80604 225334
rect 80004 189654 80604 225098
rect 80004 189418 80186 189654
rect 80422 189418 80604 189654
rect 80004 189334 80604 189418
rect 80004 189098 80186 189334
rect 80422 189098 80604 189334
rect 80004 153654 80604 189098
rect 80004 153418 80186 153654
rect 80422 153418 80604 153654
rect 80004 153334 80604 153418
rect 80004 153098 80186 153334
rect 80422 153098 80604 153334
rect 80004 117654 80604 153098
rect 80004 117418 80186 117654
rect 80422 117418 80604 117654
rect 80004 117334 80604 117418
rect 80004 117098 80186 117334
rect 80422 117098 80604 117334
rect 80004 81654 80604 117098
rect 80004 81418 80186 81654
rect 80422 81418 80604 81654
rect 80004 81334 80604 81418
rect 80004 81098 80186 81334
rect 80422 81098 80604 81334
rect 80004 45654 80604 81098
rect 80004 45418 80186 45654
rect 80422 45418 80604 45654
rect 80004 45334 80604 45418
rect 80004 45098 80186 45334
rect 80422 45098 80604 45334
rect 80004 9654 80604 45098
rect 80004 9418 80186 9654
rect 80422 9418 80604 9654
rect 80004 9334 80604 9418
rect 80004 9098 80186 9334
rect 80422 9098 80604 9334
rect 80004 -4026 80604 9098
rect 80004 -4262 80186 -4026
rect 80422 -4262 80604 -4026
rect 80004 -4346 80604 -4262
rect 80004 -4582 80186 -4346
rect 80422 -4582 80604 -4346
rect 80004 -5524 80604 -4582
rect 83604 697254 84204 709802
rect 101604 711278 102204 711300
rect 101604 711042 101786 711278
rect 102022 711042 102204 711278
rect 101604 710958 102204 711042
rect 101604 710722 101786 710958
rect 102022 710722 102204 710958
rect 98004 709438 98604 709460
rect 98004 709202 98186 709438
rect 98422 709202 98604 709438
rect 98004 709118 98604 709202
rect 98004 708882 98186 709118
rect 98422 708882 98604 709118
rect 94404 707598 95004 707620
rect 94404 707362 94586 707598
rect 94822 707362 95004 707598
rect 94404 707278 95004 707362
rect 94404 707042 94586 707278
rect 94822 707042 95004 707278
rect 83604 697018 83786 697254
rect 84022 697018 84204 697254
rect 83604 696934 84204 697018
rect 83604 696698 83786 696934
rect 84022 696698 84204 696934
rect 83604 661254 84204 696698
rect 83604 661018 83786 661254
rect 84022 661018 84204 661254
rect 83604 660934 84204 661018
rect 83604 660698 83786 660934
rect 84022 660698 84204 660934
rect 83604 625254 84204 660698
rect 83604 625018 83786 625254
rect 84022 625018 84204 625254
rect 83604 624934 84204 625018
rect 83604 624698 83786 624934
rect 84022 624698 84204 624934
rect 83604 589254 84204 624698
rect 83604 589018 83786 589254
rect 84022 589018 84204 589254
rect 83604 588934 84204 589018
rect 83604 588698 83786 588934
rect 84022 588698 84204 588934
rect 83604 553254 84204 588698
rect 83604 553018 83786 553254
rect 84022 553018 84204 553254
rect 83604 552934 84204 553018
rect 83604 552698 83786 552934
rect 84022 552698 84204 552934
rect 83604 517254 84204 552698
rect 83604 517018 83786 517254
rect 84022 517018 84204 517254
rect 83604 516934 84204 517018
rect 83604 516698 83786 516934
rect 84022 516698 84204 516934
rect 83604 481254 84204 516698
rect 83604 481018 83786 481254
rect 84022 481018 84204 481254
rect 83604 480934 84204 481018
rect 83604 480698 83786 480934
rect 84022 480698 84204 480934
rect 83604 445254 84204 480698
rect 83604 445018 83786 445254
rect 84022 445018 84204 445254
rect 83604 444934 84204 445018
rect 83604 444698 83786 444934
rect 84022 444698 84204 444934
rect 83604 409254 84204 444698
rect 83604 409018 83786 409254
rect 84022 409018 84204 409254
rect 83604 408934 84204 409018
rect 83604 408698 83786 408934
rect 84022 408698 84204 408934
rect 83604 373254 84204 408698
rect 83604 373018 83786 373254
rect 84022 373018 84204 373254
rect 83604 372934 84204 373018
rect 83604 372698 83786 372934
rect 84022 372698 84204 372934
rect 83604 337254 84204 372698
rect 83604 337018 83786 337254
rect 84022 337018 84204 337254
rect 83604 336934 84204 337018
rect 83604 336698 83786 336934
rect 84022 336698 84204 336934
rect 83604 301254 84204 336698
rect 83604 301018 83786 301254
rect 84022 301018 84204 301254
rect 83604 300934 84204 301018
rect 83604 300698 83786 300934
rect 84022 300698 84204 300934
rect 83604 265254 84204 300698
rect 83604 265018 83786 265254
rect 84022 265018 84204 265254
rect 83604 264934 84204 265018
rect 83604 264698 83786 264934
rect 84022 264698 84204 264934
rect 83604 229254 84204 264698
rect 83604 229018 83786 229254
rect 84022 229018 84204 229254
rect 83604 228934 84204 229018
rect 83604 228698 83786 228934
rect 84022 228698 84204 228934
rect 83604 193254 84204 228698
rect 83604 193018 83786 193254
rect 84022 193018 84204 193254
rect 83604 192934 84204 193018
rect 83604 192698 83786 192934
rect 84022 192698 84204 192934
rect 83604 157254 84204 192698
rect 83604 157018 83786 157254
rect 84022 157018 84204 157254
rect 83604 156934 84204 157018
rect 83604 156698 83786 156934
rect 84022 156698 84204 156934
rect 83604 121254 84204 156698
rect 83604 121018 83786 121254
rect 84022 121018 84204 121254
rect 83604 120934 84204 121018
rect 83604 120698 83786 120934
rect 84022 120698 84204 120934
rect 83604 85254 84204 120698
rect 83604 85018 83786 85254
rect 84022 85018 84204 85254
rect 83604 84934 84204 85018
rect 83604 84698 83786 84934
rect 84022 84698 84204 84934
rect 83604 49254 84204 84698
rect 83604 49018 83786 49254
rect 84022 49018 84204 49254
rect 83604 48934 84204 49018
rect 83604 48698 83786 48934
rect 84022 48698 84204 48934
rect 83604 13254 84204 48698
rect 83604 13018 83786 13254
rect 84022 13018 84204 13254
rect 83604 12934 84204 13018
rect 83604 12698 83786 12934
rect 84022 12698 84204 12934
rect 65604 -7022 65786 -6786
rect 66022 -7022 66204 -6786
rect 65604 -7106 66204 -7022
rect 65604 -7342 65786 -7106
rect 66022 -7342 66204 -7106
rect 65604 -7364 66204 -7342
rect 83604 -5866 84204 12698
rect 90804 705758 91404 705780
rect 90804 705522 90986 705758
rect 91222 705522 91404 705758
rect 90804 705438 91404 705522
rect 90804 705202 90986 705438
rect 91222 705202 91404 705438
rect 90804 668454 91404 705202
rect 90804 668218 90986 668454
rect 91222 668218 91404 668454
rect 90804 668134 91404 668218
rect 90804 667898 90986 668134
rect 91222 667898 91404 668134
rect 90804 632454 91404 667898
rect 90804 632218 90986 632454
rect 91222 632218 91404 632454
rect 90804 632134 91404 632218
rect 90804 631898 90986 632134
rect 91222 631898 91404 632134
rect 90804 596454 91404 631898
rect 90804 596218 90986 596454
rect 91222 596218 91404 596454
rect 90804 596134 91404 596218
rect 90804 595898 90986 596134
rect 91222 595898 91404 596134
rect 90804 560454 91404 595898
rect 90804 560218 90986 560454
rect 91222 560218 91404 560454
rect 90804 560134 91404 560218
rect 90804 559898 90986 560134
rect 91222 559898 91404 560134
rect 90804 524454 91404 559898
rect 90804 524218 90986 524454
rect 91222 524218 91404 524454
rect 90804 524134 91404 524218
rect 90804 523898 90986 524134
rect 91222 523898 91404 524134
rect 90804 488454 91404 523898
rect 90804 488218 90986 488454
rect 91222 488218 91404 488454
rect 90804 488134 91404 488218
rect 90804 487898 90986 488134
rect 91222 487898 91404 488134
rect 90804 452454 91404 487898
rect 90804 452218 90986 452454
rect 91222 452218 91404 452454
rect 90804 452134 91404 452218
rect 90804 451898 90986 452134
rect 91222 451898 91404 452134
rect 90804 416454 91404 451898
rect 90804 416218 90986 416454
rect 91222 416218 91404 416454
rect 90804 416134 91404 416218
rect 90804 415898 90986 416134
rect 91222 415898 91404 416134
rect 90804 380454 91404 415898
rect 90804 380218 90986 380454
rect 91222 380218 91404 380454
rect 90804 380134 91404 380218
rect 90804 379898 90986 380134
rect 91222 379898 91404 380134
rect 90804 344454 91404 379898
rect 90804 344218 90986 344454
rect 91222 344218 91404 344454
rect 90804 344134 91404 344218
rect 90804 343898 90986 344134
rect 91222 343898 91404 344134
rect 90804 308454 91404 343898
rect 90804 308218 90986 308454
rect 91222 308218 91404 308454
rect 90804 308134 91404 308218
rect 90804 307898 90986 308134
rect 91222 307898 91404 308134
rect 90804 272454 91404 307898
rect 90804 272218 90986 272454
rect 91222 272218 91404 272454
rect 90804 272134 91404 272218
rect 90804 271898 90986 272134
rect 91222 271898 91404 272134
rect 90804 236454 91404 271898
rect 90804 236218 90986 236454
rect 91222 236218 91404 236454
rect 90804 236134 91404 236218
rect 90804 235898 90986 236134
rect 91222 235898 91404 236134
rect 90804 200454 91404 235898
rect 90804 200218 90986 200454
rect 91222 200218 91404 200454
rect 90804 200134 91404 200218
rect 90804 199898 90986 200134
rect 91222 199898 91404 200134
rect 90804 164454 91404 199898
rect 90804 164218 90986 164454
rect 91222 164218 91404 164454
rect 90804 164134 91404 164218
rect 90804 163898 90986 164134
rect 91222 163898 91404 164134
rect 90804 128454 91404 163898
rect 90804 128218 90986 128454
rect 91222 128218 91404 128454
rect 90804 128134 91404 128218
rect 90804 127898 90986 128134
rect 91222 127898 91404 128134
rect 90804 92454 91404 127898
rect 90804 92218 90986 92454
rect 91222 92218 91404 92454
rect 90804 92134 91404 92218
rect 90804 91898 90986 92134
rect 91222 91898 91404 92134
rect 90804 56454 91404 91898
rect 90804 56218 90986 56454
rect 91222 56218 91404 56454
rect 90804 56134 91404 56218
rect 90804 55898 90986 56134
rect 91222 55898 91404 56134
rect 90804 20454 91404 55898
rect 90804 20218 90986 20454
rect 91222 20218 91404 20454
rect 90804 20134 91404 20218
rect 90804 19898 90986 20134
rect 91222 19898 91404 20134
rect 90804 -1266 91404 19898
rect 90804 -1502 90986 -1266
rect 91222 -1502 91404 -1266
rect 90804 -1586 91404 -1502
rect 90804 -1822 90986 -1586
rect 91222 -1822 91404 -1586
rect 90804 -1844 91404 -1822
rect 94404 672054 95004 707042
rect 94404 671818 94586 672054
rect 94822 671818 95004 672054
rect 94404 671734 95004 671818
rect 94404 671498 94586 671734
rect 94822 671498 95004 671734
rect 94404 636054 95004 671498
rect 94404 635818 94586 636054
rect 94822 635818 95004 636054
rect 94404 635734 95004 635818
rect 94404 635498 94586 635734
rect 94822 635498 95004 635734
rect 94404 600054 95004 635498
rect 94404 599818 94586 600054
rect 94822 599818 95004 600054
rect 94404 599734 95004 599818
rect 94404 599498 94586 599734
rect 94822 599498 95004 599734
rect 94404 564054 95004 599498
rect 94404 563818 94586 564054
rect 94822 563818 95004 564054
rect 94404 563734 95004 563818
rect 94404 563498 94586 563734
rect 94822 563498 95004 563734
rect 94404 528054 95004 563498
rect 94404 527818 94586 528054
rect 94822 527818 95004 528054
rect 94404 527734 95004 527818
rect 94404 527498 94586 527734
rect 94822 527498 95004 527734
rect 94404 492054 95004 527498
rect 94404 491818 94586 492054
rect 94822 491818 95004 492054
rect 94404 491734 95004 491818
rect 94404 491498 94586 491734
rect 94822 491498 95004 491734
rect 94404 456054 95004 491498
rect 94404 455818 94586 456054
rect 94822 455818 95004 456054
rect 94404 455734 95004 455818
rect 94404 455498 94586 455734
rect 94822 455498 95004 455734
rect 94404 420054 95004 455498
rect 94404 419818 94586 420054
rect 94822 419818 95004 420054
rect 94404 419734 95004 419818
rect 94404 419498 94586 419734
rect 94822 419498 95004 419734
rect 94404 384054 95004 419498
rect 94404 383818 94586 384054
rect 94822 383818 95004 384054
rect 94404 383734 95004 383818
rect 94404 383498 94586 383734
rect 94822 383498 95004 383734
rect 94404 348054 95004 383498
rect 94404 347818 94586 348054
rect 94822 347818 95004 348054
rect 94404 347734 95004 347818
rect 94404 347498 94586 347734
rect 94822 347498 95004 347734
rect 94404 312054 95004 347498
rect 94404 311818 94586 312054
rect 94822 311818 95004 312054
rect 94404 311734 95004 311818
rect 94404 311498 94586 311734
rect 94822 311498 95004 311734
rect 94404 276054 95004 311498
rect 94404 275818 94586 276054
rect 94822 275818 95004 276054
rect 94404 275734 95004 275818
rect 94404 275498 94586 275734
rect 94822 275498 95004 275734
rect 94404 240054 95004 275498
rect 94404 239818 94586 240054
rect 94822 239818 95004 240054
rect 94404 239734 95004 239818
rect 94404 239498 94586 239734
rect 94822 239498 95004 239734
rect 94404 204054 95004 239498
rect 94404 203818 94586 204054
rect 94822 203818 95004 204054
rect 94404 203734 95004 203818
rect 94404 203498 94586 203734
rect 94822 203498 95004 203734
rect 94404 168054 95004 203498
rect 94404 167818 94586 168054
rect 94822 167818 95004 168054
rect 94404 167734 95004 167818
rect 94404 167498 94586 167734
rect 94822 167498 95004 167734
rect 94404 132054 95004 167498
rect 94404 131818 94586 132054
rect 94822 131818 95004 132054
rect 94404 131734 95004 131818
rect 94404 131498 94586 131734
rect 94822 131498 95004 131734
rect 94404 96054 95004 131498
rect 94404 95818 94586 96054
rect 94822 95818 95004 96054
rect 94404 95734 95004 95818
rect 94404 95498 94586 95734
rect 94822 95498 95004 95734
rect 94404 60054 95004 95498
rect 94404 59818 94586 60054
rect 94822 59818 95004 60054
rect 94404 59734 95004 59818
rect 94404 59498 94586 59734
rect 94822 59498 95004 59734
rect 94404 24054 95004 59498
rect 94404 23818 94586 24054
rect 94822 23818 95004 24054
rect 94404 23734 95004 23818
rect 94404 23498 94586 23734
rect 94822 23498 95004 23734
rect 94404 -3106 95004 23498
rect 94404 -3342 94586 -3106
rect 94822 -3342 95004 -3106
rect 94404 -3426 95004 -3342
rect 94404 -3662 94586 -3426
rect 94822 -3662 95004 -3426
rect 94404 -3684 95004 -3662
rect 98004 675654 98604 708882
rect 98004 675418 98186 675654
rect 98422 675418 98604 675654
rect 98004 675334 98604 675418
rect 98004 675098 98186 675334
rect 98422 675098 98604 675334
rect 98004 639654 98604 675098
rect 98004 639418 98186 639654
rect 98422 639418 98604 639654
rect 98004 639334 98604 639418
rect 98004 639098 98186 639334
rect 98422 639098 98604 639334
rect 98004 603654 98604 639098
rect 98004 603418 98186 603654
rect 98422 603418 98604 603654
rect 98004 603334 98604 603418
rect 98004 603098 98186 603334
rect 98422 603098 98604 603334
rect 98004 567654 98604 603098
rect 98004 567418 98186 567654
rect 98422 567418 98604 567654
rect 98004 567334 98604 567418
rect 98004 567098 98186 567334
rect 98422 567098 98604 567334
rect 98004 531654 98604 567098
rect 98004 531418 98186 531654
rect 98422 531418 98604 531654
rect 98004 531334 98604 531418
rect 98004 531098 98186 531334
rect 98422 531098 98604 531334
rect 98004 495654 98604 531098
rect 98004 495418 98186 495654
rect 98422 495418 98604 495654
rect 98004 495334 98604 495418
rect 98004 495098 98186 495334
rect 98422 495098 98604 495334
rect 98004 459654 98604 495098
rect 98004 459418 98186 459654
rect 98422 459418 98604 459654
rect 98004 459334 98604 459418
rect 98004 459098 98186 459334
rect 98422 459098 98604 459334
rect 98004 423654 98604 459098
rect 98004 423418 98186 423654
rect 98422 423418 98604 423654
rect 98004 423334 98604 423418
rect 98004 423098 98186 423334
rect 98422 423098 98604 423334
rect 98004 387654 98604 423098
rect 98004 387418 98186 387654
rect 98422 387418 98604 387654
rect 98004 387334 98604 387418
rect 98004 387098 98186 387334
rect 98422 387098 98604 387334
rect 98004 351654 98604 387098
rect 98004 351418 98186 351654
rect 98422 351418 98604 351654
rect 98004 351334 98604 351418
rect 98004 351098 98186 351334
rect 98422 351098 98604 351334
rect 98004 315654 98604 351098
rect 98004 315418 98186 315654
rect 98422 315418 98604 315654
rect 98004 315334 98604 315418
rect 98004 315098 98186 315334
rect 98422 315098 98604 315334
rect 98004 279654 98604 315098
rect 98004 279418 98186 279654
rect 98422 279418 98604 279654
rect 98004 279334 98604 279418
rect 98004 279098 98186 279334
rect 98422 279098 98604 279334
rect 98004 243654 98604 279098
rect 98004 243418 98186 243654
rect 98422 243418 98604 243654
rect 98004 243334 98604 243418
rect 98004 243098 98186 243334
rect 98422 243098 98604 243334
rect 98004 207654 98604 243098
rect 98004 207418 98186 207654
rect 98422 207418 98604 207654
rect 98004 207334 98604 207418
rect 98004 207098 98186 207334
rect 98422 207098 98604 207334
rect 98004 171654 98604 207098
rect 98004 171418 98186 171654
rect 98422 171418 98604 171654
rect 98004 171334 98604 171418
rect 98004 171098 98186 171334
rect 98422 171098 98604 171334
rect 98004 135654 98604 171098
rect 98004 135418 98186 135654
rect 98422 135418 98604 135654
rect 98004 135334 98604 135418
rect 98004 135098 98186 135334
rect 98422 135098 98604 135334
rect 98004 99654 98604 135098
rect 98004 99418 98186 99654
rect 98422 99418 98604 99654
rect 98004 99334 98604 99418
rect 98004 99098 98186 99334
rect 98422 99098 98604 99334
rect 98004 63654 98604 99098
rect 98004 63418 98186 63654
rect 98422 63418 98604 63654
rect 98004 63334 98604 63418
rect 98004 63098 98186 63334
rect 98422 63098 98604 63334
rect 98004 27654 98604 63098
rect 98004 27418 98186 27654
rect 98422 27418 98604 27654
rect 98004 27334 98604 27418
rect 98004 27098 98186 27334
rect 98422 27098 98604 27334
rect 98004 -4946 98604 27098
rect 98004 -5182 98186 -4946
rect 98422 -5182 98604 -4946
rect 98004 -5266 98604 -5182
rect 98004 -5502 98186 -5266
rect 98422 -5502 98604 -5266
rect 98004 -5524 98604 -5502
rect 101604 679254 102204 710722
rect 119604 710358 120204 711300
rect 119604 710122 119786 710358
rect 120022 710122 120204 710358
rect 119604 710038 120204 710122
rect 119604 709802 119786 710038
rect 120022 709802 120204 710038
rect 116004 708518 116604 709460
rect 116004 708282 116186 708518
rect 116422 708282 116604 708518
rect 116004 708198 116604 708282
rect 116004 707962 116186 708198
rect 116422 707962 116604 708198
rect 112404 706678 113004 707620
rect 112404 706442 112586 706678
rect 112822 706442 113004 706678
rect 112404 706358 113004 706442
rect 112404 706122 112586 706358
rect 112822 706122 113004 706358
rect 101604 679018 101786 679254
rect 102022 679018 102204 679254
rect 101604 678934 102204 679018
rect 101604 678698 101786 678934
rect 102022 678698 102204 678934
rect 101604 643254 102204 678698
rect 101604 643018 101786 643254
rect 102022 643018 102204 643254
rect 101604 642934 102204 643018
rect 101604 642698 101786 642934
rect 102022 642698 102204 642934
rect 101604 607254 102204 642698
rect 101604 607018 101786 607254
rect 102022 607018 102204 607254
rect 101604 606934 102204 607018
rect 101604 606698 101786 606934
rect 102022 606698 102204 606934
rect 101604 571254 102204 606698
rect 101604 571018 101786 571254
rect 102022 571018 102204 571254
rect 101604 570934 102204 571018
rect 101604 570698 101786 570934
rect 102022 570698 102204 570934
rect 101604 535254 102204 570698
rect 101604 535018 101786 535254
rect 102022 535018 102204 535254
rect 101604 534934 102204 535018
rect 101604 534698 101786 534934
rect 102022 534698 102204 534934
rect 101604 499254 102204 534698
rect 101604 499018 101786 499254
rect 102022 499018 102204 499254
rect 101604 498934 102204 499018
rect 101604 498698 101786 498934
rect 102022 498698 102204 498934
rect 101604 463254 102204 498698
rect 101604 463018 101786 463254
rect 102022 463018 102204 463254
rect 101604 462934 102204 463018
rect 101604 462698 101786 462934
rect 102022 462698 102204 462934
rect 101604 427254 102204 462698
rect 101604 427018 101786 427254
rect 102022 427018 102204 427254
rect 101604 426934 102204 427018
rect 101604 426698 101786 426934
rect 102022 426698 102204 426934
rect 101604 391254 102204 426698
rect 101604 391018 101786 391254
rect 102022 391018 102204 391254
rect 101604 390934 102204 391018
rect 101604 390698 101786 390934
rect 102022 390698 102204 390934
rect 101604 355254 102204 390698
rect 101604 355018 101786 355254
rect 102022 355018 102204 355254
rect 101604 354934 102204 355018
rect 101604 354698 101786 354934
rect 102022 354698 102204 354934
rect 101604 319254 102204 354698
rect 101604 319018 101786 319254
rect 102022 319018 102204 319254
rect 101604 318934 102204 319018
rect 101604 318698 101786 318934
rect 102022 318698 102204 318934
rect 101604 283254 102204 318698
rect 101604 283018 101786 283254
rect 102022 283018 102204 283254
rect 101604 282934 102204 283018
rect 101604 282698 101786 282934
rect 102022 282698 102204 282934
rect 101604 247254 102204 282698
rect 101604 247018 101786 247254
rect 102022 247018 102204 247254
rect 101604 246934 102204 247018
rect 101604 246698 101786 246934
rect 102022 246698 102204 246934
rect 101604 211254 102204 246698
rect 101604 211018 101786 211254
rect 102022 211018 102204 211254
rect 101604 210934 102204 211018
rect 101604 210698 101786 210934
rect 102022 210698 102204 210934
rect 101604 175254 102204 210698
rect 101604 175018 101786 175254
rect 102022 175018 102204 175254
rect 101604 174934 102204 175018
rect 101604 174698 101786 174934
rect 102022 174698 102204 174934
rect 101604 139254 102204 174698
rect 101604 139018 101786 139254
rect 102022 139018 102204 139254
rect 101604 138934 102204 139018
rect 101604 138698 101786 138934
rect 102022 138698 102204 138934
rect 101604 103254 102204 138698
rect 101604 103018 101786 103254
rect 102022 103018 102204 103254
rect 101604 102934 102204 103018
rect 101604 102698 101786 102934
rect 102022 102698 102204 102934
rect 101604 67254 102204 102698
rect 101604 67018 101786 67254
rect 102022 67018 102204 67254
rect 101604 66934 102204 67018
rect 101604 66698 101786 66934
rect 102022 66698 102204 66934
rect 101604 31254 102204 66698
rect 101604 31018 101786 31254
rect 102022 31018 102204 31254
rect 101604 30934 102204 31018
rect 101604 30698 101786 30934
rect 102022 30698 102204 30934
rect 83604 -6102 83786 -5866
rect 84022 -6102 84204 -5866
rect 83604 -6186 84204 -6102
rect 83604 -6422 83786 -6186
rect 84022 -6422 84204 -6186
rect 83604 -7364 84204 -6422
rect 101604 -6786 102204 30698
rect 108804 704838 109404 705780
rect 108804 704602 108986 704838
rect 109222 704602 109404 704838
rect 108804 704518 109404 704602
rect 108804 704282 108986 704518
rect 109222 704282 109404 704518
rect 108804 686454 109404 704282
rect 108804 686218 108986 686454
rect 109222 686218 109404 686454
rect 108804 686134 109404 686218
rect 108804 685898 108986 686134
rect 109222 685898 109404 686134
rect 108804 650454 109404 685898
rect 108804 650218 108986 650454
rect 109222 650218 109404 650454
rect 108804 650134 109404 650218
rect 108804 649898 108986 650134
rect 109222 649898 109404 650134
rect 108804 614454 109404 649898
rect 108804 614218 108986 614454
rect 109222 614218 109404 614454
rect 108804 614134 109404 614218
rect 108804 613898 108986 614134
rect 109222 613898 109404 614134
rect 108804 578454 109404 613898
rect 108804 578218 108986 578454
rect 109222 578218 109404 578454
rect 108804 578134 109404 578218
rect 108804 577898 108986 578134
rect 109222 577898 109404 578134
rect 108804 542454 109404 577898
rect 108804 542218 108986 542454
rect 109222 542218 109404 542454
rect 108804 542134 109404 542218
rect 108804 541898 108986 542134
rect 109222 541898 109404 542134
rect 108804 506454 109404 541898
rect 108804 506218 108986 506454
rect 109222 506218 109404 506454
rect 108804 506134 109404 506218
rect 108804 505898 108986 506134
rect 109222 505898 109404 506134
rect 108804 470454 109404 505898
rect 108804 470218 108986 470454
rect 109222 470218 109404 470454
rect 108804 470134 109404 470218
rect 108804 469898 108986 470134
rect 109222 469898 109404 470134
rect 108804 434454 109404 469898
rect 108804 434218 108986 434454
rect 109222 434218 109404 434454
rect 108804 434134 109404 434218
rect 108804 433898 108986 434134
rect 109222 433898 109404 434134
rect 108804 398454 109404 433898
rect 108804 398218 108986 398454
rect 109222 398218 109404 398454
rect 108804 398134 109404 398218
rect 108804 397898 108986 398134
rect 109222 397898 109404 398134
rect 108804 362454 109404 397898
rect 108804 362218 108986 362454
rect 109222 362218 109404 362454
rect 108804 362134 109404 362218
rect 108804 361898 108986 362134
rect 109222 361898 109404 362134
rect 108804 326454 109404 361898
rect 108804 326218 108986 326454
rect 109222 326218 109404 326454
rect 108804 326134 109404 326218
rect 108804 325898 108986 326134
rect 109222 325898 109404 326134
rect 108804 290454 109404 325898
rect 108804 290218 108986 290454
rect 109222 290218 109404 290454
rect 108804 290134 109404 290218
rect 108804 289898 108986 290134
rect 109222 289898 109404 290134
rect 108804 254454 109404 289898
rect 108804 254218 108986 254454
rect 109222 254218 109404 254454
rect 108804 254134 109404 254218
rect 108804 253898 108986 254134
rect 109222 253898 109404 254134
rect 108804 218454 109404 253898
rect 108804 218218 108986 218454
rect 109222 218218 109404 218454
rect 108804 218134 109404 218218
rect 108804 217898 108986 218134
rect 109222 217898 109404 218134
rect 108804 182454 109404 217898
rect 108804 182218 108986 182454
rect 109222 182218 109404 182454
rect 108804 182134 109404 182218
rect 108804 181898 108986 182134
rect 109222 181898 109404 182134
rect 108804 146454 109404 181898
rect 108804 146218 108986 146454
rect 109222 146218 109404 146454
rect 108804 146134 109404 146218
rect 108804 145898 108986 146134
rect 109222 145898 109404 146134
rect 108804 110454 109404 145898
rect 108804 110218 108986 110454
rect 109222 110218 109404 110454
rect 108804 110134 109404 110218
rect 108804 109898 108986 110134
rect 109222 109898 109404 110134
rect 108804 74454 109404 109898
rect 108804 74218 108986 74454
rect 109222 74218 109404 74454
rect 108804 74134 109404 74218
rect 108804 73898 108986 74134
rect 109222 73898 109404 74134
rect 108804 38454 109404 73898
rect 108804 38218 108986 38454
rect 109222 38218 109404 38454
rect 108804 38134 109404 38218
rect 108804 37898 108986 38134
rect 109222 37898 109404 38134
rect 108804 2454 109404 37898
rect 108804 2218 108986 2454
rect 109222 2218 109404 2454
rect 108804 2134 109404 2218
rect 108804 1898 108986 2134
rect 109222 1898 109404 2134
rect 108804 -346 109404 1898
rect 108804 -582 108986 -346
rect 109222 -582 109404 -346
rect 108804 -666 109404 -582
rect 108804 -902 108986 -666
rect 109222 -902 109404 -666
rect 108804 -1844 109404 -902
rect 112404 690054 113004 706122
rect 112404 689818 112586 690054
rect 112822 689818 113004 690054
rect 112404 689734 113004 689818
rect 112404 689498 112586 689734
rect 112822 689498 113004 689734
rect 112404 654054 113004 689498
rect 112404 653818 112586 654054
rect 112822 653818 113004 654054
rect 112404 653734 113004 653818
rect 112404 653498 112586 653734
rect 112822 653498 113004 653734
rect 112404 618054 113004 653498
rect 112404 617818 112586 618054
rect 112822 617818 113004 618054
rect 112404 617734 113004 617818
rect 112404 617498 112586 617734
rect 112822 617498 113004 617734
rect 112404 582054 113004 617498
rect 112404 581818 112586 582054
rect 112822 581818 113004 582054
rect 112404 581734 113004 581818
rect 112404 581498 112586 581734
rect 112822 581498 113004 581734
rect 112404 546054 113004 581498
rect 112404 545818 112586 546054
rect 112822 545818 113004 546054
rect 112404 545734 113004 545818
rect 112404 545498 112586 545734
rect 112822 545498 113004 545734
rect 112404 510054 113004 545498
rect 112404 509818 112586 510054
rect 112822 509818 113004 510054
rect 112404 509734 113004 509818
rect 112404 509498 112586 509734
rect 112822 509498 113004 509734
rect 112404 474054 113004 509498
rect 112404 473818 112586 474054
rect 112822 473818 113004 474054
rect 112404 473734 113004 473818
rect 112404 473498 112586 473734
rect 112822 473498 113004 473734
rect 112404 438054 113004 473498
rect 112404 437818 112586 438054
rect 112822 437818 113004 438054
rect 112404 437734 113004 437818
rect 112404 437498 112586 437734
rect 112822 437498 113004 437734
rect 112404 402054 113004 437498
rect 112404 401818 112586 402054
rect 112822 401818 113004 402054
rect 112404 401734 113004 401818
rect 112404 401498 112586 401734
rect 112822 401498 113004 401734
rect 112404 366054 113004 401498
rect 112404 365818 112586 366054
rect 112822 365818 113004 366054
rect 112404 365734 113004 365818
rect 112404 365498 112586 365734
rect 112822 365498 113004 365734
rect 112404 330054 113004 365498
rect 112404 329818 112586 330054
rect 112822 329818 113004 330054
rect 112404 329734 113004 329818
rect 112404 329498 112586 329734
rect 112822 329498 113004 329734
rect 112404 294054 113004 329498
rect 112404 293818 112586 294054
rect 112822 293818 113004 294054
rect 112404 293734 113004 293818
rect 112404 293498 112586 293734
rect 112822 293498 113004 293734
rect 112404 258054 113004 293498
rect 112404 257818 112586 258054
rect 112822 257818 113004 258054
rect 112404 257734 113004 257818
rect 112404 257498 112586 257734
rect 112822 257498 113004 257734
rect 112404 222054 113004 257498
rect 112404 221818 112586 222054
rect 112822 221818 113004 222054
rect 112404 221734 113004 221818
rect 112404 221498 112586 221734
rect 112822 221498 113004 221734
rect 112404 186054 113004 221498
rect 112404 185818 112586 186054
rect 112822 185818 113004 186054
rect 112404 185734 113004 185818
rect 112404 185498 112586 185734
rect 112822 185498 113004 185734
rect 112404 150054 113004 185498
rect 112404 149818 112586 150054
rect 112822 149818 113004 150054
rect 112404 149734 113004 149818
rect 112404 149498 112586 149734
rect 112822 149498 113004 149734
rect 112404 114054 113004 149498
rect 112404 113818 112586 114054
rect 112822 113818 113004 114054
rect 112404 113734 113004 113818
rect 112404 113498 112586 113734
rect 112822 113498 113004 113734
rect 112404 78054 113004 113498
rect 112404 77818 112586 78054
rect 112822 77818 113004 78054
rect 112404 77734 113004 77818
rect 112404 77498 112586 77734
rect 112822 77498 113004 77734
rect 112404 42054 113004 77498
rect 112404 41818 112586 42054
rect 112822 41818 113004 42054
rect 112404 41734 113004 41818
rect 112404 41498 112586 41734
rect 112822 41498 113004 41734
rect 112404 6054 113004 41498
rect 112404 5818 112586 6054
rect 112822 5818 113004 6054
rect 112404 5734 113004 5818
rect 112404 5498 112586 5734
rect 112822 5498 113004 5734
rect 112404 -2186 113004 5498
rect 112404 -2422 112586 -2186
rect 112822 -2422 113004 -2186
rect 112404 -2506 113004 -2422
rect 112404 -2742 112586 -2506
rect 112822 -2742 113004 -2506
rect 112404 -3684 113004 -2742
rect 116004 693654 116604 707962
rect 116004 693418 116186 693654
rect 116422 693418 116604 693654
rect 116004 693334 116604 693418
rect 116004 693098 116186 693334
rect 116422 693098 116604 693334
rect 116004 657654 116604 693098
rect 116004 657418 116186 657654
rect 116422 657418 116604 657654
rect 116004 657334 116604 657418
rect 116004 657098 116186 657334
rect 116422 657098 116604 657334
rect 116004 621654 116604 657098
rect 116004 621418 116186 621654
rect 116422 621418 116604 621654
rect 116004 621334 116604 621418
rect 116004 621098 116186 621334
rect 116422 621098 116604 621334
rect 116004 585654 116604 621098
rect 116004 585418 116186 585654
rect 116422 585418 116604 585654
rect 116004 585334 116604 585418
rect 116004 585098 116186 585334
rect 116422 585098 116604 585334
rect 116004 549654 116604 585098
rect 116004 549418 116186 549654
rect 116422 549418 116604 549654
rect 116004 549334 116604 549418
rect 116004 549098 116186 549334
rect 116422 549098 116604 549334
rect 116004 513654 116604 549098
rect 116004 513418 116186 513654
rect 116422 513418 116604 513654
rect 116004 513334 116604 513418
rect 116004 513098 116186 513334
rect 116422 513098 116604 513334
rect 116004 477654 116604 513098
rect 116004 477418 116186 477654
rect 116422 477418 116604 477654
rect 116004 477334 116604 477418
rect 116004 477098 116186 477334
rect 116422 477098 116604 477334
rect 116004 441654 116604 477098
rect 116004 441418 116186 441654
rect 116422 441418 116604 441654
rect 116004 441334 116604 441418
rect 116004 441098 116186 441334
rect 116422 441098 116604 441334
rect 116004 405654 116604 441098
rect 116004 405418 116186 405654
rect 116422 405418 116604 405654
rect 116004 405334 116604 405418
rect 116004 405098 116186 405334
rect 116422 405098 116604 405334
rect 116004 369654 116604 405098
rect 116004 369418 116186 369654
rect 116422 369418 116604 369654
rect 116004 369334 116604 369418
rect 116004 369098 116186 369334
rect 116422 369098 116604 369334
rect 116004 333654 116604 369098
rect 116004 333418 116186 333654
rect 116422 333418 116604 333654
rect 116004 333334 116604 333418
rect 116004 333098 116186 333334
rect 116422 333098 116604 333334
rect 116004 297654 116604 333098
rect 116004 297418 116186 297654
rect 116422 297418 116604 297654
rect 116004 297334 116604 297418
rect 116004 297098 116186 297334
rect 116422 297098 116604 297334
rect 116004 261654 116604 297098
rect 116004 261418 116186 261654
rect 116422 261418 116604 261654
rect 116004 261334 116604 261418
rect 116004 261098 116186 261334
rect 116422 261098 116604 261334
rect 116004 225654 116604 261098
rect 116004 225418 116186 225654
rect 116422 225418 116604 225654
rect 116004 225334 116604 225418
rect 116004 225098 116186 225334
rect 116422 225098 116604 225334
rect 116004 189654 116604 225098
rect 116004 189418 116186 189654
rect 116422 189418 116604 189654
rect 116004 189334 116604 189418
rect 116004 189098 116186 189334
rect 116422 189098 116604 189334
rect 116004 153654 116604 189098
rect 116004 153418 116186 153654
rect 116422 153418 116604 153654
rect 116004 153334 116604 153418
rect 116004 153098 116186 153334
rect 116422 153098 116604 153334
rect 116004 117654 116604 153098
rect 116004 117418 116186 117654
rect 116422 117418 116604 117654
rect 116004 117334 116604 117418
rect 116004 117098 116186 117334
rect 116422 117098 116604 117334
rect 116004 81654 116604 117098
rect 116004 81418 116186 81654
rect 116422 81418 116604 81654
rect 116004 81334 116604 81418
rect 116004 81098 116186 81334
rect 116422 81098 116604 81334
rect 116004 45654 116604 81098
rect 116004 45418 116186 45654
rect 116422 45418 116604 45654
rect 116004 45334 116604 45418
rect 116004 45098 116186 45334
rect 116422 45098 116604 45334
rect 116004 9654 116604 45098
rect 116004 9418 116186 9654
rect 116422 9418 116604 9654
rect 116004 9334 116604 9418
rect 116004 9098 116186 9334
rect 116422 9098 116604 9334
rect 116004 -4026 116604 9098
rect 116004 -4262 116186 -4026
rect 116422 -4262 116604 -4026
rect 116004 -4346 116604 -4262
rect 116004 -4582 116186 -4346
rect 116422 -4582 116604 -4346
rect 116004 -5524 116604 -4582
rect 119604 697254 120204 709802
rect 137604 711278 138204 711300
rect 137604 711042 137786 711278
rect 138022 711042 138204 711278
rect 137604 710958 138204 711042
rect 137604 710722 137786 710958
rect 138022 710722 138204 710958
rect 134004 709438 134604 709460
rect 134004 709202 134186 709438
rect 134422 709202 134604 709438
rect 134004 709118 134604 709202
rect 134004 708882 134186 709118
rect 134422 708882 134604 709118
rect 130404 707598 131004 707620
rect 130404 707362 130586 707598
rect 130822 707362 131004 707598
rect 130404 707278 131004 707362
rect 130404 707042 130586 707278
rect 130822 707042 131004 707278
rect 119604 697018 119786 697254
rect 120022 697018 120204 697254
rect 119604 696934 120204 697018
rect 119604 696698 119786 696934
rect 120022 696698 120204 696934
rect 119604 661254 120204 696698
rect 119604 661018 119786 661254
rect 120022 661018 120204 661254
rect 119604 660934 120204 661018
rect 119604 660698 119786 660934
rect 120022 660698 120204 660934
rect 119604 625254 120204 660698
rect 119604 625018 119786 625254
rect 120022 625018 120204 625254
rect 119604 624934 120204 625018
rect 119604 624698 119786 624934
rect 120022 624698 120204 624934
rect 119604 589254 120204 624698
rect 119604 589018 119786 589254
rect 120022 589018 120204 589254
rect 119604 588934 120204 589018
rect 119604 588698 119786 588934
rect 120022 588698 120204 588934
rect 119604 553254 120204 588698
rect 119604 553018 119786 553254
rect 120022 553018 120204 553254
rect 119604 552934 120204 553018
rect 119604 552698 119786 552934
rect 120022 552698 120204 552934
rect 119604 517254 120204 552698
rect 119604 517018 119786 517254
rect 120022 517018 120204 517254
rect 119604 516934 120204 517018
rect 119604 516698 119786 516934
rect 120022 516698 120204 516934
rect 119604 481254 120204 516698
rect 119604 481018 119786 481254
rect 120022 481018 120204 481254
rect 119604 480934 120204 481018
rect 119604 480698 119786 480934
rect 120022 480698 120204 480934
rect 119604 445254 120204 480698
rect 119604 445018 119786 445254
rect 120022 445018 120204 445254
rect 119604 444934 120204 445018
rect 119604 444698 119786 444934
rect 120022 444698 120204 444934
rect 119604 409254 120204 444698
rect 119604 409018 119786 409254
rect 120022 409018 120204 409254
rect 119604 408934 120204 409018
rect 119604 408698 119786 408934
rect 120022 408698 120204 408934
rect 119604 373254 120204 408698
rect 119604 373018 119786 373254
rect 120022 373018 120204 373254
rect 119604 372934 120204 373018
rect 119604 372698 119786 372934
rect 120022 372698 120204 372934
rect 119604 337254 120204 372698
rect 119604 337018 119786 337254
rect 120022 337018 120204 337254
rect 119604 336934 120204 337018
rect 119604 336698 119786 336934
rect 120022 336698 120204 336934
rect 119604 301254 120204 336698
rect 119604 301018 119786 301254
rect 120022 301018 120204 301254
rect 119604 300934 120204 301018
rect 119604 300698 119786 300934
rect 120022 300698 120204 300934
rect 119604 265254 120204 300698
rect 119604 265018 119786 265254
rect 120022 265018 120204 265254
rect 119604 264934 120204 265018
rect 119604 264698 119786 264934
rect 120022 264698 120204 264934
rect 119604 229254 120204 264698
rect 119604 229018 119786 229254
rect 120022 229018 120204 229254
rect 119604 228934 120204 229018
rect 119604 228698 119786 228934
rect 120022 228698 120204 228934
rect 119604 193254 120204 228698
rect 119604 193018 119786 193254
rect 120022 193018 120204 193254
rect 119604 192934 120204 193018
rect 119604 192698 119786 192934
rect 120022 192698 120204 192934
rect 119604 157254 120204 192698
rect 119604 157018 119786 157254
rect 120022 157018 120204 157254
rect 119604 156934 120204 157018
rect 119604 156698 119786 156934
rect 120022 156698 120204 156934
rect 119604 121254 120204 156698
rect 119604 121018 119786 121254
rect 120022 121018 120204 121254
rect 119604 120934 120204 121018
rect 119604 120698 119786 120934
rect 120022 120698 120204 120934
rect 119604 85254 120204 120698
rect 119604 85018 119786 85254
rect 120022 85018 120204 85254
rect 119604 84934 120204 85018
rect 119604 84698 119786 84934
rect 120022 84698 120204 84934
rect 119604 49254 120204 84698
rect 119604 49018 119786 49254
rect 120022 49018 120204 49254
rect 119604 48934 120204 49018
rect 119604 48698 119786 48934
rect 120022 48698 120204 48934
rect 119604 13254 120204 48698
rect 119604 13018 119786 13254
rect 120022 13018 120204 13254
rect 119604 12934 120204 13018
rect 119604 12698 119786 12934
rect 120022 12698 120204 12934
rect 101604 -7022 101786 -6786
rect 102022 -7022 102204 -6786
rect 101604 -7106 102204 -7022
rect 101604 -7342 101786 -7106
rect 102022 -7342 102204 -7106
rect 101604 -7364 102204 -7342
rect 119604 -5866 120204 12698
rect 126804 705758 127404 705780
rect 126804 705522 126986 705758
rect 127222 705522 127404 705758
rect 126804 705438 127404 705522
rect 126804 705202 126986 705438
rect 127222 705202 127404 705438
rect 126804 668454 127404 705202
rect 126804 668218 126986 668454
rect 127222 668218 127404 668454
rect 126804 668134 127404 668218
rect 126804 667898 126986 668134
rect 127222 667898 127404 668134
rect 126804 632454 127404 667898
rect 126804 632218 126986 632454
rect 127222 632218 127404 632454
rect 126804 632134 127404 632218
rect 126804 631898 126986 632134
rect 127222 631898 127404 632134
rect 126804 596454 127404 631898
rect 126804 596218 126986 596454
rect 127222 596218 127404 596454
rect 126804 596134 127404 596218
rect 126804 595898 126986 596134
rect 127222 595898 127404 596134
rect 126804 560454 127404 595898
rect 126804 560218 126986 560454
rect 127222 560218 127404 560454
rect 126804 560134 127404 560218
rect 126804 559898 126986 560134
rect 127222 559898 127404 560134
rect 126804 524454 127404 559898
rect 126804 524218 126986 524454
rect 127222 524218 127404 524454
rect 126804 524134 127404 524218
rect 126804 523898 126986 524134
rect 127222 523898 127404 524134
rect 126804 488454 127404 523898
rect 126804 488218 126986 488454
rect 127222 488218 127404 488454
rect 126804 488134 127404 488218
rect 126804 487898 126986 488134
rect 127222 487898 127404 488134
rect 126804 452454 127404 487898
rect 126804 452218 126986 452454
rect 127222 452218 127404 452454
rect 126804 452134 127404 452218
rect 126804 451898 126986 452134
rect 127222 451898 127404 452134
rect 126804 416454 127404 451898
rect 126804 416218 126986 416454
rect 127222 416218 127404 416454
rect 126804 416134 127404 416218
rect 126804 415898 126986 416134
rect 127222 415898 127404 416134
rect 126804 380454 127404 415898
rect 126804 380218 126986 380454
rect 127222 380218 127404 380454
rect 126804 380134 127404 380218
rect 126804 379898 126986 380134
rect 127222 379898 127404 380134
rect 126804 344454 127404 379898
rect 126804 344218 126986 344454
rect 127222 344218 127404 344454
rect 126804 344134 127404 344218
rect 126804 343898 126986 344134
rect 127222 343898 127404 344134
rect 126804 308454 127404 343898
rect 126804 308218 126986 308454
rect 127222 308218 127404 308454
rect 126804 308134 127404 308218
rect 126804 307898 126986 308134
rect 127222 307898 127404 308134
rect 126804 272454 127404 307898
rect 126804 272218 126986 272454
rect 127222 272218 127404 272454
rect 126804 272134 127404 272218
rect 126804 271898 126986 272134
rect 127222 271898 127404 272134
rect 126804 236454 127404 271898
rect 126804 236218 126986 236454
rect 127222 236218 127404 236454
rect 126804 236134 127404 236218
rect 126804 235898 126986 236134
rect 127222 235898 127404 236134
rect 126804 200454 127404 235898
rect 126804 200218 126986 200454
rect 127222 200218 127404 200454
rect 126804 200134 127404 200218
rect 126804 199898 126986 200134
rect 127222 199898 127404 200134
rect 126804 164454 127404 199898
rect 126804 164218 126986 164454
rect 127222 164218 127404 164454
rect 126804 164134 127404 164218
rect 126804 163898 126986 164134
rect 127222 163898 127404 164134
rect 126804 128454 127404 163898
rect 126804 128218 126986 128454
rect 127222 128218 127404 128454
rect 126804 128134 127404 128218
rect 126804 127898 126986 128134
rect 127222 127898 127404 128134
rect 126804 92454 127404 127898
rect 126804 92218 126986 92454
rect 127222 92218 127404 92454
rect 126804 92134 127404 92218
rect 126804 91898 126986 92134
rect 127222 91898 127404 92134
rect 126804 56454 127404 91898
rect 126804 56218 126986 56454
rect 127222 56218 127404 56454
rect 126804 56134 127404 56218
rect 126804 55898 126986 56134
rect 127222 55898 127404 56134
rect 126804 20454 127404 55898
rect 126804 20218 126986 20454
rect 127222 20218 127404 20454
rect 126804 20134 127404 20218
rect 126804 19898 126986 20134
rect 127222 19898 127404 20134
rect 126804 -1266 127404 19898
rect 126804 -1502 126986 -1266
rect 127222 -1502 127404 -1266
rect 126804 -1586 127404 -1502
rect 126804 -1822 126986 -1586
rect 127222 -1822 127404 -1586
rect 126804 -1844 127404 -1822
rect 130404 672054 131004 707042
rect 130404 671818 130586 672054
rect 130822 671818 131004 672054
rect 130404 671734 131004 671818
rect 130404 671498 130586 671734
rect 130822 671498 131004 671734
rect 130404 636054 131004 671498
rect 130404 635818 130586 636054
rect 130822 635818 131004 636054
rect 130404 635734 131004 635818
rect 130404 635498 130586 635734
rect 130822 635498 131004 635734
rect 130404 600054 131004 635498
rect 130404 599818 130586 600054
rect 130822 599818 131004 600054
rect 130404 599734 131004 599818
rect 130404 599498 130586 599734
rect 130822 599498 131004 599734
rect 130404 564054 131004 599498
rect 130404 563818 130586 564054
rect 130822 563818 131004 564054
rect 130404 563734 131004 563818
rect 130404 563498 130586 563734
rect 130822 563498 131004 563734
rect 130404 528054 131004 563498
rect 130404 527818 130586 528054
rect 130822 527818 131004 528054
rect 130404 527734 131004 527818
rect 130404 527498 130586 527734
rect 130822 527498 131004 527734
rect 130404 492054 131004 527498
rect 130404 491818 130586 492054
rect 130822 491818 131004 492054
rect 130404 491734 131004 491818
rect 130404 491498 130586 491734
rect 130822 491498 131004 491734
rect 130404 456054 131004 491498
rect 130404 455818 130586 456054
rect 130822 455818 131004 456054
rect 130404 455734 131004 455818
rect 130404 455498 130586 455734
rect 130822 455498 131004 455734
rect 130404 420054 131004 455498
rect 130404 419818 130586 420054
rect 130822 419818 131004 420054
rect 130404 419734 131004 419818
rect 130404 419498 130586 419734
rect 130822 419498 131004 419734
rect 130404 384054 131004 419498
rect 130404 383818 130586 384054
rect 130822 383818 131004 384054
rect 130404 383734 131004 383818
rect 130404 383498 130586 383734
rect 130822 383498 131004 383734
rect 130404 348054 131004 383498
rect 130404 347818 130586 348054
rect 130822 347818 131004 348054
rect 130404 347734 131004 347818
rect 130404 347498 130586 347734
rect 130822 347498 131004 347734
rect 130404 312054 131004 347498
rect 130404 311818 130586 312054
rect 130822 311818 131004 312054
rect 130404 311734 131004 311818
rect 130404 311498 130586 311734
rect 130822 311498 131004 311734
rect 130404 276054 131004 311498
rect 130404 275818 130586 276054
rect 130822 275818 131004 276054
rect 130404 275734 131004 275818
rect 130404 275498 130586 275734
rect 130822 275498 131004 275734
rect 130404 240054 131004 275498
rect 130404 239818 130586 240054
rect 130822 239818 131004 240054
rect 130404 239734 131004 239818
rect 130404 239498 130586 239734
rect 130822 239498 131004 239734
rect 130404 204054 131004 239498
rect 130404 203818 130586 204054
rect 130822 203818 131004 204054
rect 130404 203734 131004 203818
rect 130404 203498 130586 203734
rect 130822 203498 131004 203734
rect 130404 168054 131004 203498
rect 130404 167818 130586 168054
rect 130822 167818 131004 168054
rect 130404 167734 131004 167818
rect 130404 167498 130586 167734
rect 130822 167498 131004 167734
rect 130404 132054 131004 167498
rect 130404 131818 130586 132054
rect 130822 131818 131004 132054
rect 130404 131734 131004 131818
rect 130404 131498 130586 131734
rect 130822 131498 131004 131734
rect 130404 96054 131004 131498
rect 130404 95818 130586 96054
rect 130822 95818 131004 96054
rect 130404 95734 131004 95818
rect 130404 95498 130586 95734
rect 130822 95498 131004 95734
rect 130404 60054 131004 95498
rect 130404 59818 130586 60054
rect 130822 59818 131004 60054
rect 130404 59734 131004 59818
rect 130404 59498 130586 59734
rect 130822 59498 131004 59734
rect 130404 24054 131004 59498
rect 130404 23818 130586 24054
rect 130822 23818 131004 24054
rect 130404 23734 131004 23818
rect 130404 23498 130586 23734
rect 130822 23498 131004 23734
rect 130404 -3106 131004 23498
rect 130404 -3342 130586 -3106
rect 130822 -3342 131004 -3106
rect 130404 -3426 131004 -3342
rect 130404 -3662 130586 -3426
rect 130822 -3662 131004 -3426
rect 130404 -3684 131004 -3662
rect 134004 675654 134604 708882
rect 134004 675418 134186 675654
rect 134422 675418 134604 675654
rect 134004 675334 134604 675418
rect 134004 675098 134186 675334
rect 134422 675098 134604 675334
rect 134004 639654 134604 675098
rect 134004 639418 134186 639654
rect 134422 639418 134604 639654
rect 134004 639334 134604 639418
rect 134004 639098 134186 639334
rect 134422 639098 134604 639334
rect 134004 603654 134604 639098
rect 134004 603418 134186 603654
rect 134422 603418 134604 603654
rect 134004 603334 134604 603418
rect 134004 603098 134186 603334
rect 134422 603098 134604 603334
rect 134004 567654 134604 603098
rect 134004 567418 134186 567654
rect 134422 567418 134604 567654
rect 134004 567334 134604 567418
rect 134004 567098 134186 567334
rect 134422 567098 134604 567334
rect 134004 531654 134604 567098
rect 134004 531418 134186 531654
rect 134422 531418 134604 531654
rect 134004 531334 134604 531418
rect 134004 531098 134186 531334
rect 134422 531098 134604 531334
rect 134004 495654 134604 531098
rect 134004 495418 134186 495654
rect 134422 495418 134604 495654
rect 134004 495334 134604 495418
rect 134004 495098 134186 495334
rect 134422 495098 134604 495334
rect 134004 459654 134604 495098
rect 134004 459418 134186 459654
rect 134422 459418 134604 459654
rect 134004 459334 134604 459418
rect 134004 459098 134186 459334
rect 134422 459098 134604 459334
rect 134004 423654 134604 459098
rect 134004 423418 134186 423654
rect 134422 423418 134604 423654
rect 134004 423334 134604 423418
rect 134004 423098 134186 423334
rect 134422 423098 134604 423334
rect 134004 387654 134604 423098
rect 134004 387418 134186 387654
rect 134422 387418 134604 387654
rect 134004 387334 134604 387418
rect 134004 387098 134186 387334
rect 134422 387098 134604 387334
rect 134004 351654 134604 387098
rect 134004 351418 134186 351654
rect 134422 351418 134604 351654
rect 134004 351334 134604 351418
rect 134004 351098 134186 351334
rect 134422 351098 134604 351334
rect 134004 315654 134604 351098
rect 134004 315418 134186 315654
rect 134422 315418 134604 315654
rect 134004 315334 134604 315418
rect 134004 315098 134186 315334
rect 134422 315098 134604 315334
rect 134004 279654 134604 315098
rect 134004 279418 134186 279654
rect 134422 279418 134604 279654
rect 134004 279334 134604 279418
rect 134004 279098 134186 279334
rect 134422 279098 134604 279334
rect 134004 243654 134604 279098
rect 134004 243418 134186 243654
rect 134422 243418 134604 243654
rect 134004 243334 134604 243418
rect 134004 243098 134186 243334
rect 134422 243098 134604 243334
rect 134004 207654 134604 243098
rect 134004 207418 134186 207654
rect 134422 207418 134604 207654
rect 134004 207334 134604 207418
rect 134004 207098 134186 207334
rect 134422 207098 134604 207334
rect 134004 171654 134604 207098
rect 134004 171418 134186 171654
rect 134422 171418 134604 171654
rect 134004 171334 134604 171418
rect 134004 171098 134186 171334
rect 134422 171098 134604 171334
rect 134004 135654 134604 171098
rect 134004 135418 134186 135654
rect 134422 135418 134604 135654
rect 134004 135334 134604 135418
rect 134004 135098 134186 135334
rect 134422 135098 134604 135334
rect 134004 99654 134604 135098
rect 134004 99418 134186 99654
rect 134422 99418 134604 99654
rect 134004 99334 134604 99418
rect 134004 99098 134186 99334
rect 134422 99098 134604 99334
rect 134004 63654 134604 99098
rect 134004 63418 134186 63654
rect 134422 63418 134604 63654
rect 134004 63334 134604 63418
rect 134004 63098 134186 63334
rect 134422 63098 134604 63334
rect 134004 27654 134604 63098
rect 134004 27418 134186 27654
rect 134422 27418 134604 27654
rect 134004 27334 134604 27418
rect 134004 27098 134186 27334
rect 134422 27098 134604 27334
rect 134004 -4946 134604 27098
rect 134004 -5182 134186 -4946
rect 134422 -5182 134604 -4946
rect 134004 -5266 134604 -5182
rect 134004 -5502 134186 -5266
rect 134422 -5502 134604 -5266
rect 134004 -5524 134604 -5502
rect 137604 679254 138204 710722
rect 155604 710358 156204 711300
rect 155604 710122 155786 710358
rect 156022 710122 156204 710358
rect 155604 710038 156204 710122
rect 155604 709802 155786 710038
rect 156022 709802 156204 710038
rect 152004 708518 152604 709460
rect 152004 708282 152186 708518
rect 152422 708282 152604 708518
rect 152004 708198 152604 708282
rect 152004 707962 152186 708198
rect 152422 707962 152604 708198
rect 148404 706678 149004 707620
rect 148404 706442 148586 706678
rect 148822 706442 149004 706678
rect 148404 706358 149004 706442
rect 148404 706122 148586 706358
rect 148822 706122 149004 706358
rect 137604 679018 137786 679254
rect 138022 679018 138204 679254
rect 137604 678934 138204 679018
rect 137604 678698 137786 678934
rect 138022 678698 138204 678934
rect 137604 643254 138204 678698
rect 137604 643018 137786 643254
rect 138022 643018 138204 643254
rect 137604 642934 138204 643018
rect 137604 642698 137786 642934
rect 138022 642698 138204 642934
rect 137604 607254 138204 642698
rect 137604 607018 137786 607254
rect 138022 607018 138204 607254
rect 137604 606934 138204 607018
rect 137604 606698 137786 606934
rect 138022 606698 138204 606934
rect 137604 571254 138204 606698
rect 137604 571018 137786 571254
rect 138022 571018 138204 571254
rect 137604 570934 138204 571018
rect 137604 570698 137786 570934
rect 138022 570698 138204 570934
rect 137604 535254 138204 570698
rect 137604 535018 137786 535254
rect 138022 535018 138204 535254
rect 137604 534934 138204 535018
rect 137604 534698 137786 534934
rect 138022 534698 138204 534934
rect 137604 499254 138204 534698
rect 137604 499018 137786 499254
rect 138022 499018 138204 499254
rect 137604 498934 138204 499018
rect 137604 498698 137786 498934
rect 138022 498698 138204 498934
rect 137604 463254 138204 498698
rect 137604 463018 137786 463254
rect 138022 463018 138204 463254
rect 137604 462934 138204 463018
rect 137604 462698 137786 462934
rect 138022 462698 138204 462934
rect 137604 427254 138204 462698
rect 137604 427018 137786 427254
rect 138022 427018 138204 427254
rect 137604 426934 138204 427018
rect 137604 426698 137786 426934
rect 138022 426698 138204 426934
rect 137604 391254 138204 426698
rect 137604 391018 137786 391254
rect 138022 391018 138204 391254
rect 137604 390934 138204 391018
rect 137604 390698 137786 390934
rect 138022 390698 138204 390934
rect 137604 355254 138204 390698
rect 137604 355018 137786 355254
rect 138022 355018 138204 355254
rect 137604 354934 138204 355018
rect 137604 354698 137786 354934
rect 138022 354698 138204 354934
rect 137604 319254 138204 354698
rect 137604 319018 137786 319254
rect 138022 319018 138204 319254
rect 137604 318934 138204 319018
rect 137604 318698 137786 318934
rect 138022 318698 138204 318934
rect 137604 283254 138204 318698
rect 137604 283018 137786 283254
rect 138022 283018 138204 283254
rect 137604 282934 138204 283018
rect 137604 282698 137786 282934
rect 138022 282698 138204 282934
rect 137604 247254 138204 282698
rect 137604 247018 137786 247254
rect 138022 247018 138204 247254
rect 137604 246934 138204 247018
rect 137604 246698 137786 246934
rect 138022 246698 138204 246934
rect 137604 211254 138204 246698
rect 137604 211018 137786 211254
rect 138022 211018 138204 211254
rect 137604 210934 138204 211018
rect 137604 210698 137786 210934
rect 138022 210698 138204 210934
rect 137604 175254 138204 210698
rect 137604 175018 137786 175254
rect 138022 175018 138204 175254
rect 137604 174934 138204 175018
rect 137604 174698 137786 174934
rect 138022 174698 138204 174934
rect 137604 139254 138204 174698
rect 137604 139018 137786 139254
rect 138022 139018 138204 139254
rect 137604 138934 138204 139018
rect 137604 138698 137786 138934
rect 138022 138698 138204 138934
rect 137604 103254 138204 138698
rect 137604 103018 137786 103254
rect 138022 103018 138204 103254
rect 137604 102934 138204 103018
rect 137604 102698 137786 102934
rect 138022 102698 138204 102934
rect 137604 67254 138204 102698
rect 137604 67018 137786 67254
rect 138022 67018 138204 67254
rect 137604 66934 138204 67018
rect 137604 66698 137786 66934
rect 138022 66698 138204 66934
rect 137604 31254 138204 66698
rect 137604 31018 137786 31254
rect 138022 31018 138204 31254
rect 137604 30934 138204 31018
rect 137604 30698 137786 30934
rect 138022 30698 138204 30934
rect 119604 -6102 119786 -5866
rect 120022 -6102 120204 -5866
rect 119604 -6186 120204 -6102
rect 119604 -6422 119786 -6186
rect 120022 -6422 120204 -6186
rect 119604 -7364 120204 -6422
rect 137604 -6786 138204 30698
rect 144804 704838 145404 705780
rect 144804 704602 144986 704838
rect 145222 704602 145404 704838
rect 144804 704518 145404 704602
rect 144804 704282 144986 704518
rect 145222 704282 145404 704518
rect 144804 686454 145404 704282
rect 144804 686218 144986 686454
rect 145222 686218 145404 686454
rect 144804 686134 145404 686218
rect 144804 685898 144986 686134
rect 145222 685898 145404 686134
rect 144804 650454 145404 685898
rect 144804 650218 144986 650454
rect 145222 650218 145404 650454
rect 144804 650134 145404 650218
rect 144804 649898 144986 650134
rect 145222 649898 145404 650134
rect 144804 614454 145404 649898
rect 144804 614218 144986 614454
rect 145222 614218 145404 614454
rect 144804 614134 145404 614218
rect 144804 613898 144986 614134
rect 145222 613898 145404 614134
rect 144804 578454 145404 613898
rect 144804 578218 144986 578454
rect 145222 578218 145404 578454
rect 144804 578134 145404 578218
rect 144804 577898 144986 578134
rect 145222 577898 145404 578134
rect 144804 542454 145404 577898
rect 144804 542218 144986 542454
rect 145222 542218 145404 542454
rect 144804 542134 145404 542218
rect 144804 541898 144986 542134
rect 145222 541898 145404 542134
rect 144804 506454 145404 541898
rect 144804 506218 144986 506454
rect 145222 506218 145404 506454
rect 144804 506134 145404 506218
rect 144804 505898 144986 506134
rect 145222 505898 145404 506134
rect 144804 470454 145404 505898
rect 144804 470218 144986 470454
rect 145222 470218 145404 470454
rect 144804 470134 145404 470218
rect 144804 469898 144986 470134
rect 145222 469898 145404 470134
rect 144804 434454 145404 469898
rect 144804 434218 144986 434454
rect 145222 434218 145404 434454
rect 144804 434134 145404 434218
rect 144804 433898 144986 434134
rect 145222 433898 145404 434134
rect 144804 398454 145404 433898
rect 144804 398218 144986 398454
rect 145222 398218 145404 398454
rect 144804 398134 145404 398218
rect 144804 397898 144986 398134
rect 145222 397898 145404 398134
rect 144804 362454 145404 397898
rect 144804 362218 144986 362454
rect 145222 362218 145404 362454
rect 144804 362134 145404 362218
rect 144804 361898 144986 362134
rect 145222 361898 145404 362134
rect 144804 326454 145404 361898
rect 144804 326218 144986 326454
rect 145222 326218 145404 326454
rect 144804 326134 145404 326218
rect 144804 325898 144986 326134
rect 145222 325898 145404 326134
rect 144804 290454 145404 325898
rect 144804 290218 144986 290454
rect 145222 290218 145404 290454
rect 144804 290134 145404 290218
rect 144804 289898 144986 290134
rect 145222 289898 145404 290134
rect 144804 254454 145404 289898
rect 144804 254218 144986 254454
rect 145222 254218 145404 254454
rect 144804 254134 145404 254218
rect 144804 253898 144986 254134
rect 145222 253898 145404 254134
rect 144804 218454 145404 253898
rect 144804 218218 144986 218454
rect 145222 218218 145404 218454
rect 144804 218134 145404 218218
rect 144804 217898 144986 218134
rect 145222 217898 145404 218134
rect 144804 182454 145404 217898
rect 144804 182218 144986 182454
rect 145222 182218 145404 182454
rect 144804 182134 145404 182218
rect 144804 181898 144986 182134
rect 145222 181898 145404 182134
rect 144804 146454 145404 181898
rect 144804 146218 144986 146454
rect 145222 146218 145404 146454
rect 144804 146134 145404 146218
rect 144804 145898 144986 146134
rect 145222 145898 145404 146134
rect 144804 110454 145404 145898
rect 144804 110218 144986 110454
rect 145222 110218 145404 110454
rect 144804 110134 145404 110218
rect 144804 109898 144986 110134
rect 145222 109898 145404 110134
rect 144804 74454 145404 109898
rect 144804 74218 144986 74454
rect 145222 74218 145404 74454
rect 144804 74134 145404 74218
rect 144804 73898 144986 74134
rect 145222 73898 145404 74134
rect 144804 38454 145404 73898
rect 144804 38218 144986 38454
rect 145222 38218 145404 38454
rect 144804 38134 145404 38218
rect 144804 37898 144986 38134
rect 145222 37898 145404 38134
rect 144804 2454 145404 37898
rect 144804 2218 144986 2454
rect 145222 2218 145404 2454
rect 144804 2134 145404 2218
rect 144804 1898 144986 2134
rect 145222 1898 145404 2134
rect 144804 -346 145404 1898
rect 144804 -582 144986 -346
rect 145222 -582 145404 -346
rect 144804 -666 145404 -582
rect 144804 -902 144986 -666
rect 145222 -902 145404 -666
rect 144804 -1844 145404 -902
rect 148404 690054 149004 706122
rect 148404 689818 148586 690054
rect 148822 689818 149004 690054
rect 148404 689734 149004 689818
rect 148404 689498 148586 689734
rect 148822 689498 149004 689734
rect 148404 654054 149004 689498
rect 148404 653818 148586 654054
rect 148822 653818 149004 654054
rect 148404 653734 149004 653818
rect 148404 653498 148586 653734
rect 148822 653498 149004 653734
rect 148404 618054 149004 653498
rect 148404 617818 148586 618054
rect 148822 617818 149004 618054
rect 148404 617734 149004 617818
rect 148404 617498 148586 617734
rect 148822 617498 149004 617734
rect 148404 582054 149004 617498
rect 148404 581818 148586 582054
rect 148822 581818 149004 582054
rect 148404 581734 149004 581818
rect 148404 581498 148586 581734
rect 148822 581498 149004 581734
rect 148404 546054 149004 581498
rect 148404 545818 148586 546054
rect 148822 545818 149004 546054
rect 148404 545734 149004 545818
rect 148404 545498 148586 545734
rect 148822 545498 149004 545734
rect 148404 510054 149004 545498
rect 148404 509818 148586 510054
rect 148822 509818 149004 510054
rect 148404 509734 149004 509818
rect 148404 509498 148586 509734
rect 148822 509498 149004 509734
rect 148404 474054 149004 509498
rect 148404 473818 148586 474054
rect 148822 473818 149004 474054
rect 148404 473734 149004 473818
rect 148404 473498 148586 473734
rect 148822 473498 149004 473734
rect 148404 438054 149004 473498
rect 148404 437818 148586 438054
rect 148822 437818 149004 438054
rect 148404 437734 149004 437818
rect 148404 437498 148586 437734
rect 148822 437498 149004 437734
rect 148404 402054 149004 437498
rect 148404 401818 148586 402054
rect 148822 401818 149004 402054
rect 148404 401734 149004 401818
rect 148404 401498 148586 401734
rect 148822 401498 149004 401734
rect 148404 366054 149004 401498
rect 148404 365818 148586 366054
rect 148822 365818 149004 366054
rect 148404 365734 149004 365818
rect 148404 365498 148586 365734
rect 148822 365498 149004 365734
rect 148404 330054 149004 365498
rect 148404 329818 148586 330054
rect 148822 329818 149004 330054
rect 148404 329734 149004 329818
rect 148404 329498 148586 329734
rect 148822 329498 149004 329734
rect 148404 294054 149004 329498
rect 148404 293818 148586 294054
rect 148822 293818 149004 294054
rect 148404 293734 149004 293818
rect 148404 293498 148586 293734
rect 148822 293498 149004 293734
rect 148404 258054 149004 293498
rect 148404 257818 148586 258054
rect 148822 257818 149004 258054
rect 148404 257734 149004 257818
rect 148404 257498 148586 257734
rect 148822 257498 149004 257734
rect 148404 222054 149004 257498
rect 148404 221818 148586 222054
rect 148822 221818 149004 222054
rect 148404 221734 149004 221818
rect 148404 221498 148586 221734
rect 148822 221498 149004 221734
rect 148404 186054 149004 221498
rect 148404 185818 148586 186054
rect 148822 185818 149004 186054
rect 148404 185734 149004 185818
rect 148404 185498 148586 185734
rect 148822 185498 149004 185734
rect 148404 150054 149004 185498
rect 148404 149818 148586 150054
rect 148822 149818 149004 150054
rect 148404 149734 149004 149818
rect 148404 149498 148586 149734
rect 148822 149498 149004 149734
rect 148404 114054 149004 149498
rect 148404 113818 148586 114054
rect 148822 113818 149004 114054
rect 148404 113734 149004 113818
rect 148404 113498 148586 113734
rect 148822 113498 149004 113734
rect 148404 78054 149004 113498
rect 148404 77818 148586 78054
rect 148822 77818 149004 78054
rect 148404 77734 149004 77818
rect 148404 77498 148586 77734
rect 148822 77498 149004 77734
rect 148404 42054 149004 77498
rect 148404 41818 148586 42054
rect 148822 41818 149004 42054
rect 148404 41734 149004 41818
rect 148404 41498 148586 41734
rect 148822 41498 149004 41734
rect 148404 6054 149004 41498
rect 148404 5818 148586 6054
rect 148822 5818 149004 6054
rect 148404 5734 149004 5818
rect 148404 5498 148586 5734
rect 148822 5498 149004 5734
rect 148404 -2186 149004 5498
rect 148404 -2422 148586 -2186
rect 148822 -2422 149004 -2186
rect 148404 -2506 149004 -2422
rect 148404 -2742 148586 -2506
rect 148822 -2742 149004 -2506
rect 148404 -3684 149004 -2742
rect 152004 693654 152604 707962
rect 152004 693418 152186 693654
rect 152422 693418 152604 693654
rect 152004 693334 152604 693418
rect 152004 693098 152186 693334
rect 152422 693098 152604 693334
rect 152004 657654 152604 693098
rect 152004 657418 152186 657654
rect 152422 657418 152604 657654
rect 152004 657334 152604 657418
rect 152004 657098 152186 657334
rect 152422 657098 152604 657334
rect 152004 621654 152604 657098
rect 152004 621418 152186 621654
rect 152422 621418 152604 621654
rect 152004 621334 152604 621418
rect 152004 621098 152186 621334
rect 152422 621098 152604 621334
rect 152004 585654 152604 621098
rect 152004 585418 152186 585654
rect 152422 585418 152604 585654
rect 152004 585334 152604 585418
rect 152004 585098 152186 585334
rect 152422 585098 152604 585334
rect 152004 549654 152604 585098
rect 152004 549418 152186 549654
rect 152422 549418 152604 549654
rect 152004 549334 152604 549418
rect 152004 549098 152186 549334
rect 152422 549098 152604 549334
rect 152004 513654 152604 549098
rect 152004 513418 152186 513654
rect 152422 513418 152604 513654
rect 152004 513334 152604 513418
rect 152004 513098 152186 513334
rect 152422 513098 152604 513334
rect 152004 477654 152604 513098
rect 152004 477418 152186 477654
rect 152422 477418 152604 477654
rect 152004 477334 152604 477418
rect 152004 477098 152186 477334
rect 152422 477098 152604 477334
rect 152004 441654 152604 477098
rect 152004 441418 152186 441654
rect 152422 441418 152604 441654
rect 152004 441334 152604 441418
rect 152004 441098 152186 441334
rect 152422 441098 152604 441334
rect 152004 405654 152604 441098
rect 152004 405418 152186 405654
rect 152422 405418 152604 405654
rect 152004 405334 152604 405418
rect 152004 405098 152186 405334
rect 152422 405098 152604 405334
rect 152004 369654 152604 405098
rect 152004 369418 152186 369654
rect 152422 369418 152604 369654
rect 152004 369334 152604 369418
rect 152004 369098 152186 369334
rect 152422 369098 152604 369334
rect 152004 333654 152604 369098
rect 152004 333418 152186 333654
rect 152422 333418 152604 333654
rect 152004 333334 152604 333418
rect 152004 333098 152186 333334
rect 152422 333098 152604 333334
rect 152004 297654 152604 333098
rect 152004 297418 152186 297654
rect 152422 297418 152604 297654
rect 152004 297334 152604 297418
rect 152004 297098 152186 297334
rect 152422 297098 152604 297334
rect 152004 261654 152604 297098
rect 152004 261418 152186 261654
rect 152422 261418 152604 261654
rect 152004 261334 152604 261418
rect 152004 261098 152186 261334
rect 152422 261098 152604 261334
rect 152004 225654 152604 261098
rect 152004 225418 152186 225654
rect 152422 225418 152604 225654
rect 152004 225334 152604 225418
rect 152004 225098 152186 225334
rect 152422 225098 152604 225334
rect 152004 189654 152604 225098
rect 152004 189418 152186 189654
rect 152422 189418 152604 189654
rect 152004 189334 152604 189418
rect 152004 189098 152186 189334
rect 152422 189098 152604 189334
rect 152004 153654 152604 189098
rect 152004 153418 152186 153654
rect 152422 153418 152604 153654
rect 152004 153334 152604 153418
rect 152004 153098 152186 153334
rect 152422 153098 152604 153334
rect 152004 117654 152604 153098
rect 152004 117418 152186 117654
rect 152422 117418 152604 117654
rect 152004 117334 152604 117418
rect 152004 117098 152186 117334
rect 152422 117098 152604 117334
rect 152004 81654 152604 117098
rect 152004 81418 152186 81654
rect 152422 81418 152604 81654
rect 152004 81334 152604 81418
rect 152004 81098 152186 81334
rect 152422 81098 152604 81334
rect 152004 45654 152604 81098
rect 152004 45418 152186 45654
rect 152422 45418 152604 45654
rect 152004 45334 152604 45418
rect 152004 45098 152186 45334
rect 152422 45098 152604 45334
rect 152004 9654 152604 45098
rect 152004 9418 152186 9654
rect 152422 9418 152604 9654
rect 152004 9334 152604 9418
rect 152004 9098 152186 9334
rect 152422 9098 152604 9334
rect 152004 -4026 152604 9098
rect 152004 -4262 152186 -4026
rect 152422 -4262 152604 -4026
rect 152004 -4346 152604 -4262
rect 152004 -4582 152186 -4346
rect 152422 -4582 152604 -4346
rect 152004 -5524 152604 -4582
rect 155604 697254 156204 709802
rect 173604 711278 174204 711300
rect 173604 711042 173786 711278
rect 174022 711042 174204 711278
rect 173604 710958 174204 711042
rect 173604 710722 173786 710958
rect 174022 710722 174204 710958
rect 170004 709438 170604 709460
rect 170004 709202 170186 709438
rect 170422 709202 170604 709438
rect 170004 709118 170604 709202
rect 170004 708882 170186 709118
rect 170422 708882 170604 709118
rect 166404 707598 167004 707620
rect 166404 707362 166586 707598
rect 166822 707362 167004 707598
rect 166404 707278 167004 707362
rect 166404 707042 166586 707278
rect 166822 707042 167004 707278
rect 155604 697018 155786 697254
rect 156022 697018 156204 697254
rect 155604 696934 156204 697018
rect 155604 696698 155786 696934
rect 156022 696698 156204 696934
rect 155604 661254 156204 696698
rect 155604 661018 155786 661254
rect 156022 661018 156204 661254
rect 155604 660934 156204 661018
rect 155604 660698 155786 660934
rect 156022 660698 156204 660934
rect 155604 625254 156204 660698
rect 155604 625018 155786 625254
rect 156022 625018 156204 625254
rect 155604 624934 156204 625018
rect 155604 624698 155786 624934
rect 156022 624698 156204 624934
rect 155604 589254 156204 624698
rect 155604 589018 155786 589254
rect 156022 589018 156204 589254
rect 155604 588934 156204 589018
rect 155604 588698 155786 588934
rect 156022 588698 156204 588934
rect 155604 553254 156204 588698
rect 155604 553018 155786 553254
rect 156022 553018 156204 553254
rect 155604 552934 156204 553018
rect 155604 552698 155786 552934
rect 156022 552698 156204 552934
rect 155604 517254 156204 552698
rect 155604 517018 155786 517254
rect 156022 517018 156204 517254
rect 155604 516934 156204 517018
rect 155604 516698 155786 516934
rect 156022 516698 156204 516934
rect 155604 481254 156204 516698
rect 155604 481018 155786 481254
rect 156022 481018 156204 481254
rect 155604 480934 156204 481018
rect 155604 480698 155786 480934
rect 156022 480698 156204 480934
rect 155604 445254 156204 480698
rect 155604 445018 155786 445254
rect 156022 445018 156204 445254
rect 155604 444934 156204 445018
rect 155604 444698 155786 444934
rect 156022 444698 156204 444934
rect 155604 409254 156204 444698
rect 155604 409018 155786 409254
rect 156022 409018 156204 409254
rect 155604 408934 156204 409018
rect 155604 408698 155786 408934
rect 156022 408698 156204 408934
rect 155604 373254 156204 408698
rect 155604 373018 155786 373254
rect 156022 373018 156204 373254
rect 155604 372934 156204 373018
rect 155604 372698 155786 372934
rect 156022 372698 156204 372934
rect 155604 337254 156204 372698
rect 155604 337018 155786 337254
rect 156022 337018 156204 337254
rect 155604 336934 156204 337018
rect 155604 336698 155786 336934
rect 156022 336698 156204 336934
rect 155604 301254 156204 336698
rect 155604 301018 155786 301254
rect 156022 301018 156204 301254
rect 155604 300934 156204 301018
rect 155604 300698 155786 300934
rect 156022 300698 156204 300934
rect 155604 265254 156204 300698
rect 155604 265018 155786 265254
rect 156022 265018 156204 265254
rect 155604 264934 156204 265018
rect 155604 264698 155786 264934
rect 156022 264698 156204 264934
rect 155604 229254 156204 264698
rect 155604 229018 155786 229254
rect 156022 229018 156204 229254
rect 155604 228934 156204 229018
rect 155604 228698 155786 228934
rect 156022 228698 156204 228934
rect 155604 193254 156204 228698
rect 155604 193018 155786 193254
rect 156022 193018 156204 193254
rect 155604 192934 156204 193018
rect 155604 192698 155786 192934
rect 156022 192698 156204 192934
rect 155604 157254 156204 192698
rect 155604 157018 155786 157254
rect 156022 157018 156204 157254
rect 155604 156934 156204 157018
rect 155604 156698 155786 156934
rect 156022 156698 156204 156934
rect 155604 121254 156204 156698
rect 155604 121018 155786 121254
rect 156022 121018 156204 121254
rect 155604 120934 156204 121018
rect 155604 120698 155786 120934
rect 156022 120698 156204 120934
rect 155604 85254 156204 120698
rect 155604 85018 155786 85254
rect 156022 85018 156204 85254
rect 155604 84934 156204 85018
rect 155604 84698 155786 84934
rect 156022 84698 156204 84934
rect 155604 49254 156204 84698
rect 155604 49018 155786 49254
rect 156022 49018 156204 49254
rect 155604 48934 156204 49018
rect 155604 48698 155786 48934
rect 156022 48698 156204 48934
rect 155604 13254 156204 48698
rect 155604 13018 155786 13254
rect 156022 13018 156204 13254
rect 155604 12934 156204 13018
rect 155604 12698 155786 12934
rect 156022 12698 156204 12934
rect 137604 -7022 137786 -6786
rect 138022 -7022 138204 -6786
rect 137604 -7106 138204 -7022
rect 137604 -7342 137786 -7106
rect 138022 -7342 138204 -7106
rect 137604 -7364 138204 -7342
rect 155604 -5866 156204 12698
rect 162804 705758 163404 705780
rect 162804 705522 162986 705758
rect 163222 705522 163404 705758
rect 162804 705438 163404 705522
rect 162804 705202 162986 705438
rect 163222 705202 163404 705438
rect 162804 668454 163404 705202
rect 162804 668218 162986 668454
rect 163222 668218 163404 668454
rect 162804 668134 163404 668218
rect 162804 667898 162986 668134
rect 163222 667898 163404 668134
rect 162804 632454 163404 667898
rect 162804 632218 162986 632454
rect 163222 632218 163404 632454
rect 162804 632134 163404 632218
rect 162804 631898 162986 632134
rect 163222 631898 163404 632134
rect 162804 596454 163404 631898
rect 162804 596218 162986 596454
rect 163222 596218 163404 596454
rect 162804 596134 163404 596218
rect 162804 595898 162986 596134
rect 163222 595898 163404 596134
rect 162804 560454 163404 595898
rect 162804 560218 162986 560454
rect 163222 560218 163404 560454
rect 162804 560134 163404 560218
rect 162804 559898 162986 560134
rect 163222 559898 163404 560134
rect 162804 524454 163404 559898
rect 162804 524218 162986 524454
rect 163222 524218 163404 524454
rect 162804 524134 163404 524218
rect 162804 523898 162986 524134
rect 163222 523898 163404 524134
rect 162804 488454 163404 523898
rect 162804 488218 162986 488454
rect 163222 488218 163404 488454
rect 162804 488134 163404 488218
rect 162804 487898 162986 488134
rect 163222 487898 163404 488134
rect 162804 452454 163404 487898
rect 162804 452218 162986 452454
rect 163222 452218 163404 452454
rect 162804 452134 163404 452218
rect 162804 451898 162986 452134
rect 163222 451898 163404 452134
rect 162804 416454 163404 451898
rect 162804 416218 162986 416454
rect 163222 416218 163404 416454
rect 162804 416134 163404 416218
rect 162804 415898 162986 416134
rect 163222 415898 163404 416134
rect 162804 380454 163404 415898
rect 162804 380218 162986 380454
rect 163222 380218 163404 380454
rect 162804 380134 163404 380218
rect 162804 379898 162986 380134
rect 163222 379898 163404 380134
rect 162804 344454 163404 379898
rect 162804 344218 162986 344454
rect 163222 344218 163404 344454
rect 162804 344134 163404 344218
rect 162804 343898 162986 344134
rect 163222 343898 163404 344134
rect 162804 308454 163404 343898
rect 162804 308218 162986 308454
rect 163222 308218 163404 308454
rect 162804 308134 163404 308218
rect 162804 307898 162986 308134
rect 163222 307898 163404 308134
rect 162804 272454 163404 307898
rect 162804 272218 162986 272454
rect 163222 272218 163404 272454
rect 162804 272134 163404 272218
rect 162804 271898 162986 272134
rect 163222 271898 163404 272134
rect 162804 236454 163404 271898
rect 162804 236218 162986 236454
rect 163222 236218 163404 236454
rect 162804 236134 163404 236218
rect 162804 235898 162986 236134
rect 163222 235898 163404 236134
rect 162804 200454 163404 235898
rect 162804 200218 162986 200454
rect 163222 200218 163404 200454
rect 162804 200134 163404 200218
rect 162804 199898 162986 200134
rect 163222 199898 163404 200134
rect 162804 164454 163404 199898
rect 162804 164218 162986 164454
rect 163222 164218 163404 164454
rect 162804 164134 163404 164218
rect 162804 163898 162986 164134
rect 163222 163898 163404 164134
rect 162804 128454 163404 163898
rect 162804 128218 162986 128454
rect 163222 128218 163404 128454
rect 162804 128134 163404 128218
rect 162804 127898 162986 128134
rect 163222 127898 163404 128134
rect 162804 92454 163404 127898
rect 162804 92218 162986 92454
rect 163222 92218 163404 92454
rect 162804 92134 163404 92218
rect 162804 91898 162986 92134
rect 163222 91898 163404 92134
rect 162804 56454 163404 91898
rect 162804 56218 162986 56454
rect 163222 56218 163404 56454
rect 162804 56134 163404 56218
rect 162804 55898 162986 56134
rect 163222 55898 163404 56134
rect 162804 20454 163404 55898
rect 162804 20218 162986 20454
rect 163222 20218 163404 20454
rect 162804 20134 163404 20218
rect 162804 19898 162986 20134
rect 163222 19898 163404 20134
rect 162804 -1266 163404 19898
rect 162804 -1502 162986 -1266
rect 163222 -1502 163404 -1266
rect 162804 -1586 163404 -1502
rect 162804 -1822 162986 -1586
rect 163222 -1822 163404 -1586
rect 162804 -1844 163404 -1822
rect 166404 672054 167004 707042
rect 166404 671818 166586 672054
rect 166822 671818 167004 672054
rect 166404 671734 167004 671818
rect 166404 671498 166586 671734
rect 166822 671498 167004 671734
rect 166404 636054 167004 671498
rect 166404 635818 166586 636054
rect 166822 635818 167004 636054
rect 166404 635734 167004 635818
rect 166404 635498 166586 635734
rect 166822 635498 167004 635734
rect 166404 600054 167004 635498
rect 166404 599818 166586 600054
rect 166822 599818 167004 600054
rect 166404 599734 167004 599818
rect 166404 599498 166586 599734
rect 166822 599498 167004 599734
rect 166404 564054 167004 599498
rect 166404 563818 166586 564054
rect 166822 563818 167004 564054
rect 166404 563734 167004 563818
rect 166404 563498 166586 563734
rect 166822 563498 167004 563734
rect 166404 528054 167004 563498
rect 166404 527818 166586 528054
rect 166822 527818 167004 528054
rect 166404 527734 167004 527818
rect 166404 527498 166586 527734
rect 166822 527498 167004 527734
rect 166404 492054 167004 527498
rect 166404 491818 166586 492054
rect 166822 491818 167004 492054
rect 166404 491734 167004 491818
rect 166404 491498 166586 491734
rect 166822 491498 167004 491734
rect 166404 456054 167004 491498
rect 166404 455818 166586 456054
rect 166822 455818 167004 456054
rect 166404 455734 167004 455818
rect 166404 455498 166586 455734
rect 166822 455498 167004 455734
rect 166404 420054 167004 455498
rect 166404 419818 166586 420054
rect 166822 419818 167004 420054
rect 166404 419734 167004 419818
rect 166404 419498 166586 419734
rect 166822 419498 167004 419734
rect 166404 384054 167004 419498
rect 166404 383818 166586 384054
rect 166822 383818 167004 384054
rect 166404 383734 167004 383818
rect 166404 383498 166586 383734
rect 166822 383498 167004 383734
rect 166404 348054 167004 383498
rect 166404 347818 166586 348054
rect 166822 347818 167004 348054
rect 166404 347734 167004 347818
rect 166404 347498 166586 347734
rect 166822 347498 167004 347734
rect 166404 312054 167004 347498
rect 166404 311818 166586 312054
rect 166822 311818 167004 312054
rect 166404 311734 167004 311818
rect 166404 311498 166586 311734
rect 166822 311498 167004 311734
rect 166404 276054 167004 311498
rect 166404 275818 166586 276054
rect 166822 275818 167004 276054
rect 166404 275734 167004 275818
rect 166404 275498 166586 275734
rect 166822 275498 167004 275734
rect 166404 240054 167004 275498
rect 166404 239818 166586 240054
rect 166822 239818 167004 240054
rect 166404 239734 167004 239818
rect 166404 239498 166586 239734
rect 166822 239498 167004 239734
rect 166404 204054 167004 239498
rect 166404 203818 166586 204054
rect 166822 203818 167004 204054
rect 166404 203734 167004 203818
rect 166404 203498 166586 203734
rect 166822 203498 167004 203734
rect 166404 168054 167004 203498
rect 166404 167818 166586 168054
rect 166822 167818 167004 168054
rect 166404 167734 167004 167818
rect 166404 167498 166586 167734
rect 166822 167498 167004 167734
rect 166404 132054 167004 167498
rect 166404 131818 166586 132054
rect 166822 131818 167004 132054
rect 166404 131734 167004 131818
rect 166404 131498 166586 131734
rect 166822 131498 167004 131734
rect 166404 96054 167004 131498
rect 166404 95818 166586 96054
rect 166822 95818 167004 96054
rect 166404 95734 167004 95818
rect 166404 95498 166586 95734
rect 166822 95498 167004 95734
rect 166404 60054 167004 95498
rect 166404 59818 166586 60054
rect 166822 59818 167004 60054
rect 166404 59734 167004 59818
rect 166404 59498 166586 59734
rect 166822 59498 167004 59734
rect 166404 24054 167004 59498
rect 166404 23818 166586 24054
rect 166822 23818 167004 24054
rect 166404 23734 167004 23818
rect 166404 23498 166586 23734
rect 166822 23498 167004 23734
rect 166404 -3106 167004 23498
rect 166404 -3342 166586 -3106
rect 166822 -3342 167004 -3106
rect 166404 -3426 167004 -3342
rect 166404 -3662 166586 -3426
rect 166822 -3662 167004 -3426
rect 166404 -3684 167004 -3662
rect 170004 675654 170604 708882
rect 170004 675418 170186 675654
rect 170422 675418 170604 675654
rect 170004 675334 170604 675418
rect 170004 675098 170186 675334
rect 170422 675098 170604 675334
rect 170004 639654 170604 675098
rect 170004 639418 170186 639654
rect 170422 639418 170604 639654
rect 170004 639334 170604 639418
rect 170004 639098 170186 639334
rect 170422 639098 170604 639334
rect 170004 603654 170604 639098
rect 170004 603418 170186 603654
rect 170422 603418 170604 603654
rect 170004 603334 170604 603418
rect 170004 603098 170186 603334
rect 170422 603098 170604 603334
rect 170004 567654 170604 603098
rect 170004 567418 170186 567654
rect 170422 567418 170604 567654
rect 170004 567334 170604 567418
rect 170004 567098 170186 567334
rect 170422 567098 170604 567334
rect 170004 531654 170604 567098
rect 170004 531418 170186 531654
rect 170422 531418 170604 531654
rect 170004 531334 170604 531418
rect 170004 531098 170186 531334
rect 170422 531098 170604 531334
rect 170004 495654 170604 531098
rect 173604 679254 174204 710722
rect 191604 710358 192204 711300
rect 191604 710122 191786 710358
rect 192022 710122 192204 710358
rect 191604 710038 192204 710122
rect 191604 709802 191786 710038
rect 192022 709802 192204 710038
rect 188004 708518 188604 709460
rect 188004 708282 188186 708518
rect 188422 708282 188604 708518
rect 188004 708198 188604 708282
rect 188004 707962 188186 708198
rect 188422 707962 188604 708198
rect 184404 706678 185004 707620
rect 184404 706442 184586 706678
rect 184822 706442 185004 706678
rect 184404 706358 185004 706442
rect 184404 706122 184586 706358
rect 184822 706122 185004 706358
rect 173604 679018 173786 679254
rect 174022 679018 174204 679254
rect 173604 678934 174204 679018
rect 173604 678698 173786 678934
rect 174022 678698 174204 678934
rect 173604 643254 174204 678698
rect 173604 643018 173786 643254
rect 174022 643018 174204 643254
rect 173604 642934 174204 643018
rect 173604 642698 173786 642934
rect 174022 642698 174204 642934
rect 173604 607254 174204 642698
rect 173604 607018 173786 607254
rect 174022 607018 174204 607254
rect 173604 606934 174204 607018
rect 173604 606698 173786 606934
rect 174022 606698 174204 606934
rect 173604 571254 174204 606698
rect 173604 571018 173786 571254
rect 174022 571018 174204 571254
rect 173604 570934 174204 571018
rect 173604 570698 173786 570934
rect 174022 570698 174204 570934
rect 173604 535254 174204 570698
rect 173604 535018 173786 535254
rect 174022 535018 174204 535254
rect 173604 534934 174204 535018
rect 173604 534698 173786 534934
rect 174022 534698 174204 534934
rect 173387 519348 173453 519349
rect 173387 519284 173388 519348
rect 173452 519284 173453 519348
rect 173387 519283 173453 519284
rect 170004 495418 170186 495654
rect 170422 495418 170604 495654
rect 170004 495334 170604 495418
rect 170004 495098 170186 495334
rect 170422 495098 170604 495334
rect 170004 459654 170604 495098
rect 170004 459418 170186 459654
rect 170422 459418 170604 459654
rect 170004 459334 170604 459418
rect 170004 459098 170186 459334
rect 170422 459098 170604 459334
rect 170004 423654 170604 459098
rect 170004 423418 170186 423654
rect 170422 423418 170604 423654
rect 170004 423334 170604 423418
rect 170004 423098 170186 423334
rect 170422 423098 170604 423334
rect 170004 387654 170604 423098
rect 170004 387418 170186 387654
rect 170422 387418 170604 387654
rect 170004 387334 170604 387418
rect 170004 387098 170186 387334
rect 170422 387098 170604 387334
rect 170004 351654 170604 387098
rect 170004 351418 170186 351654
rect 170422 351418 170604 351654
rect 170004 351334 170604 351418
rect 170004 351098 170186 351334
rect 170422 351098 170604 351334
rect 170004 315654 170604 351098
rect 170004 315418 170186 315654
rect 170422 315418 170604 315654
rect 170004 315334 170604 315418
rect 170004 315098 170186 315334
rect 170422 315098 170604 315334
rect 170004 279654 170604 315098
rect 170004 279418 170186 279654
rect 170422 279418 170604 279654
rect 170004 279334 170604 279418
rect 170004 279098 170186 279334
rect 170422 279098 170604 279334
rect 170004 243654 170604 279098
rect 170004 243418 170186 243654
rect 170422 243418 170604 243654
rect 170004 243334 170604 243418
rect 170004 243098 170186 243334
rect 170422 243098 170604 243334
rect 170004 207654 170604 243098
rect 170004 207418 170186 207654
rect 170422 207418 170604 207654
rect 170004 207334 170604 207418
rect 170004 207098 170186 207334
rect 170422 207098 170604 207334
rect 170004 171654 170604 207098
rect 170004 171418 170186 171654
rect 170422 171418 170604 171654
rect 170004 171334 170604 171418
rect 170004 171098 170186 171334
rect 170422 171098 170604 171334
rect 170004 135654 170604 171098
rect 170004 135418 170186 135654
rect 170422 135418 170604 135654
rect 170004 135334 170604 135418
rect 170004 135098 170186 135334
rect 170422 135098 170604 135334
rect 170004 99654 170604 135098
rect 170004 99418 170186 99654
rect 170422 99418 170604 99654
rect 170004 99334 170604 99418
rect 170004 99098 170186 99334
rect 170422 99098 170604 99334
rect 170004 63654 170604 99098
rect 170004 63418 170186 63654
rect 170422 63418 170604 63654
rect 170004 63334 170604 63418
rect 170004 63098 170186 63334
rect 170422 63098 170604 63334
rect 170004 27654 170604 63098
rect 173390 40357 173450 519283
rect 173604 499254 174204 534698
rect 180804 704838 181404 705780
rect 180804 704602 180986 704838
rect 181222 704602 181404 704838
rect 180804 704518 181404 704602
rect 180804 704282 180986 704518
rect 181222 704282 181404 704518
rect 180804 686454 181404 704282
rect 180804 686218 180986 686454
rect 181222 686218 181404 686454
rect 180804 686134 181404 686218
rect 180804 685898 180986 686134
rect 181222 685898 181404 686134
rect 180804 650454 181404 685898
rect 180804 650218 180986 650454
rect 181222 650218 181404 650454
rect 180804 650134 181404 650218
rect 180804 649898 180986 650134
rect 181222 649898 181404 650134
rect 180804 614454 181404 649898
rect 180804 614218 180986 614454
rect 181222 614218 181404 614454
rect 180804 614134 181404 614218
rect 180804 613898 180986 614134
rect 181222 613898 181404 614134
rect 180804 578454 181404 613898
rect 180804 578218 180986 578454
rect 181222 578218 181404 578454
rect 180804 578134 181404 578218
rect 180804 577898 180986 578134
rect 181222 577898 181404 578134
rect 180804 542454 181404 577898
rect 180804 542218 180986 542454
rect 181222 542218 181404 542454
rect 180804 542134 181404 542218
rect 180804 541898 180986 542134
rect 181222 541898 181404 542134
rect 176515 517988 176581 517989
rect 176515 517924 176516 517988
rect 176580 517924 176581 517988
rect 176515 517923 176581 517924
rect 176699 517988 176765 517989
rect 176699 517924 176700 517988
rect 176764 517924 176765 517988
rect 176699 517923 176765 517924
rect 176518 517850 176578 517923
rect 176702 517850 176762 517923
rect 176518 517790 176762 517850
rect 173604 499018 173786 499254
rect 174022 499018 174204 499254
rect 173604 498934 174204 499018
rect 173604 498698 173786 498934
rect 174022 498698 174204 498934
rect 173604 463254 174204 498698
rect 173604 463018 173786 463254
rect 174022 463018 174204 463254
rect 173604 462934 174204 463018
rect 173604 462698 173786 462934
rect 174022 462698 174204 462934
rect 173604 427254 174204 462698
rect 173604 427018 173786 427254
rect 174022 427018 174204 427254
rect 173604 426934 174204 427018
rect 173604 426698 173786 426934
rect 174022 426698 174204 426934
rect 173604 391254 174204 426698
rect 173604 391018 173786 391254
rect 174022 391018 174204 391254
rect 173604 390934 174204 391018
rect 173604 390698 173786 390934
rect 174022 390698 174204 390934
rect 173604 355254 174204 390698
rect 173604 355018 173786 355254
rect 174022 355018 174204 355254
rect 173604 354934 174204 355018
rect 173604 354698 173786 354934
rect 174022 354698 174204 354934
rect 173604 319254 174204 354698
rect 173604 319018 173786 319254
rect 174022 319018 174204 319254
rect 173604 318934 174204 319018
rect 173604 318698 173786 318934
rect 174022 318698 174204 318934
rect 173604 283254 174204 318698
rect 173604 283018 173786 283254
rect 174022 283018 174204 283254
rect 173604 282934 174204 283018
rect 173604 282698 173786 282934
rect 174022 282698 174204 282934
rect 173604 247254 174204 282698
rect 173604 247018 173786 247254
rect 174022 247018 174204 247254
rect 173604 246934 174204 247018
rect 173604 246698 173786 246934
rect 174022 246698 174204 246934
rect 173604 211254 174204 246698
rect 173604 211018 173786 211254
rect 174022 211018 174204 211254
rect 173604 210934 174204 211018
rect 173604 210698 173786 210934
rect 174022 210698 174204 210934
rect 173604 175254 174204 210698
rect 173604 175018 173786 175254
rect 174022 175018 174204 175254
rect 173604 174934 174204 175018
rect 173604 174698 173786 174934
rect 174022 174698 174204 174934
rect 173604 139254 174204 174698
rect 173604 139018 173786 139254
rect 174022 139018 174204 139254
rect 173604 138934 174204 139018
rect 173604 138698 173786 138934
rect 174022 138698 174204 138934
rect 173604 103254 174204 138698
rect 173604 103018 173786 103254
rect 174022 103018 174204 103254
rect 173604 102934 174204 103018
rect 173604 102698 173786 102934
rect 174022 102698 174204 102934
rect 173604 67254 174204 102698
rect 173604 67018 173786 67254
rect 174022 67018 174204 67254
rect 173604 66934 174204 67018
rect 173604 66698 173786 66934
rect 174022 66698 174204 66934
rect 173387 40356 173453 40357
rect 173387 40292 173388 40356
rect 173452 40292 173453 40356
rect 173387 40291 173453 40292
rect 170004 27418 170186 27654
rect 170422 27418 170604 27654
rect 170004 27334 170604 27418
rect 170004 27098 170186 27334
rect 170422 27098 170604 27334
rect 170004 -4946 170604 27098
rect 170004 -5182 170186 -4946
rect 170422 -5182 170604 -4946
rect 170004 -5266 170604 -5182
rect 170004 -5502 170186 -5266
rect 170422 -5502 170604 -5266
rect 170004 -5524 170604 -5502
rect 173604 31254 174204 66698
rect 173604 31018 173786 31254
rect 174022 31018 174204 31254
rect 173604 30934 174204 31018
rect 173604 30698 173786 30934
rect 174022 30698 174204 30934
rect 155604 -6102 155786 -5866
rect 156022 -6102 156204 -5866
rect 155604 -6186 156204 -6102
rect 155604 -6422 155786 -6186
rect 156022 -6422 156204 -6186
rect 155604 -7364 156204 -6422
rect 173604 -6786 174204 30698
rect 180804 506454 181404 541898
rect 184404 690054 185004 706122
rect 184404 689818 184586 690054
rect 184822 689818 185004 690054
rect 184404 689734 185004 689818
rect 184404 689498 184586 689734
rect 184822 689498 185004 689734
rect 184404 654054 185004 689498
rect 184404 653818 184586 654054
rect 184822 653818 185004 654054
rect 184404 653734 185004 653818
rect 184404 653498 184586 653734
rect 184822 653498 185004 653734
rect 184404 618054 185004 653498
rect 184404 617818 184586 618054
rect 184822 617818 185004 618054
rect 184404 617734 185004 617818
rect 184404 617498 184586 617734
rect 184822 617498 185004 617734
rect 184404 582054 185004 617498
rect 184404 581818 184586 582054
rect 184822 581818 185004 582054
rect 184404 581734 185004 581818
rect 184404 581498 184586 581734
rect 184822 581498 185004 581734
rect 184404 546054 185004 581498
rect 184404 545818 184586 546054
rect 184822 545818 185004 546054
rect 184404 545734 185004 545818
rect 184404 545498 184586 545734
rect 184822 545498 185004 545734
rect 182219 518532 182285 518533
rect 182219 518468 182220 518532
rect 182284 518468 182285 518532
rect 182219 518467 182285 518468
rect 182222 517989 182282 518467
rect 182219 517988 182285 517989
rect 182219 517924 182220 517988
rect 182284 517924 182285 517988
rect 182219 517923 182285 517924
rect 180804 506218 180986 506454
rect 181222 506218 181404 506454
rect 180804 506134 181404 506218
rect 180804 505898 180986 506134
rect 181222 505898 181404 506134
rect 180804 470454 181404 505898
rect 180804 470218 180986 470454
rect 181222 470218 181404 470454
rect 180804 470134 181404 470218
rect 180804 469898 180986 470134
rect 181222 469898 181404 470134
rect 180804 434454 181404 469898
rect 180804 434218 180986 434454
rect 181222 434218 181404 434454
rect 180804 434134 181404 434218
rect 180804 433898 180986 434134
rect 181222 433898 181404 434134
rect 180804 398454 181404 433898
rect 180804 398218 180986 398454
rect 181222 398218 181404 398454
rect 180804 398134 181404 398218
rect 180804 397898 180986 398134
rect 181222 397898 181404 398134
rect 180804 362454 181404 397898
rect 180804 362218 180986 362454
rect 181222 362218 181404 362454
rect 180804 362134 181404 362218
rect 180804 361898 180986 362134
rect 181222 361898 181404 362134
rect 180804 326454 181404 361898
rect 180804 326218 180986 326454
rect 181222 326218 181404 326454
rect 180804 326134 181404 326218
rect 180804 325898 180986 326134
rect 181222 325898 181404 326134
rect 180804 290454 181404 325898
rect 180804 290218 180986 290454
rect 181222 290218 181404 290454
rect 180804 290134 181404 290218
rect 180804 289898 180986 290134
rect 181222 289898 181404 290134
rect 180804 254454 181404 289898
rect 180804 254218 180986 254454
rect 181222 254218 181404 254454
rect 180804 254134 181404 254218
rect 180804 253898 180986 254134
rect 181222 253898 181404 254134
rect 180804 218454 181404 253898
rect 180804 218218 180986 218454
rect 181222 218218 181404 218454
rect 180804 218134 181404 218218
rect 180804 217898 180986 218134
rect 181222 217898 181404 218134
rect 180804 182454 181404 217898
rect 180804 182218 180986 182454
rect 181222 182218 181404 182454
rect 180804 182134 181404 182218
rect 180804 181898 180986 182134
rect 181222 181898 181404 182134
rect 180804 146454 181404 181898
rect 180804 146218 180986 146454
rect 181222 146218 181404 146454
rect 180804 146134 181404 146218
rect 180804 145898 180986 146134
rect 181222 145898 181404 146134
rect 180804 110454 181404 145898
rect 180804 110218 180986 110454
rect 181222 110218 181404 110454
rect 180804 110134 181404 110218
rect 180804 109898 180986 110134
rect 181222 109898 181404 110134
rect 180804 74454 181404 109898
rect 180804 74218 180986 74454
rect 181222 74218 181404 74454
rect 180804 74134 181404 74218
rect 180804 73898 180986 74134
rect 181222 73898 181404 74134
rect 180804 38454 181404 73898
rect 180804 38218 180986 38454
rect 181222 38218 181404 38454
rect 180804 38134 181404 38218
rect 180804 37898 180986 38134
rect 181222 37898 181404 38134
rect 180804 2454 181404 37898
rect 180804 2218 180986 2454
rect 181222 2218 181404 2454
rect 180804 2134 181404 2218
rect 180804 1898 180986 2134
rect 181222 1898 181404 2134
rect 180804 -346 181404 1898
rect 180804 -582 180986 -346
rect 181222 -582 181404 -346
rect 180804 -666 181404 -582
rect 180804 -902 180986 -666
rect 181222 -902 181404 -666
rect 180804 -1844 181404 -902
rect 184404 510054 185004 545498
rect 184404 509818 184586 510054
rect 184822 509818 185004 510054
rect 184404 509734 185004 509818
rect 184404 509498 184586 509734
rect 184822 509498 185004 509734
rect 184404 474054 185004 509498
rect 184404 473818 184586 474054
rect 184822 473818 185004 474054
rect 184404 473734 185004 473818
rect 184404 473498 184586 473734
rect 184822 473498 185004 473734
rect 184404 438054 185004 473498
rect 184404 437818 184586 438054
rect 184822 437818 185004 438054
rect 184404 437734 185004 437818
rect 184404 437498 184586 437734
rect 184822 437498 185004 437734
rect 184404 402054 185004 437498
rect 184404 401818 184586 402054
rect 184822 401818 185004 402054
rect 184404 401734 185004 401818
rect 184404 401498 184586 401734
rect 184822 401498 185004 401734
rect 184404 366054 185004 401498
rect 184404 365818 184586 366054
rect 184822 365818 185004 366054
rect 184404 365734 185004 365818
rect 184404 365498 184586 365734
rect 184822 365498 185004 365734
rect 184404 330054 185004 365498
rect 184404 329818 184586 330054
rect 184822 329818 185004 330054
rect 184404 329734 185004 329818
rect 184404 329498 184586 329734
rect 184822 329498 185004 329734
rect 184404 294054 185004 329498
rect 184404 293818 184586 294054
rect 184822 293818 185004 294054
rect 184404 293734 185004 293818
rect 184404 293498 184586 293734
rect 184822 293498 185004 293734
rect 184404 258054 185004 293498
rect 184404 257818 184586 258054
rect 184822 257818 185004 258054
rect 184404 257734 185004 257818
rect 184404 257498 184586 257734
rect 184822 257498 185004 257734
rect 184404 222054 185004 257498
rect 184404 221818 184586 222054
rect 184822 221818 185004 222054
rect 184404 221734 185004 221818
rect 184404 221498 184586 221734
rect 184822 221498 185004 221734
rect 184404 186054 185004 221498
rect 184404 185818 184586 186054
rect 184822 185818 185004 186054
rect 184404 185734 185004 185818
rect 184404 185498 184586 185734
rect 184822 185498 185004 185734
rect 184404 150054 185004 185498
rect 184404 149818 184586 150054
rect 184822 149818 185004 150054
rect 184404 149734 185004 149818
rect 184404 149498 184586 149734
rect 184822 149498 185004 149734
rect 184404 114054 185004 149498
rect 184404 113818 184586 114054
rect 184822 113818 185004 114054
rect 184404 113734 185004 113818
rect 184404 113498 184586 113734
rect 184822 113498 185004 113734
rect 184404 78054 185004 113498
rect 184404 77818 184586 78054
rect 184822 77818 185004 78054
rect 184404 77734 185004 77818
rect 184404 77498 184586 77734
rect 184822 77498 185004 77734
rect 184404 42054 185004 77498
rect 184404 41818 184586 42054
rect 184822 41818 185004 42054
rect 184404 41734 185004 41818
rect 184404 41498 184586 41734
rect 184822 41498 185004 41734
rect 184404 6054 185004 41498
rect 184404 5818 184586 6054
rect 184822 5818 185004 6054
rect 184404 5734 185004 5818
rect 184404 5498 184586 5734
rect 184822 5498 185004 5734
rect 184404 -2186 185004 5498
rect 184404 -2422 184586 -2186
rect 184822 -2422 185004 -2186
rect 184404 -2506 185004 -2422
rect 184404 -2742 184586 -2506
rect 184822 -2742 185004 -2506
rect 184404 -3684 185004 -2742
rect 188004 693654 188604 707962
rect 188004 693418 188186 693654
rect 188422 693418 188604 693654
rect 188004 693334 188604 693418
rect 188004 693098 188186 693334
rect 188422 693098 188604 693334
rect 188004 657654 188604 693098
rect 188004 657418 188186 657654
rect 188422 657418 188604 657654
rect 188004 657334 188604 657418
rect 188004 657098 188186 657334
rect 188422 657098 188604 657334
rect 188004 621654 188604 657098
rect 188004 621418 188186 621654
rect 188422 621418 188604 621654
rect 188004 621334 188604 621418
rect 188004 621098 188186 621334
rect 188422 621098 188604 621334
rect 188004 585654 188604 621098
rect 188004 585418 188186 585654
rect 188422 585418 188604 585654
rect 188004 585334 188604 585418
rect 188004 585098 188186 585334
rect 188422 585098 188604 585334
rect 188004 549654 188604 585098
rect 188004 549418 188186 549654
rect 188422 549418 188604 549654
rect 188004 549334 188604 549418
rect 188004 549098 188186 549334
rect 188422 549098 188604 549334
rect 188004 513654 188604 549098
rect 188004 513418 188186 513654
rect 188422 513418 188604 513654
rect 188004 513334 188604 513418
rect 188004 513098 188186 513334
rect 188422 513098 188604 513334
rect 188004 477654 188604 513098
rect 188004 477418 188186 477654
rect 188422 477418 188604 477654
rect 188004 477334 188604 477418
rect 188004 477098 188186 477334
rect 188422 477098 188604 477334
rect 188004 441654 188604 477098
rect 188004 441418 188186 441654
rect 188422 441418 188604 441654
rect 188004 441334 188604 441418
rect 188004 441098 188186 441334
rect 188422 441098 188604 441334
rect 188004 405654 188604 441098
rect 188004 405418 188186 405654
rect 188422 405418 188604 405654
rect 188004 405334 188604 405418
rect 188004 405098 188186 405334
rect 188422 405098 188604 405334
rect 188004 369654 188604 405098
rect 188004 369418 188186 369654
rect 188422 369418 188604 369654
rect 188004 369334 188604 369418
rect 188004 369098 188186 369334
rect 188422 369098 188604 369334
rect 188004 333654 188604 369098
rect 188004 333418 188186 333654
rect 188422 333418 188604 333654
rect 188004 333334 188604 333418
rect 188004 333098 188186 333334
rect 188422 333098 188604 333334
rect 188004 297654 188604 333098
rect 188004 297418 188186 297654
rect 188422 297418 188604 297654
rect 188004 297334 188604 297418
rect 188004 297098 188186 297334
rect 188422 297098 188604 297334
rect 188004 261654 188604 297098
rect 188004 261418 188186 261654
rect 188422 261418 188604 261654
rect 188004 261334 188604 261418
rect 188004 261098 188186 261334
rect 188422 261098 188604 261334
rect 188004 225654 188604 261098
rect 188004 225418 188186 225654
rect 188422 225418 188604 225654
rect 188004 225334 188604 225418
rect 188004 225098 188186 225334
rect 188422 225098 188604 225334
rect 188004 189654 188604 225098
rect 188004 189418 188186 189654
rect 188422 189418 188604 189654
rect 188004 189334 188604 189418
rect 188004 189098 188186 189334
rect 188422 189098 188604 189334
rect 188004 153654 188604 189098
rect 188004 153418 188186 153654
rect 188422 153418 188604 153654
rect 188004 153334 188604 153418
rect 188004 153098 188186 153334
rect 188422 153098 188604 153334
rect 188004 117654 188604 153098
rect 188004 117418 188186 117654
rect 188422 117418 188604 117654
rect 188004 117334 188604 117418
rect 188004 117098 188186 117334
rect 188422 117098 188604 117334
rect 188004 81654 188604 117098
rect 188004 81418 188186 81654
rect 188422 81418 188604 81654
rect 188004 81334 188604 81418
rect 188004 81098 188186 81334
rect 188422 81098 188604 81334
rect 188004 45654 188604 81098
rect 188004 45418 188186 45654
rect 188422 45418 188604 45654
rect 188004 45334 188604 45418
rect 188004 45098 188186 45334
rect 188422 45098 188604 45334
rect 188004 9654 188604 45098
rect 188004 9418 188186 9654
rect 188422 9418 188604 9654
rect 188004 9334 188604 9418
rect 188004 9098 188186 9334
rect 188422 9098 188604 9334
rect 188004 -4026 188604 9098
rect 188004 -4262 188186 -4026
rect 188422 -4262 188604 -4026
rect 188004 -4346 188604 -4262
rect 188004 -4582 188186 -4346
rect 188422 -4582 188604 -4346
rect 188004 -5524 188604 -4582
rect 191604 697254 192204 709802
rect 209604 711278 210204 711300
rect 209604 711042 209786 711278
rect 210022 711042 210204 711278
rect 209604 710958 210204 711042
rect 209604 710722 209786 710958
rect 210022 710722 210204 710958
rect 206004 709438 206604 709460
rect 206004 709202 206186 709438
rect 206422 709202 206604 709438
rect 206004 709118 206604 709202
rect 206004 708882 206186 709118
rect 206422 708882 206604 709118
rect 202404 707598 203004 707620
rect 202404 707362 202586 707598
rect 202822 707362 203004 707598
rect 202404 707278 203004 707362
rect 202404 707042 202586 707278
rect 202822 707042 203004 707278
rect 191604 697018 191786 697254
rect 192022 697018 192204 697254
rect 191604 696934 192204 697018
rect 191604 696698 191786 696934
rect 192022 696698 192204 696934
rect 191604 661254 192204 696698
rect 191604 661018 191786 661254
rect 192022 661018 192204 661254
rect 191604 660934 192204 661018
rect 191604 660698 191786 660934
rect 192022 660698 192204 660934
rect 191604 625254 192204 660698
rect 191604 625018 191786 625254
rect 192022 625018 192204 625254
rect 191604 624934 192204 625018
rect 191604 624698 191786 624934
rect 192022 624698 192204 624934
rect 191604 589254 192204 624698
rect 191604 589018 191786 589254
rect 192022 589018 192204 589254
rect 191604 588934 192204 589018
rect 191604 588698 191786 588934
rect 192022 588698 192204 588934
rect 191604 553254 192204 588698
rect 191604 553018 191786 553254
rect 192022 553018 192204 553254
rect 191604 552934 192204 553018
rect 191604 552698 191786 552934
rect 192022 552698 192204 552934
rect 191604 517254 192204 552698
rect 198804 705758 199404 705780
rect 198804 705522 198986 705758
rect 199222 705522 199404 705758
rect 198804 705438 199404 705522
rect 198804 705202 198986 705438
rect 199222 705202 199404 705438
rect 198804 668454 199404 705202
rect 198804 668218 198986 668454
rect 199222 668218 199404 668454
rect 198804 668134 199404 668218
rect 198804 667898 198986 668134
rect 199222 667898 199404 668134
rect 198804 632454 199404 667898
rect 198804 632218 198986 632454
rect 199222 632218 199404 632454
rect 198804 632134 199404 632218
rect 198804 631898 198986 632134
rect 199222 631898 199404 632134
rect 198804 596454 199404 631898
rect 198804 596218 198986 596454
rect 199222 596218 199404 596454
rect 198804 596134 199404 596218
rect 198804 595898 198986 596134
rect 199222 595898 199404 596134
rect 198804 560454 199404 595898
rect 198804 560218 198986 560454
rect 199222 560218 199404 560454
rect 198804 560134 199404 560218
rect 198804 559898 198986 560134
rect 199222 559898 199404 560134
rect 198804 524454 199404 559898
rect 198804 524218 198986 524454
rect 199222 524218 199404 524454
rect 198804 524134 199404 524218
rect 198804 523898 198986 524134
rect 199222 523898 199404 524134
rect 193075 519348 193141 519349
rect 193075 519284 193076 519348
rect 193140 519284 193141 519348
rect 193075 519283 193141 519284
rect 195099 519348 195165 519349
rect 195099 519284 195100 519348
rect 195164 519284 195165 519348
rect 195099 519283 195165 519284
rect 198411 519348 198477 519349
rect 198411 519284 198412 519348
rect 198476 519284 198477 519348
rect 198411 519283 198477 519284
rect 193078 518125 193138 519283
rect 195102 518261 195162 519283
rect 198414 518397 198474 519283
rect 198411 518396 198477 518397
rect 198411 518332 198412 518396
rect 198476 518332 198477 518396
rect 198411 518331 198477 518332
rect 195099 518260 195165 518261
rect 195099 518196 195100 518260
rect 195164 518196 195165 518260
rect 195099 518195 195165 518196
rect 193075 518124 193141 518125
rect 193075 518060 193076 518124
rect 193140 518060 193141 518124
rect 193075 518059 193141 518060
rect 196019 517988 196085 517989
rect 196019 517924 196020 517988
rect 196084 517924 196085 517988
rect 196019 517923 196085 517924
rect 195835 517852 195901 517853
rect 195835 517788 195836 517852
rect 195900 517850 195901 517852
rect 196022 517850 196082 517923
rect 195900 517790 196082 517850
rect 195900 517788 195901 517790
rect 195835 517787 195901 517788
rect 191604 517018 191786 517254
rect 192022 517018 192204 517254
rect 191604 516934 192204 517018
rect 191604 516698 191786 516934
rect 192022 516698 192204 516934
rect 191604 481254 192204 516698
rect 191604 481018 191786 481254
rect 192022 481018 192204 481254
rect 191604 480934 192204 481018
rect 191604 480698 191786 480934
rect 192022 480698 192204 480934
rect 191604 445254 192204 480698
rect 191604 445018 191786 445254
rect 192022 445018 192204 445254
rect 191604 444934 192204 445018
rect 191604 444698 191786 444934
rect 192022 444698 192204 444934
rect 191604 409254 192204 444698
rect 191604 409018 191786 409254
rect 192022 409018 192204 409254
rect 191604 408934 192204 409018
rect 191604 408698 191786 408934
rect 192022 408698 192204 408934
rect 191604 373254 192204 408698
rect 191604 373018 191786 373254
rect 192022 373018 192204 373254
rect 191604 372934 192204 373018
rect 191604 372698 191786 372934
rect 192022 372698 192204 372934
rect 191604 337254 192204 372698
rect 191604 337018 191786 337254
rect 192022 337018 192204 337254
rect 191604 336934 192204 337018
rect 191604 336698 191786 336934
rect 192022 336698 192204 336934
rect 191604 301254 192204 336698
rect 191604 301018 191786 301254
rect 192022 301018 192204 301254
rect 191604 300934 192204 301018
rect 191604 300698 191786 300934
rect 192022 300698 192204 300934
rect 191604 265254 192204 300698
rect 191604 265018 191786 265254
rect 192022 265018 192204 265254
rect 191604 264934 192204 265018
rect 191604 264698 191786 264934
rect 192022 264698 192204 264934
rect 191604 229254 192204 264698
rect 191604 229018 191786 229254
rect 192022 229018 192204 229254
rect 191604 228934 192204 229018
rect 191604 228698 191786 228934
rect 192022 228698 192204 228934
rect 191604 193254 192204 228698
rect 191604 193018 191786 193254
rect 192022 193018 192204 193254
rect 191604 192934 192204 193018
rect 191604 192698 191786 192934
rect 192022 192698 192204 192934
rect 191604 157254 192204 192698
rect 191604 157018 191786 157254
rect 192022 157018 192204 157254
rect 191604 156934 192204 157018
rect 191604 156698 191786 156934
rect 192022 156698 192204 156934
rect 191604 121254 192204 156698
rect 198804 488454 199404 523898
rect 202404 672054 203004 707042
rect 202404 671818 202586 672054
rect 202822 671818 203004 672054
rect 202404 671734 203004 671818
rect 202404 671498 202586 671734
rect 202822 671498 203004 671734
rect 202404 636054 203004 671498
rect 202404 635818 202586 636054
rect 202822 635818 203004 636054
rect 202404 635734 203004 635818
rect 202404 635498 202586 635734
rect 202822 635498 203004 635734
rect 202404 600054 203004 635498
rect 202404 599818 202586 600054
rect 202822 599818 203004 600054
rect 202404 599734 203004 599818
rect 202404 599498 202586 599734
rect 202822 599498 203004 599734
rect 202404 564054 203004 599498
rect 202404 563818 202586 564054
rect 202822 563818 203004 564054
rect 202404 563734 203004 563818
rect 202404 563498 202586 563734
rect 202822 563498 203004 563734
rect 202404 528054 203004 563498
rect 202404 527818 202586 528054
rect 202822 527818 203004 528054
rect 202404 527734 203004 527818
rect 202404 527498 202586 527734
rect 202822 527498 203004 527734
rect 199883 519348 199949 519349
rect 199883 519284 199884 519348
rect 199948 519284 199949 519348
rect 199883 519283 199949 519284
rect 199886 518533 199946 519283
rect 199883 518532 199949 518533
rect 199883 518468 199884 518532
rect 199948 518468 199949 518532
rect 199883 518467 199949 518468
rect 198804 488218 198986 488454
rect 199222 488218 199404 488454
rect 198804 488134 199404 488218
rect 198804 487898 198986 488134
rect 199222 487898 199404 488134
rect 198804 452454 199404 487898
rect 198804 452218 198986 452454
rect 199222 452218 199404 452454
rect 198804 452134 199404 452218
rect 198804 451898 198986 452134
rect 199222 451898 199404 452134
rect 198804 416454 199404 451898
rect 198804 416218 198986 416454
rect 199222 416218 199404 416454
rect 198804 416134 199404 416218
rect 198804 415898 198986 416134
rect 199222 415898 199404 416134
rect 198804 380454 199404 415898
rect 198804 380218 198986 380454
rect 199222 380218 199404 380454
rect 198804 380134 199404 380218
rect 198804 379898 198986 380134
rect 199222 379898 199404 380134
rect 198804 344454 199404 379898
rect 198804 344218 198986 344454
rect 199222 344218 199404 344454
rect 198804 344134 199404 344218
rect 198804 343898 198986 344134
rect 199222 343898 199404 344134
rect 198804 308454 199404 343898
rect 198804 308218 198986 308454
rect 199222 308218 199404 308454
rect 198804 308134 199404 308218
rect 198804 307898 198986 308134
rect 199222 307898 199404 308134
rect 198804 272454 199404 307898
rect 198804 272218 198986 272454
rect 199222 272218 199404 272454
rect 198804 272134 199404 272218
rect 198804 271898 198986 272134
rect 199222 271898 199404 272134
rect 198804 236454 199404 271898
rect 198804 236218 198986 236454
rect 199222 236218 199404 236454
rect 198804 236134 199404 236218
rect 198804 235898 198986 236134
rect 199222 235898 199404 236134
rect 198804 200454 199404 235898
rect 198804 200218 198986 200454
rect 199222 200218 199404 200454
rect 198804 200134 199404 200218
rect 198804 199898 198986 200134
rect 199222 199898 199404 200134
rect 198804 164454 199404 199898
rect 198804 164218 198986 164454
rect 199222 164218 199404 164454
rect 198804 164134 199404 164218
rect 198804 163898 198986 164134
rect 199222 163898 199404 164134
rect 194915 143580 194981 143581
rect 194915 143516 194916 143580
rect 194980 143516 194981 143580
rect 194915 143515 194981 143516
rect 194918 142221 194978 143515
rect 194915 142220 194981 142221
rect 194915 142156 194916 142220
rect 194980 142156 194981 142220
rect 194915 142155 194981 142156
rect 191604 121018 191786 121254
rect 192022 121018 192204 121254
rect 191604 120934 192204 121018
rect 191604 120698 191786 120934
rect 192022 120698 192204 120934
rect 191604 85254 192204 120698
rect 191604 85018 191786 85254
rect 192022 85018 192204 85254
rect 191604 84934 192204 85018
rect 191604 84698 191786 84934
rect 192022 84698 192204 84934
rect 191604 49254 192204 84698
rect 198804 128454 199404 163898
rect 198804 128218 198986 128454
rect 199222 128218 199404 128454
rect 198804 128134 199404 128218
rect 198804 127898 198986 128134
rect 199222 127898 199404 128134
rect 198804 92454 199404 127898
rect 198804 92218 198986 92454
rect 199222 92218 199404 92454
rect 198804 92134 199404 92218
rect 198804 91898 198986 92134
rect 199222 91898 199404 92134
rect 195099 66196 195165 66197
rect 195099 66132 195100 66196
rect 195164 66132 195165 66196
rect 195099 66131 195165 66132
rect 195102 57901 195162 66131
rect 195099 57900 195165 57901
rect 195099 57836 195100 57900
rect 195164 57836 195165 57900
rect 195099 57835 195165 57836
rect 191604 49018 191786 49254
rect 192022 49018 192204 49254
rect 191604 48934 192204 49018
rect 191604 48698 191786 48934
rect 192022 48698 192204 48934
rect 191604 13254 192204 48698
rect 191604 13018 191786 13254
rect 192022 13018 192204 13254
rect 191604 12934 192204 13018
rect 191604 12698 191786 12934
rect 192022 12698 192204 12934
rect 173604 -7022 173786 -6786
rect 174022 -7022 174204 -6786
rect 173604 -7106 174204 -7022
rect 173604 -7342 173786 -7106
rect 174022 -7342 174204 -7106
rect 173604 -7364 174204 -7342
rect 191604 -5866 192204 12698
rect 198804 56454 199404 91898
rect 198804 56218 198986 56454
rect 199222 56218 199404 56454
rect 198804 56134 199404 56218
rect 198804 55898 198986 56134
rect 199222 55898 199404 56134
rect 198804 20454 199404 55898
rect 198804 20218 198986 20454
rect 199222 20218 199404 20454
rect 198804 20134 199404 20218
rect 198804 19898 198986 20134
rect 199222 19898 199404 20134
rect 198804 -1266 199404 19898
rect 198804 -1502 198986 -1266
rect 199222 -1502 199404 -1266
rect 198804 -1586 199404 -1502
rect 198804 -1822 198986 -1586
rect 199222 -1822 199404 -1586
rect 198804 -1844 199404 -1822
rect 202404 492054 203004 527498
rect 206004 675654 206604 708882
rect 206004 675418 206186 675654
rect 206422 675418 206604 675654
rect 206004 675334 206604 675418
rect 206004 675098 206186 675334
rect 206422 675098 206604 675334
rect 206004 639654 206604 675098
rect 206004 639418 206186 639654
rect 206422 639418 206604 639654
rect 206004 639334 206604 639418
rect 206004 639098 206186 639334
rect 206422 639098 206604 639334
rect 206004 603654 206604 639098
rect 206004 603418 206186 603654
rect 206422 603418 206604 603654
rect 206004 603334 206604 603418
rect 206004 603098 206186 603334
rect 206422 603098 206604 603334
rect 206004 567654 206604 603098
rect 206004 567418 206186 567654
rect 206422 567418 206604 567654
rect 206004 567334 206604 567418
rect 206004 567098 206186 567334
rect 206422 567098 206604 567334
rect 206004 531654 206604 567098
rect 206004 531418 206186 531654
rect 206422 531418 206604 531654
rect 206004 531334 206604 531418
rect 206004 531098 206186 531334
rect 206422 531098 206604 531334
rect 205219 519348 205285 519349
rect 205219 519284 205220 519348
rect 205284 519284 205285 519348
rect 205219 519283 205285 519284
rect 205222 517853 205282 519283
rect 205219 517852 205285 517853
rect 205219 517788 205220 517852
rect 205284 517788 205285 517852
rect 205219 517787 205285 517788
rect 202404 491818 202586 492054
rect 202822 491818 203004 492054
rect 202404 491734 203004 491818
rect 202404 491498 202586 491734
rect 202822 491498 203004 491734
rect 202404 456054 203004 491498
rect 202404 455818 202586 456054
rect 202822 455818 203004 456054
rect 202404 455734 203004 455818
rect 202404 455498 202586 455734
rect 202822 455498 203004 455734
rect 202404 420054 203004 455498
rect 202404 419818 202586 420054
rect 202822 419818 203004 420054
rect 202404 419734 203004 419818
rect 202404 419498 202586 419734
rect 202822 419498 203004 419734
rect 202404 384054 203004 419498
rect 202404 383818 202586 384054
rect 202822 383818 203004 384054
rect 202404 383734 203004 383818
rect 202404 383498 202586 383734
rect 202822 383498 203004 383734
rect 202404 348054 203004 383498
rect 202404 347818 202586 348054
rect 202822 347818 203004 348054
rect 202404 347734 203004 347818
rect 202404 347498 202586 347734
rect 202822 347498 203004 347734
rect 202404 312054 203004 347498
rect 202404 311818 202586 312054
rect 202822 311818 203004 312054
rect 202404 311734 203004 311818
rect 202404 311498 202586 311734
rect 202822 311498 203004 311734
rect 202404 276054 203004 311498
rect 202404 275818 202586 276054
rect 202822 275818 203004 276054
rect 202404 275734 203004 275818
rect 202404 275498 202586 275734
rect 202822 275498 203004 275734
rect 202404 240054 203004 275498
rect 202404 239818 202586 240054
rect 202822 239818 203004 240054
rect 202404 239734 203004 239818
rect 202404 239498 202586 239734
rect 202822 239498 203004 239734
rect 202404 204054 203004 239498
rect 202404 203818 202586 204054
rect 202822 203818 203004 204054
rect 202404 203734 203004 203818
rect 202404 203498 202586 203734
rect 202822 203498 203004 203734
rect 202404 168054 203004 203498
rect 202404 167818 202586 168054
rect 202822 167818 203004 168054
rect 202404 167734 203004 167818
rect 202404 167498 202586 167734
rect 202822 167498 203004 167734
rect 202404 132054 203004 167498
rect 202404 131818 202586 132054
rect 202822 131818 203004 132054
rect 202404 131734 203004 131818
rect 202404 131498 202586 131734
rect 202822 131498 203004 131734
rect 202404 96054 203004 131498
rect 202404 95818 202586 96054
rect 202822 95818 203004 96054
rect 202404 95734 203004 95818
rect 202404 95498 202586 95734
rect 202822 95498 203004 95734
rect 202404 60054 203004 95498
rect 202404 59818 202586 60054
rect 202822 59818 203004 60054
rect 202404 59734 203004 59818
rect 202404 59498 202586 59734
rect 202822 59498 203004 59734
rect 202404 24054 203004 59498
rect 202404 23818 202586 24054
rect 202822 23818 203004 24054
rect 202404 23734 203004 23818
rect 202404 23498 202586 23734
rect 202822 23498 203004 23734
rect 202404 -3106 203004 23498
rect 202404 -3342 202586 -3106
rect 202822 -3342 203004 -3106
rect 202404 -3426 203004 -3342
rect 202404 -3662 202586 -3426
rect 202822 -3662 203004 -3426
rect 202404 -3684 203004 -3662
rect 206004 495654 206604 531098
rect 206004 495418 206186 495654
rect 206422 495418 206604 495654
rect 206004 495334 206604 495418
rect 206004 495098 206186 495334
rect 206422 495098 206604 495334
rect 206004 459654 206604 495098
rect 206004 459418 206186 459654
rect 206422 459418 206604 459654
rect 206004 459334 206604 459418
rect 206004 459098 206186 459334
rect 206422 459098 206604 459334
rect 206004 423654 206604 459098
rect 206004 423418 206186 423654
rect 206422 423418 206604 423654
rect 206004 423334 206604 423418
rect 206004 423098 206186 423334
rect 206422 423098 206604 423334
rect 206004 387654 206604 423098
rect 206004 387418 206186 387654
rect 206422 387418 206604 387654
rect 206004 387334 206604 387418
rect 206004 387098 206186 387334
rect 206422 387098 206604 387334
rect 206004 351654 206604 387098
rect 206004 351418 206186 351654
rect 206422 351418 206604 351654
rect 206004 351334 206604 351418
rect 206004 351098 206186 351334
rect 206422 351098 206604 351334
rect 206004 315654 206604 351098
rect 206004 315418 206186 315654
rect 206422 315418 206604 315654
rect 206004 315334 206604 315418
rect 206004 315098 206186 315334
rect 206422 315098 206604 315334
rect 206004 279654 206604 315098
rect 206004 279418 206186 279654
rect 206422 279418 206604 279654
rect 206004 279334 206604 279418
rect 206004 279098 206186 279334
rect 206422 279098 206604 279334
rect 206004 243654 206604 279098
rect 206004 243418 206186 243654
rect 206422 243418 206604 243654
rect 206004 243334 206604 243418
rect 206004 243098 206186 243334
rect 206422 243098 206604 243334
rect 206004 207654 206604 243098
rect 206004 207418 206186 207654
rect 206422 207418 206604 207654
rect 206004 207334 206604 207418
rect 206004 207098 206186 207334
rect 206422 207098 206604 207334
rect 206004 171654 206604 207098
rect 206004 171418 206186 171654
rect 206422 171418 206604 171654
rect 206004 171334 206604 171418
rect 206004 171098 206186 171334
rect 206422 171098 206604 171334
rect 206004 135654 206604 171098
rect 206004 135418 206186 135654
rect 206422 135418 206604 135654
rect 206004 135334 206604 135418
rect 206004 135098 206186 135334
rect 206422 135098 206604 135334
rect 206004 99654 206604 135098
rect 206004 99418 206186 99654
rect 206422 99418 206604 99654
rect 206004 99334 206604 99418
rect 206004 99098 206186 99334
rect 206422 99098 206604 99334
rect 206004 63654 206604 99098
rect 206004 63418 206186 63654
rect 206422 63418 206604 63654
rect 206004 63334 206604 63418
rect 206004 63098 206186 63334
rect 206422 63098 206604 63334
rect 206004 27654 206604 63098
rect 206004 27418 206186 27654
rect 206422 27418 206604 27654
rect 206004 27334 206604 27418
rect 206004 27098 206186 27334
rect 206422 27098 206604 27334
rect 206004 -4946 206604 27098
rect 206004 -5182 206186 -4946
rect 206422 -5182 206604 -4946
rect 206004 -5266 206604 -5182
rect 206004 -5502 206186 -5266
rect 206422 -5502 206604 -5266
rect 206004 -5524 206604 -5502
rect 209604 679254 210204 710722
rect 227604 710358 228204 711300
rect 227604 710122 227786 710358
rect 228022 710122 228204 710358
rect 227604 710038 228204 710122
rect 227604 709802 227786 710038
rect 228022 709802 228204 710038
rect 224004 708518 224604 709460
rect 224004 708282 224186 708518
rect 224422 708282 224604 708518
rect 224004 708198 224604 708282
rect 224004 707962 224186 708198
rect 224422 707962 224604 708198
rect 220404 706678 221004 707620
rect 220404 706442 220586 706678
rect 220822 706442 221004 706678
rect 220404 706358 221004 706442
rect 220404 706122 220586 706358
rect 220822 706122 221004 706358
rect 209604 679018 209786 679254
rect 210022 679018 210204 679254
rect 209604 678934 210204 679018
rect 209604 678698 209786 678934
rect 210022 678698 210204 678934
rect 209604 643254 210204 678698
rect 209604 643018 209786 643254
rect 210022 643018 210204 643254
rect 209604 642934 210204 643018
rect 209604 642698 209786 642934
rect 210022 642698 210204 642934
rect 209604 607254 210204 642698
rect 209604 607018 209786 607254
rect 210022 607018 210204 607254
rect 209604 606934 210204 607018
rect 209604 606698 209786 606934
rect 210022 606698 210204 606934
rect 209604 571254 210204 606698
rect 209604 571018 209786 571254
rect 210022 571018 210204 571254
rect 209604 570934 210204 571018
rect 209604 570698 209786 570934
rect 210022 570698 210204 570934
rect 209604 535254 210204 570698
rect 209604 535018 209786 535254
rect 210022 535018 210204 535254
rect 209604 534934 210204 535018
rect 209604 534698 209786 534934
rect 210022 534698 210204 534934
rect 209604 499254 210204 534698
rect 216804 704838 217404 705780
rect 216804 704602 216986 704838
rect 217222 704602 217404 704838
rect 216804 704518 217404 704602
rect 216804 704282 216986 704518
rect 217222 704282 217404 704518
rect 216804 686454 217404 704282
rect 216804 686218 216986 686454
rect 217222 686218 217404 686454
rect 216804 686134 217404 686218
rect 216804 685898 216986 686134
rect 217222 685898 217404 686134
rect 216804 650454 217404 685898
rect 216804 650218 216986 650454
rect 217222 650218 217404 650454
rect 216804 650134 217404 650218
rect 216804 649898 216986 650134
rect 217222 649898 217404 650134
rect 216804 614454 217404 649898
rect 216804 614218 216986 614454
rect 217222 614218 217404 614454
rect 216804 614134 217404 614218
rect 216804 613898 216986 614134
rect 217222 613898 217404 614134
rect 216804 578454 217404 613898
rect 216804 578218 216986 578454
rect 217222 578218 217404 578454
rect 216804 578134 217404 578218
rect 216804 577898 216986 578134
rect 217222 577898 217404 578134
rect 216804 542454 217404 577898
rect 216804 542218 216986 542454
rect 217222 542218 217404 542454
rect 216804 542134 217404 542218
rect 216804 541898 216986 542134
rect 217222 541898 217404 542134
rect 210371 519348 210437 519349
rect 210371 519284 210372 519348
rect 210436 519284 210437 519348
rect 210371 519283 210437 519284
rect 210374 518669 210434 519283
rect 210371 518668 210437 518669
rect 210371 518604 210372 518668
rect 210436 518604 210437 518668
rect 210371 518603 210437 518604
rect 210371 517988 210437 517989
rect 210371 517938 210372 517988
rect 210436 517938 210437 517988
rect 209604 499018 209786 499254
rect 210022 499018 210204 499254
rect 209604 498934 210204 499018
rect 209604 498698 209786 498934
rect 210022 498698 210204 498934
rect 209604 463254 210204 498698
rect 209604 463018 209786 463254
rect 210022 463018 210204 463254
rect 209604 462934 210204 463018
rect 209604 462698 209786 462934
rect 210022 462698 210204 462934
rect 209604 427254 210204 462698
rect 209604 427018 209786 427254
rect 210022 427018 210204 427254
rect 209604 426934 210204 427018
rect 209604 426698 209786 426934
rect 210022 426698 210204 426934
rect 209604 391254 210204 426698
rect 209604 391018 209786 391254
rect 210022 391018 210204 391254
rect 209604 390934 210204 391018
rect 209604 390698 209786 390934
rect 210022 390698 210204 390934
rect 209604 355254 210204 390698
rect 209604 355018 209786 355254
rect 210022 355018 210204 355254
rect 209604 354934 210204 355018
rect 209604 354698 209786 354934
rect 210022 354698 210204 354934
rect 209604 319254 210204 354698
rect 209604 319018 209786 319254
rect 210022 319018 210204 319254
rect 209604 318934 210204 319018
rect 209604 318698 209786 318934
rect 210022 318698 210204 318934
rect 209604 283254 210204 318698
rect 209604 283018 209786 283254
rect 210022 283018 210204 283254
rect 209604 282934 210204 283018
rect 209604 282698 209786 282934
rect 210022 282698 210204 282934
rect 209604 247254 210204 282698
rect 209604 247018 209786 247254
rect 210022 247018 210204 247254
rect 209604 246934 210204 247018
rect 209604 246698 209786 246934
rect 210022 246698 210204 246934
rect 209604 211254 210204 246698
rect 209604 211018 209786 211254
rect 210022 211018 210204 211254
rect 209604 210934 210204 211018
rect 209604 210698 209786 210934
rect 210022 210698 210204 210934
rect 209604 175254 210204 210698
rect 209604 175018 209786 175254
rect 210022 175018 210204 175254
rect 209604 174934 210204 175018
rect 209604 174698 209786 174934
rect 210022 174698 210204 174934
rect 209604 139254 210204 174698
rect 209604 139018 209786 139254
rect 210022 139018 210204 139254
rect 209604 138934 210204 139018
rect 209604 138698 209786 138934
rect 210022 138698 210204 138934
rect 209604 103254 210204 138698
rect 209604 103018 209786 103254
rect 210022 103018 210204 103254
rect 209604 102934 210204 103018
rect 209604 102698 209786 102934
rect 210022 102698 210204 102934
rect 209604 67254 210204 102698
rect 209604 67018 209786 67254
rect 210022 67018 210204 67254
rect 209604 66934 210204 67018
rect 209604 66698 209786 66934
rect 210022 66698 210204 66934
rect 209604 31254 210204 66698
rect 209604 31018 209786 31254
rect 210022 31018 210204 31254
rect 209604 30934 210204 31018
rect 209604 30698 209786 30934
rect 210022 30698 210204 30934
rect 191604 -6102 191786 -5866
rect 192022 -6102 192204 -5866
rect 191604 -6186 192204 -6102
rect 191604 -6422 191786 -6186
rect 192022 -6422 192204 -6186
rect 191604 -7364 192204 -6422
rect 209604 -6786 210204 30698
rect 216804 506454 217404 541898
rect 220404 690054 221004 706122
rect 220404 689818 220586 690054
rect 220822 689818 221004 690054
rect 220404 689734 221004 689818
rect 220404 689498 220586 689734
rect 220822 689498 221004 689734
rect 220404 654054 221004 689498
rect 220404 653818 220586 654054
rect 220822 653818 221004 654054
rect 220404 653734 221004 653818
rect 220404 653498 220586 653734
rect 220822 653498 221004 653734
rect 220404 618054 221004 653498
rect 220404 617818 220586 618054
rect 220822 617818 221004 618054
rect 220404 617734 221004 617818
rect 220404 617498 220586 617734
rect 220822 617498 221004 617734
rect 220404 582054 221004 617498
rect 220404 581818 220586 582054
rect 220822 581818 221004 582054
rect 220404 581734 221004 581818
rect 220404 581498 220586 581734
rect 220822 581498 221004 581734
rect 220404 546054 221004 581498
rect 220404 545818 220586 546054
rect 220822 545818 221004 546054
rect 220404 545734 221004 545818
rect 220404 545498 220586 545734
rect 220822 545498 221004 545734
rect 219203 517988 219269 517989
rect 219203 517938 219204 517988
rect 219268 517938 219269 517988
rect 216804 506218 216986 506454
rect 217222 506218 217404 506454
rect 216804 506134 217404 506218
rect 216804 505898 216986 506134
rect 217222 505898 217404 506134
rect 216804 470454 217404 505898
rect 216804 470218 216986 470454
rect 217222 470218 217404 470454
rect 216804 470134 217404 470218
rect 216804 469898 216986 470134
rect 217222 469898 217404 470134
rect 216804 434454 217404 469898
rect 216804 434218 216986 434454
rect 217222 434218 217404 434454
rect 216804 434134 217404 434218
rect 216804 433898 216986 434134
rect 217222 433898 217404 434134
rect 216804 398454 217404 433898
rect 216804 398218 216986 398454
rect 217222 398218 217404 398454
rect 216804 398134 217404 398218
rect 216804 397898 216986 398134
rect 217222 397898 217404 398134
rect 216804 362454 217404 397898
rect 216804 362218 216986 362454
rect 217222 362218 217404 362454
rect 216804 362134 217404 362218
rect 216804 361898 216986 362134
rect 217222 361898 217404 362134
rect 216804 326454 217404 361898
rect 216804 326218 216986 326454
rect 217222 326218 217404 326454
rect 216804 326134 217404 326218
rect 216804 325898 216986 326134
rect 217222 325898 217404 326134
rect 216804 290454 217404 325898
rect 216804 290218 216986 290454
rect 217222 290218 217404 290454
rect 216804 290134 217404 290218
rect 216804 289898 216986 290134
rect 217222 289898 217404 290134
rect 216804 254454 217404 289898
rect 216804 254218 216986 254454
rect 217222 254218 217404 254454
rect 216804 254134 217404 254218
rect 216804 253898 216986 254134
rect 217222 253898 217404 254134
rect 216804 218454 217404 253898
rect 216804 218218 216986 218454
rect 217222 218218 217404 218454
rect 216804 218134 217404 218218
rect 216804 217898 216986 218134
rect 217222 217898 217404 218134
rect 216804 182454 217404 217898
rect 216804 182218 216986 182454
rect 217222 182218 217404 182454
rect 216804 182134 217404 182218
rect 216804 181898 216986 182134
rect 217222 181898 217404 182134
rect 216804 146454 217404 181898
rect 216804 146218 216986 146454
rect 217222 146218 217404 146454
rect 216804 146134 217404 146218
rect 216804 145898 216986 146134
rect 217222 145898 217404 146134
rect 216804 110454 217404 145898
rect 216804 110218 216986 110454
rect 217222 110218 217404 110454
rect 216804 110134 217404 110218
rect 216804 109898 216986 110134
rect 217222 109898 217404 110134
rect 216804 74454 217404 109898
rect 216804 74218 216986 74454
rect 217222 74218 217404 74454
rect 216804 74134 217404 74218
rect 216804 73898 216986 74134
rect 217222 73898 217404 74134
rect 216804 38454 217404 73898
rect 216804 38218 216986 38454
rect 217222 38218 217404 38454
rect 216804 38134 217404 38218
rect 216804 37898 216986 38134
rect 217222 37898 217404 38134
rect 216804 2454 217404 37898
rect 216804 2218 216986 2454
rect 217222 2218 217404 2454
rect 216804 2134 217404 2218
rect 216804 1898 216986 2134
rect 217222 1898 217404 2134
rect 216804 -346 217404 1898
rect 216804 -582 216986 -346
rect 217222 -582 217404 -346
rect 216804 -666 217404 -582
rect 216804 -902 216986 -666
rect 217222 -902 217404 -666
rect 216804 -1844 217404 -902
rect 220404 510054 221004 545498
rect 220404 509818 220586 510054
rect 220822 509818 221004 510054
rect 220404 509734 221004 509818
rect 220404 509498 220586 509734
rect 220822 509498 221004 509734
rect 220404 474054 221004 509498
rect 220404 473818 220586 474054
rect 220822 473818 221004 474054
rect 220404 473734 221004 473818
rect 220404 473498 220586 473734
rect 220822 473498 221004 473734
rect 220404 438054 221004 473498
rect 220404 437818 220586 438054
rect 220822 437818 221004 438054
rect 220404 437734 221004 437818
rect 220404 437498 220586 437734
rect 220822 437498 221004 437734
rect 220404 402054 221004 437498
rect 220404 401818 220586 402054
rect 220822 401818 221004 402054
rect 220404 401734 221004 401818
rect 220404 401498 220586 401734
rect 220822 401498 221004 401734
rect 220404 366054 221004 401498
rect 220404 365818 220586 366054
rect 220822 365818 221004 366054
rect 220404 365734 221004 365818
rect 220404 365498 220586 365734
rect 220822 365498 221004 365734
rect 220404 330054 221004 365498
rect 220404 329818 220586 330054
rect 220822 329818 221004 330054
rect 220404 329734 221004 329818
rect 220404 329498 220586 329734
rect 220822 329498 221004 329734
rect 220404 294054 221004 329498
rect 220404 293818 220586 294054
rect 220822 293818 221004 294054
rect 220404 293734 221004 293818
rect 220404 293498 220586 293734
rect 220822 293498 221004 293734
rect 220404 258054 221004 293498
rect 220404 257818 220586 258054
rect 220822 257818 221004 258054
rect 220404 257734 221004 257818
rect 220404 257498 220586 257734
rect 220822 257498 221004 257734
rect 220404 222054 221004 257498
rect 220404 221818 220586 222054
rect 220822 221818 221004 222054
rect 220404 221734 221004 221818
rect 220404 221498 220586 221734
rect 220822 221498 221004 221734
rect 220404 186054 221004 221498
rect 220404 185818 220586 186054
rect 220822 185818 221004 186054
rect 220404 185734 221004 185818
rect 220404 185498 220586 185734
rect 220822 185498 221004 185734
rect 220404 150054 221004 185498
rect 220404 149818 220586 150054
rect 220822 149818 221004 150054
rect 220404 149734 221004 149818
rect 220404 149498 220586 149734
rect 220822 149498 221004 149734
rect 220404 114054 221004 149498
rect 220404 113818 220586 114054
rect 220822 113818 221004 114054
rect 220404 113734 221004 113818
rect 220404 113498 220586 113734
rect 220822 113498 221004 113734
rect 220404 78054 221004 113498
rect 220404 77818 220586 78054
rect 220822 77818 221004 78054
rect 220404 77734 221004 77818
rect 220404 77498 220586 77734
rect 220822 77498 221004 77734
rect 220404 42054 221004 77498
rect 220404 41818 220586 42054
rect 220822 41818 221004 42054
rect 220404 41734 221004 41818
rect 220404 41498 220586 41734
rect 220822 41498 221004 41734
rect 220404 6054 221004 41498
rect 220404 5818 220586 6054
rect 220822 5818 221004 6054
rect 220404 5734 221004 5818
rect 220404 5498 220586 5734
rect 220822 5498 221004 5734
rect 220404 -2186 221004 5498
rect 220404 -2422 220586 -2186
rect 220822 -2422 221004 -2186
rect 220404 -2506 221004 -2422
rect 220404 -2742 220586 -2506
rect 220822 -2742 221004 -2506
rect 220404 -3684 221004 -2742
rect 224004 693654 224604 707962
rect 224004 693418 224186 693654
rect 224422 693418 224604 693654
rect 224004 693334 224604 693418
rect 224004 693098 224186 693334
rect 224422 693098 224604 693334
rect 224004 657654 224604 693098
rect 224004 657418 224186 657654
rect 224422 657418 224604 657654
rect 224004 657334 224604 657418
rect 224004 657098 224186 657334
rect 224422 657098 224604 657334
rect 224004 621654 224604 657098
rect 224004 621418 224186 621654
rect 224422 621418 224604 621654
rect 224004 621334 224604 621418
rect 224004 621098 224186 621334
rect 224422 621098 224604 621334
rect 224004 585654 224604 621098
rect 224004 585418 224186 585654
rect 224422 585418 224604 585654
rect 224004 585334 224604 585418
rect 224004 585098 224186 585334
rect 224422 585098 224604 585334
rect 224004 549654 224604 585098
rect 224004 549418 224186 549654
rect 224422 549418 224604 549654
rect 224004 549334 224604 549418
rect 224004 549098 224186 549334
rect 224422 549098 224604 549334
rect 224004 513654 224604 549098
rect 224004 513418 224186 513654
rect 224422 513418 224604 513654
rect 224004 513334 224604 513418
rect 224004 513098 224186 513334
rect 224422 513098 224604 513334
rect 224004 477654 224604 513098
rect 224004 477418 224186 477654
rect 224422 477418 224604 477654
rect 224004 477334 224604 477418
rect 224004 477098 224186 477334
rect 224422 477098 224604 477334
rect 224004 441654 224604 477098
rect 224004 441418 224186 441654
rect 224422 441418 224604 441654
rect 224004 441334 224604 441418
rect 224004 441098 224186 441334
rect 224422 441098 224604 441334
rect 224004 405654 224604 441098
rect 224004 405418 224186 405654
rect 224422 405418 224604 405654
rect 224004 405334 224604 405418
rect 224004 405098 224186 405334
rect 224422 405098 224604 405334
rect 224004 369654 224604 405098
rect 224004 369418 224186 369654
rect 224422 369418 224604 369654
rect 224004 369334 224604 369418
rect 224004 369098 224186 369334
rect 224422 369098 224604 369334
rect 224004 333654 224604 369098
rect 224004 333418 224186 333654
rect 224422 333418 224604 333654
rect 224004 333334 224604 333418
rect 224004 333098 224186 333334
rect 224422 333098 224604 333334
rect 224004 297654 224604 333098
rect 224004 297418 224186 297654
rect 224422 297418 224604 297654
rect 224004 297334 224604 297418
rect 224004 297098 224186 297334
rect 224422 297098 224604 297334
rect 224004 261654 224604 297098
rect 224004 261418 224186 261654
rect 224422 261418 224604 261654
rect 224004 261334 224604 261418
rect 224004 261098 224186 261334
rect 224422 261098 224604 261334
rect 224004 225654 224604 261098
rect 224004 225418 224186 225654
rect 224422 225418 224604 225654
rect 224004 225334 224604 225418
rect 224004 225098 224186 225334
rect 224422 225098 224604 225334
rect 224004 189654 224604 225098
rect 224004 189418 224186 189654
rect 224422 189418 224604 189654
rect 224004 189334 224604 189418
rect 224004 189098 224186 189334
rect 224422 189098 224604 189334
rect 224004 153654 224604 189098
rect 224004 153418 224186 153654
rect 224422 153418 224604 153654
rect 224004 153334 224604 153418
rect 224004 153098 224186 153334
rect 224422 153098 224604 153334
rect 224004 117654 224604 153098
rect 224004 117418 224186 117654
rect 224422 117418 224604 117654
rect 224004 117334 224604 117418
rect 224004 117098 224186 117334
rect 224422 117098 224604 117334
rect 224004 81654 224604 117098
rect 224004 81418 224186 81654
rect 224422 81418 224604 81654
rect 224004 81334 224604 81418
rect 224004 81098 224186 81334
rect 224422 81098 224604 81334
rect 224004 45654 224604 81098
rect 224004 45418 224186 45654
rect 224422 45418 224604 45654
rect 224004 45334 224604 45418
rect 224004 45098 224186 45334
rect 224422 45098 224604 45334
rect 224004 9654 224604 45098
rect 224004 9418 224186 9654
rect 224422 9418 224604 9654
rect 224004 9334 224604 9418
rect 224004 9098 224186 9334
rect 224422 9098 224604 9334
rect 224004 -4026 224604 9098
rect 224004 -4262 224186 -4026
rect 224422 -4262 224604 -4026
rect 224004 -4346 224604 -4262
rect 224004 -4582 224186 -4346
rect 224422 -4582 224604 -4346
rect 224004 -5524 224604 -4582
rect 227604 697254 228204 709802
rect 245604 711278 246204 711300
rect 245604 711042 245786 711278
rect 246022 711042 246204 711278
rect 245604 710958 246204 711042
rect 245604 710722 245786 710958
rect 246022 710722 246204 710958
rect 242004 709438 242604 709460
rect 242004 709202 242186 709438
rect 242422 709202 242604 709438
rect 242004 709118 242604 709202
rect 242004 708882 242186 709118
rect 242422 708882 242604 709118
rect 238404 707598 239004 707620
rect 238404 707362 238586 707598
rect 238822 707362 239004 707598
rect 238404 707278 239004 707362
rect 238404 707042 238586 707278
rect 238822 707042 239004 707278
rect 227604 697018 227786 697254
rect 228022 697018 228204 697254
rect 227604 696934 228204 697018
rect 227604 696698 227786 696934
rect 228022 696698 228204 696934
rect 227604 661254 228204 696698
rect 227604 661018 227786 661254
rect 228022 661018 228204 661254
rect 227604 660934 228204 661018
rect 227604 660698 227786 660934
rect 228022 660698 228204 660934
rect 227604 625254 228204 660698
rect 227604 625018 227786 625254
rect 228022 625018 228204 625254
rect 227604 624934 228204 625018
rect 227604 624698 227786 624934
rect 228022 624698 228204 624934
rect 227604 589254 228204 624698
rect 227604 589018 227786 589254
rect 228022 589018 228204 589254
rect 227604 588934 228204 589018
rect 227604 588698 227786 588934
rect 228022 588698 228204 588934
rect 227604 553254 228204 588698
rect 227604 553018 227786 553254
rect 228022 553018 228204 553254
rect 227604 552934 228204 553018
rect 227604 552698 227786 552934
rect 228022 552698 228204 552934
rect 227604 517254 228204 552698
rect 234804 705758 235404 705780
rect 234804 705522 234986 705758
rect 235222 705522 235404 705758
rect 234804 705438 235404 705522
rect 234804 705202 234986 705438
rect 235222 705202 235404 705438
rect 234804 668454 235404 705202
rect 234804 668218 234986 668454
rect 235222 668218 235404 668454
rect 234804 668134 235404 668218
rect 234804 667898 234986 668134
rect 235222 667898 235404 668134
rect 234804 632454 235404 667898
rect 234804 632218 234986 632454
rect 235222 632218 235404 632454
rect 234804 632134 235404 632218
rect 234804 631898 234986 632134
rect 235222 631898 235404 632134
rect 234804 596454 235404 631898
rect 234804 596218 234986 596454
rect 235222 596218 235404 596454
rect 234804 596134 235404 596218
rect 234804 595898 234986 596134
rect 235222 595898 235404 596134
rect 234804 560454 235404 595898
rect 234804 560218 234986 560454
rect 235222 560218 235404 560454
rect 234804 560134 235404 560218
rect 234804 559898 234986 560134
rect 235222 559898 235404 560134
rect 234804 524454 235404 559898
rect 234804 524218 234986 524454
rect 235222 524218 235404 524454
rect 234804 524134 235404 524218
rect 234804 523898 234986 524134
rect 235222 523898 235404 524134
rect 234291 519348 234357 519349
rect 234291 519284 234292 519348
rect 234356 519284 234357 519348
rect 234291 519283 234357 519284
rect 234294 518397 234354 519283
rect 234475 519212 234541 519213
rect 234475 519148 234476 519212
rect 234540 519148 234541 519212
rect 234475 519147 234541 519148
rect 234478 518669 234538 519147
rect 234475 518668 234541 518669
rect 234475 518604 234476 518668
rect 234540 518604 234541 518668
rect 234475 518603 234541 518604
rect 234291 518396 234357 518397
rect 234291 518332 234292 518396
rect 234356 518332 234357 518396
rect 234291 518331 234357 518332
rect 234659 518396 234725 518397
rect 234659 518332 234660 518396
rect 234724 518332 234725 518396
rect 234659 518331 234725 518332
rect 234662 518125 234722 518331
rect 234659 518124 234725 518125
rect 234659 518060 234660 518124
rect 234724 518060 234725 518124
rect 234659 518059 234725 518060
rect 234475 517988 234541 517989
rect 234475 517938 234476 517988
rect 234540 517938 234541 517988
rect 227604 517018 227786 517254
rect 228022 517018 228204 517254
rect 227604 516934 228204 517018
rect 227604 516698 227786 516934
rect 228022 516698 228204 516934
rect 227604 481254 228204 516698
rect 227604 481018 227786 481254
rect 228022 481018 228204 481254
rect 227604 480934 228204 481018
rect 227604 480698 227786 480934
rect 228022 480698 228204 480934
rect 227604 445254 228204 480698
rect 227604 445018 227786 445254
rect 228022 445018 228204 445254
rect 227604 444934 228204 445018
rect 227604 444698 227786 444934
rect 228022 444698 228204 444934
rect 227604 409254 228204 444698
rect 227604 409018 227786 409254
rect 228022 409018 228204 409254
rect 227604 408934 228204 409018
rect 227604 408698 227786 408934
rect 228022 408698 228204 408934
rect 227604 373254 228204 408698
rect 227604 373018 227786 373254
rect 228022 373018 228204 373254
rect 227604 372934 228204 373018
rect 227604 372698 227786 372934
rect 228022 372698 228204 372934
rect 227604 337254 228204 372698
rect 227604 337018 227786 337254
rect 228022 337018 228204 337254
rect 227604 336934 228204 337018
rect 227604 336698 227786 336934
rect 228022 336698 228204 336934
rect 227604 301254 228204 336698
rect 227604 301018 227786 301254
rect 228022 301018 228204 301254
rect 227604 300934 228204 301018
rect 227604 300698 227786 300934
rect 228022 300698 228204 300934
rect 227604 265254 228204 300698
rect 227604 265018 227786 265254
rect 228022 265018 228204 265254
rect 227604 264934 228204 265018
rect 227604 264698 227786 264934
rect 228022 264698 228204 264934
rect 227604 229254 228204 264698
rect 227604 229018 227786 229254
rect 228022 229018 228204 229254
rect 227604 228934 228204 229018
rect 227604 228698 227786 228934
rect 228022 228698 228204 228934
rect 227604 193254 228204 228698
rect 227604 193018 227786 193254
rect 228022 193018 228204 193254
rect 227604 192934 228204 193018
rect 227604 192698 227786 192934
rect 228022 192698 228204 192934
rect 227604 157254 228204 192698
rect 227604 157018 227786 157254
rect 228022 157018 228204 157254
rect 227604 156934 228204 157018
rect 227604 156698 227786 156934
rect 228022 156698 228204 156934
rect 227604 121254 228204 156698
rect 227604 121018 227786 121254
rect 228022 121018 228204 121254
rect 227604 120934 228204 121018
rect 227604 120698 227786 120934
rect 228022 120698 228204 120934
rect 227604 85254 228204 120698
rect 227604 85018 227786 85254
rect 228022 85018 228204 85254
rect 227604 84934 228204 85018
rect 227604 84698 227786 84934
rect 228022 84698 228204 84934
rect 227604 49254 228204 84698
rect 227604 49018 227786 49254
rect 228022 49018 228204 49254
rect 227604 48934 228204 49018
rect 227604 48698 227786 48934
rect 228022 48698 228204 48934
rect 227604 13254 228204 48698
rect 227604 13018 227786 13254
rect 228022 13018 228204 13254
rect 227604 12934 228204 13018
rect 227604 12698 227786 12934
rect 228022 12698 228204 12934
rect 209604 -7022 209786 -6786
rect 210022 -7022 210204 -6786
rect 209604 -7106 210204 -7022
rect 209604 -7342 209786 -7106
rect 210022 -7342 210204 -7106
rect 209604 -7364 210204 -7342
rect 227604 -5866 228204 12698
rect 234804 488454 235404 523898
rect 238404 672054 239004 707042
rect 238404 671818 238586 672054
rect 238822 671818 239004 672054
rect 238404 671734 239004 671818
rect 238404 671498 238586 671734
rect 238822 671498 239004 671734
rect 238404 636054 239004 671498
rect 238404 635818 238586 636054
rect 238822 635818 239004 636054
rect 238404 635734 239004 635818
rect 238404 635498 238586 635734
rect 238822 635498 239004 635734
rect 238404 600054 239004 635498
rect 238404 599818 238586 600054
rect 238822 599818 239004 600054
rect 238404 599734 239004 599818
rect 238404 599498 238586 599734
rect 238822 599498 239004 599734
rect 238404 564054 239004 599498
rect 238404 563818 238586 564054
rect 238822 563818 239004 564054
rect 238404 563734 239004 563818
rect 238404 563498 238586 563734
rect 238822 563498 239004 563734
rect 238404 528054 239004 563498
rect 238404 527818 238586 528054
rect 238822 527818 239004 528054
rect 238404 527734 239004 527818
rect 238404 527498 238586 527734
rect 238822 527498 239004 527734
rect 236499 519348 236565 519349
rect 236499 519284 236500 519348
rect 236564 519284 236565 519348
rect 236499 519283 236565 519284
rect 236502 518397 236562 519283
rect 236683 519212 236749 519213
rect 236683 519148 236684 519212
rect 236748 519148 236749 519212
rect 236683 519147 236749 519148
rect 236315 518396 236381 518397
rect 236315 518332 236316 518396
rect 236380 518332 236381 518396
rect 236315 518331 236381 518332
rect 236499 518396 236565 518397
rect 236499 518332 236500 518396
rect 236564 518332 236565 518396
rect 236499 518331 236565 518332
rect 236318 518125 236378 518331
rect 236315 518124 236381 518125
rect 236315 518060 236316 518124
rect 236380 518060 236381 518124
rect 236315 518059 236381 518060
rect 236686 517989 236746 519147
rect 236867 519076 236933 519077
rect 236867 519012 236868 519076
rect 236932 519012 236933 519076
rect 236867 519011 236933 519012
rect 236870 518669 236930 519011
rect 236867 518668 236933 518669
rect 236867 518604 236868 518668
rect 236932 518604 236933 518668
rect 236867 518603 236933 518604
rect 236683 517988 236749 517989
rect 236683 517924 236684 517988
rect 236748 517924 236749 517988
rect 236683 517923 236749 517924
rect 234804 488218 234986 488454
rect 235222 488218 235404 488454
rect 234804 488134 235404 488218
rect 234804 487898 234986 488134
rect 235222 487898 235404 488134
rect 234804 452454 235404 487898
rect 234804 452218 234986 452454
rect 235222 452218 235404 452454
rect 234804 452134 235404 452218
rect 234804 451898 234986 452134
rect 235222 451898 235404 452134
rect 234804 416454 235404 451898
rect 234804 416218 234986 416454
rect 235222 416218 235404 416454
rect 234804 416134 235404 416218
rect 234804 415898 234986 416134
rect 235222 415898 235404 416134
rect 234804 380454 235404 415898
rect 234804 380218 234986 380454
rect 235222 380218 235404 380454
rect 234804 380134 235404 380218
rect 234804 379898 234986 380134
rect 235222 379898 235404 380134
rect 234804 344454 235404 379898
rect 234804 344218 234986 344454
rect 235222 344218 235404 344454
rect 234804 344134 235404 344218
rect 234804 343898 234986 344134
rect 235222 343898 235404 344134
rect 234804 308454 235404 343898
rect 234804 308218 234986 308454
rect 235222 308218 235404 308454
rect 234804 308134 235404 308218
rect 234804 307898 234986 308134
rect 235222 307898 235404 308134
rect 234804 272454 235404 307898
rect 234804 272218 234986 272454
rect 235222 272218 235404 272454
rect 234804 272134 235404 272218
rect 234804 271898 234986 272134
rect 235222 271898 235404 272134
rect 234804 236454 235404 271898
rect 234804 236218 234986 236454
rect 235222 236218 235404 236454
rect 234804 236134 235404 236218
rect 234804 235898 234986 236134
rect 235222 235898 235404 236134
rect 234804 200454 235404 235898
rect 234804 200218 234986 200454
rect 235222 200218 235404 200454
rect 234804 200134 235404 200218
rect 234804 199898 234986 200134
rect 235222 199898 235404 200134
rect 234804 164454 235404 199898
rect 234804 164218 234986 164454
rect 235222 164218 235404 164454
rect 234804 164134 235404 164218
rect 234804 163898 234986 164134
rect 235222 163898 235404 164134
rect 234804 128454 235404 163898
rect 234804 128218 234986 128454
rect 235222 128218 235404 128454
rect 234804 128134 235404 128218
rect 234804 127898 234986 128134
rect 235222 127898 235404 128134
rect 234804 92454 235404 127898
rect 234804 92218 234986 92454
rect 235222 92218 235404 92454
rect 234804 92134 235404 92218
rect 234804 91898 234986 92134
rect 235222 91898 235404 92134
rect 234804 56454 235404 91898
rect 234804 56218 234986 56454
rect 235222 56218 235404 56454
rect 234804 56134 235404 56218
rect 234804 55898 234986 56134
rect 235222 55898 235404 56134
rect 234804 20454 235404 55898
rect 234804 20218 234986 20454
rect 235222 20218 235404 20454
rect 234804 20134 235404 20218
rect 234804 19898 234986 20134
rect 235222 19898 235404 20134
rect 234804 -1266 235404 19898
rect 234804 -1502 234986 -1266
rect 235222 -1502 235404 -1266
rect 234804 -1586 235404 -1502
rect 234804 -1822 234986 -1586
rect 235222 -1822 235404 -1586
rect 234804 -1844 235404 -1822
rect 238404 492054 239004 527498
rect 242004 675654 242604 708882
rect 242004 675418 242186 675654
rect 242422 675418 242604 675654
rect 242004 675334 242604 675418
rect 242004 675098 242186 675334
rect 242422 675098 242604 675334
rect 242004 639654 242604 675098
rect 242004 639418 242186 639654
rect 242422 639418 242604 639654
rect 242004 639334 242604 639418
rect 242004 639098 242186 639334
rect 242422 639098 242604 639334
rect 242004 603654 242604 639098
rect 242004 603418 242186 603654
rect 242422 603418 242604 603654
rect 242004 603334 242604 603418
rect 242004 603098 242186 603334
rect 242422 603098 242604 603334
rect 242004 567654 242604 603098
rect 242004 567418 242186 567654
rect 242422 567418 242604 567654
rect 242004 567334 242604 567418
rect 242004 567098 242186 567334
rect 242422 567098 242604 567334
rect 242004 531654 242604 567098
rect 242004 531418 242186 531654
rect 242422 531418 242604 531654
rect 242004 531334 242604 531418
rect 242004 531098 242186 531334
rect 242422 531098 242604 531334
rect 241467 519212 241533 519213
rect 241467 519148 241468 519212
rect 241532 519148 241533 519212
rect 241467 519147 241533 519148
rect 241470 518805 241530 519147
rect 241467 518804 241533 518805
rect 241467 518740 241468 518804
rect 241532 518740 241533 518804
rect 241467 518739 241533 518740
rect 238404 491818 238586 492054
rect 238822 491818 239004 492054
rect 238404 491734 239004 491818
rect 238404 491498 238586 491734
rect 238822 491498 239004 491734
rect 238404 456054 239004 491498
rect 238404 455818 238586 456054
rect 238822 455818 239004 456054
rect 238404 455734 239004 455818
rect 238404 455498 238586 455734
rect 238822 455498 239004 455734
rect 238404 420054 239004 455498
rect 238404 419818 238586 420054
rect 238822 419818 239004 420054
rect 238404 419734 239004 419818
rect 238404 419498 238586 419734
rect 238822 419498 239004 419734
rect 238404 384054 239004 419498
rect 238404 383818 238586 384054
rect 238822 383818 239004 384054
rect 238404 383734 239004 383818
rect 238404 383498 238586 383734
rect 238822 383498 239004 383734
rect 238404 348054 239004 383498
rect 238404 347818 238586 348054
rect 238822 347818 239004 348054
rect 238404 347734 239004 347818
rect 238404 347498 238586 347734
rect 238822 347498 239004 347734
rect 238404 312054 239004 347498
rect 238404 311818 238586 312054
rect 238822 311818 239004 312054
rect 238404 311734 239004 311818
rect 238404 311498 238586 311734
rect 238822 311498 239004 311734
rect 238404 276054 239004 311498
rect 238404 275818 238586 276054
rect 238822 275818 239004 276054
rect 238404 275734 239004 275818
rect 238404 275498 238586 275734
rect 238822 275498 239004 275734
rect 238404 240054 239004 275498
rect 238404 239818 238586 240054
rect 238822 239818 239004 240054
rect 238404 239734 239004 239818
rect 238404 239498 238586 239734
rect 238822 239498 239004 239734
rect 238404 204054 239004 239498
rect 238404 203818 238586 204054
rect 238822 203818 239004 204054
rect 238404 203734 239004 203818
rect 238404 203498 238586 203734
rect 238822 203498 239004 203734
rect 238404 168054 239004 203498
rect 238404 167818 238586 168054
rect 238822 167818 239004 168054
rect 238404 167734 239004 167818
rect 238404 167498 238586 167734
rect 238822 167498 239004 167734
rect 238404 132054 239004 167498
rect 238404 131818 238586 132054
rect 238822 131818 239004 132054
rect 238404 131734 239004 131818
rect 238404 131498 238586 131734
rect 238822 131498 239004 131734
rect 238404 96054 239004 131498
rect 238404 95818 238586 96054
rect 238822 95818 239004 96054
rect 238404 95734 239004 95818
rect 238404 95498 238586 95734
rect 238822 95498 239004 95734
rect 238404 60054 239004 95498
rect 238404 59818 238586 60054
rect 238822 59818 239004 60054
rect 238404 59734 239004 59818
rect 238404 59498 238586 59734
rect 238822 59498 239004 59734
rect 238404 24054 239004 59498
rect 238404 23818 238586 24054
rect 238822 23818 239004 24054
rect 238404 23734 239004 23818
rect 238404 23498 238586 23734
rect 238822 23498 239004 23734
rect 238404 -3106 239004 23498
rect 238404 -3342 238586 -3106
rect 238822 -3342 239004 -3106
rect 238404 -3426 239004 -3342
rect 238404 -3662 238586 -3426
rect 238822 -3662 239004 -3426
rect 238404 -3684 239004 -3662
rect 242004 495654 242604 531098
rect 245604 679254 246204 710722
rect 263604 710358 264204 711300
rect 263604 710122 263786 710358
rect 264022 710122 264204 710358
rect 263604 710038 264204 710122
rect 263604 709802 263786 710038
rect 264022 709802 264204 710038
rect 260004 708518 260604 709460
rect 260004 708282 260186 708518
rect 260422 708282 260604 708518
rect 260004 708198 260604 708282
rect 260004 707962 260186 708198
rect 260422 707962 260604 708198
rect 256404 706678 257004 707620
rect 256404 706442 256586 706678
rect 256822 706442 257004 706678
rect 256404 706358 257004 706442
rect 256404 706122 256586 706358
rect 256822 706122 257004 706358
rect 245604 679018 245786 679254
rect 246022 679018 246204 679254
rect 245604 678934 246204 679018
rect 245604 678698 245786 678934
rect 246022 678698 246204 678934
rect 245604 643254 246204 678698
rect 245604 643018 245786 643254
rect 246022 643018 246204 643254
rect 245604 642934 246204 643018
rect 245604 642698 245786 642934
rect 246022 642698 246204 642934
rect 245604 607254 246204 642698
rect 245604 607018 245786 607254
rect 246022 607018 246204 607254
rect 245604 606934 246204 607018
rect 245604 606698 245786 606934
rect 246022 606698 246204 606934
rect 245604 571254 246204 606698
rect 245604 571018 245786 571254
rect 246022 571018 246204 571254
rect 245604 570934 246204 571018
rect 245604 570698 245786 570934
rect 246022 570698 246204 570934
rect 245604 535254 246204 570698
rect 245604 535018 245786 535254
rect 246022 535018 246204 535254
rect 245604 534934 246204 535018
rect 245604 534698 245786 534934
rect 246022 534698 246204 534934
rect 243859 518668 243925 518669
rect 243859 518666 243860 518668
rect 243310 518606 243860 518666
rect 243310 517989 243370 518606
rect 243859 518604 243860 518606
rect 243924 518604 243925 518668
rect 243859 518603 243925 518604
rect 244227 518668 244293 518669
rect 244227 518604 244228 518668
rect 244292 518604 244293 518668
rect 244227 518603 244293 518604
rect 244230 518530 244290 518603
rect 244230 518470 244474 518530
rect 244414 517989 244474 518470
rect 243307 517988 243373 517989
rect 243307 517924 243308 517988
rect 243372 517924 243373 517988
rect 243675 517988 243741 517989
rect 243675 517938 243676 517988
rect 243740 517938 243741 517988
rect 244227 517988 244293 517989
rect 243307 517923 243373 517924
rect 244227 517924 244228 517988
rect 244292 517924 244293 517988
rect 244227 517923 244293 517924
rect 244411 517988 244477 517989
rect 244411 517924 244412 517988
rect 244476 517924 244477 517988
rect 244411 517923 244477 517924
rect 244230 517850 244290 517923
rect 244230 517790 244694 517850
rect 242004 495418 242186 495654
rect 242422 495418 242604 495654
rect 242004 495334 242604 495418
rect 242004 495098 242186 495334
rect 242422 495098 242604 495334
rect 242004 459654 242604 495098
rect 242004 459418 242186 459654
rect 242422 459418 242604 459654
rect 242004 459334 242604 459418
rect 242004 459098 242186 459334
rect 242422 459098 242604 459334
rect 242004 423654 242604 459098
rect 242004 423418 242186 423654
rect 242422 423418 242604 423654
rect 242004 423334 242604 423418
rect 242004 423098 242186 423334
rect 242422 423098 242604 423334
rect 242004 387654 242604 423098
rect 242004 387418 242186 387654
rect 242422 387418 242604 387654
rect 242004 387334 242604 387418
rect 242004 387098 242186 387334
rect 242422 387098 242604 387334
rect 242004 351654 242604 387098
rect 242004 351418 242186 351654
rect 242422 351418 242604 351654
rect 242004 351334 242604 351418
rect 242004 351098 242186 351334
rect 242422 351098 242604 351334
rect 242004 315654 242604 351098
rect 242004 315418 242186 315654
rect 242422 315418 242604 315654
rect 242004 315334 242604 315418
rect 242004 315098 242186 315334
rect 242422 315098 242604 315334
rect 242004 279654 242604 315098
rect 242004 279418 242186 279654
rect 242422 279418 242604 279654
rect 242004 279334 242604 279418
rect 242004 279098 242186 279334
rect 242422 279098 242604 279334
rect 242004 243654 242604 279098
rect 242004 243418 242186 243654
rect 242422 243418 242604 243654
rect 242004 243334 242604 243418
rect 242004 243098 242186 243334
rect 242422 243098 242604 243334
rect 242004 207654 242604 243098
rect 242004 207418 242186 207654
rect 242422 207418 242604 207654
rect 242004 207334 242604 207418
rect 242004 207098 242186 207334
rect 242422 207098 242604 207334
rect 242004 171654 242604 207098
rect 242004 171418 242186 171654
rect 242422 171418 242604 171654
rect 242004 171334 242604 171418
rect 242004 171098 242186 171334
rect 242422 171098 242604 171334
rect 242004 135654 242604 171098
rect 242004 135418 242186 135654
rect 242422 135418 242604 135654
rect 242004 135334 242604 135418
rect 242004 135098 242186 135334
rect 242422 135098 242604 135334
rect 242004 99654 242604 135098
rect 242004 99418 242186 99654
rect 242422 99418 242604 99654
rect 242004 99334 242604 99418
rect 242004 99098 242186 99334
rect 242422 99098 242604 99334
rect 242004 63654 242604 99098
rect 242004 63418 242186 63654
rect 242422 63418 242604 63654
rect 242004 63334 242604 63418
rect 242004 63098 242186 63334
rect 242422 63098 242604 63334
rect 242004 27654 242604 63098
rect 242004 27418 242186 27654
rect 242422 27418 242604 27654
rect 242004 27334 242604 27418
rect 242004 27098 242186 27334
rect 242422 27098 242604 27334
rect 242004 -4946 242604 27098
rect 242004 -5182 242186 -4946
rect 242422 -5182 242604 -4946
rect 242004 -5266 242604 -5182
rect 242004 -5502 242186 -5266
rect 242422 -5502 242604 -5266
rect 242004 -5524 242604 -5502
rect 245604 499254 246204 534698
rect 252804 704838 253404 705780
rect 252804 704602 252986 704838
rect 253222 704602 253404 704838
rect 252804 704518 253404 704602
rect 252804 704282 252986 704518
rect 253222 704282 253404 704518
rect 252804 686454 253404 704282
rect 252804 686218 252986 686454
rect 253222 686218 253404 686454
rect 252804 686134 253404 686218
rect 252804 685898 252986 686134
rect 253222 685898 253404 686134
rect 252804 650454 253404 685898
rect 252804 650218 252986 650454
rect 253222 650218 253404 650454
rect 252804 650134 253404 650218
rect 252804 649898 252986 650134
rect 253222 649898 253404 650134
rect 252804 614454 253404 649898
rect 252804 614218 252986 614454
rect 253222 614218 253404 614454
rect 252804 614134 253404 614218
rect 252804 613898 252986 614134
rect 253222 613898 253404 614134
rect 252804 578454 253404 613898
rect 252804 578218 252986 578454
rect 253222 578218 253404 578454
rect 252804 578134 253404 578218
rect 252804 577898 252986 578134
rect 253222 577898 253404 578134
rect 252804 542454 253404 577898
rect 252804 542218 252986 542454
rect 253222 542218 253404 542454
rect 252804 542134 253404 542218
rect 252804 541898 252986 542134
rect 253222 541898 253404 542134
rect 246435 519212 246501 519213
rect 246435 519148 246436 519212
rect 246500 519148 246501 519212
rect 246435 519147 246501 519148
rect 246438 518805 246498 519147
rect 246435 518804 246501 518805
rect 246435 518740 246436 518804
rect 246500 518740 246501 518804
rect 246435 518739 246501 518740
rect 245604 499018 245786 499254
rect 246022 499018 246204 499254
rect 245604 498934 246204 499018
rect 245604 498698 245786 498934
rect 246022 498698 246204 498934
rect 245604 463254 246204 498698
rect 245604 463018 245786 463254
rect 246022 463018 246204 463254
rect 245604 462934 246204 463018
rect 245604 462698 245786 462934
rect 246022 462698 246204 462934
rect 245604 427254 246204 462698
rect 245604 427018 245786 427254
rect 246022 427018 246204 427254
rect 245604 426934 246204 427018
rect 245604 426698 245786 426934
rect 246022 426698 246204 426934
rect 245604 391254 246204 426698
rect 245604 391018 245786 391254
rect 246022 391018 246204 391254
rect 245604 390934 246204 391018
rect 245604 390698 245786 390934
rect 246022 390698 246204 390934
rect 245604 355254 246204 390698
rect 245604 355018 245786 355254
rect 246022 355018 246204 355254
rect 245604 354934 246204 355018
rect 245604 354698 245786 354934
rect 246022 354698 246204 354934
rect 245604 319254 246204 354698
rect 245604 319018 245786 319254
rect 246022 319018 246204 319254
rect 245604 318934 246204 319018
rect 245604 318698 245786 318934
rect 246022 318698 246204 318934
rect 245604 283254 246204 318698
rect 245604 283018 245786 283254
rect 246022 283018 246204 283254
rect 245604 282934 246204 283018
rect 245604 282698 245786 282934
rect 246022 282698 246204 282934
rect 245604 247254 246204 282698
rect 245604 247018 245786 247254
rect 246022 247018 246204 247254
rect 245604 246934 246204 247018
rect 245604 246698 245786 246934
rect 246022 246698 246204 246934
rect 245604 211254 246204 246698
rect 245604 211018 245786 211254
rect 246022 211018 246204 211254
rect 245604 210934 246204 211018
rect 245604 210698 245786 210934
rect 246022 210698 246204 210934
rect 245604 175254 246204 210698
rect 245604 175018 245786 175254
rect 246022 175018 246204 175254
rect 245604 174934 246204 175018
rect 245604 174698 245786 174934
rect 246022 174698 246204 174934
rect 245604 139254 246204 174698
rect 245604 139018 245786 139254
rect 246022 139018 246204 139254
rect 245604 138934 246204 139018
rect 245604 138698 245786 138934
rect 246022 138698 246204 138934
rect 245604 103254 246204 138698
rect 245604 103018 245786 103254
rect 246022 103018 246204 103254
rect 245604 102934 246204 103018
rect 245604 102698 245786 102934
rect 246022 102698 246204 102934
rect 245604 67254 246204 102698
rect 245604 67018 245786 67254
rect 246022 67018 246204 67254
rect 245604 66934 246204 67018
rect 245604 66698 245786 66934
rect 246022 66698 246204 66934
rect 245604 31254 246204 66698
rect 245604 31018 245786 31254
rect 246022 31018 246204 31254
rect 245604 30934 246204 31018
rect 245604 30698 245786 30934
rect 246022 30698 246204 30934
rect 227604 -6102 227786 -5866
rect 228022 -6102 228204 -5866
rect 227604 -6186 228204 -6102
rect 227604 -6422 227786 -6186
rect 228022 -6422 228204 -6186
rect 227604 -7364 228204 -6422
rect 245604 -6786 246204 30698
rect 252804 506454 253404 541898
rect 256404 690054 257004 706122
rect 256404 689818 256586 690054
rect 256822 689818 257004 690054
rect 256404 689734 257004 689818
rect 256404 689498 256586 689734
rect 256822 689498 257004 689734
rect 256404 654054 257004 689498
rect 256404 653818 256586 654054
rect 256822 653818 257004 654054
rect 256404 653734 257004 653818
rect 256404 653498 256586 653734
rect 256822 653498 257004 653734
rect 256404 618054 257004 653498
rect 256404 617818 256586 618054
rect 256822 617818 257004 618054
rect 256404 617734 257004 617818
rect 256404 617498 256586 617734
rect 256822 617498 257004 617734
rect 256404 582054 257004 617498
rect 256404 581818 256586 582054
rect 256822 581818 257004 582054
rect 256404 581734 257004 581818
rect 256404 581498 256586 581734
rect 256822 581498 257004 581734
rect 256404 546054 257004 581498
rect 256404 545818 256586 546054
rect 256822 545818 257004 546054
rect 256404 545734 257004 545818
rect 256404 545498 256586 545734
rect 256822 545498 257004 545734
rect 253611 518940 253677 518941
rect 253611 518876 253612 518940
rect 253676 518876 253677 518940
rect 253611 518875 253677 518876
rect 253614 518669 253674 518875
rect 253611 518668 253677 518669
rect 253611 518604 253612 518668
rect 253676 518604 253677 518668
rect 253611 518603 253677 518604
rect 253795 518668 253861 518669
rect 253795 518604 253796 518668
rect 253860 518604 253861 518668
rect 253795 518603 253861 518604
rect 253798 517989 253858 518603
rect 253795 517988 253861 517989
rect 253795 517924 253796 517988
rect 253860 517924 253861 517988
rect 254163 517988 254229 517989
rect 254163 517938 254164 517988
rect 254228 517938 254229 517988
rect 253795 517923 253861 517924
rect 252804 506218 252986 506454
rect 253222 506218 253404 506454
rect 252804 506134 253404 506218
rect 252804 505898 252986 506134
rect 253222 505898 253404 506134
rect 252804 470454 253404 505898
rect 252804 470218 252986 470454
rect 253222 470218 253404 470454
rect 252804 470134 253404 470218
rect 252804 469898 252986 470134
rect 253222 469898 253404 470134
rect 252804 434454 253404 469898
rect 252804 434218 252986 434454
rect 253222 434218 253404 434454
rect 252804 434134 253404 434218
rect 252804 433898 252986 434134
rect 253222 433898 253404 434134
rect 252804 398454 253404 433898
rect 252804 398218 252986 398454
rect 253222 398218 253404 398454
rect 252804 398134 253404 398218
rect 252804 397898 252986 398134
rect 253222 397898 253404 398134
rect 252804 362454 253404 397898
rect 252804 362218 252986 362454
rect 253222 362218 253404 362454
rect 252804 362134 253404 362218
rect 252804 361898 252986 362134
rect 253222 361898 253404 362134
rect 252804 326454 253404 361898
rect 252804 326218 252986 326454
rect 253222 326218 253404 326454
rect 252804 326134 253404 326218
rect 252804 325898 252986 326134
rect 253222 325898 253404 326134
rect 252804 290454 253404 325898
rect 252804 290218 252986 290454
rect 253222 290218 253404 290454
rect 252804 290134 253404 290218
rect 252804 289898 252986 290134
rect 253222 289898 253404 290134
rect 252804 254454 253404 289898
rect 252804 254218 252986 254454
rect 253222 254218 253404 254454
rect 252804 254134 253404 254218
rect 252804 253898 252986 254134
rect 253222 253898 253404 254134
rect 252804 218454 253404 253898
rect 252804 218218 252986 218454
rect 253222 218218 253404 218454
rect 252804 218134 253404 218218
rect 252804 217898 252986 218134
rect 253222 217898 253404 218134
rect 252804 182454 253404 217898
rect 252804 182218 252986 182454
rect 253222 182218 253404 182454
rect 252804 182134 253404 182218
rect 252804 181898 252986 182134
rect 253222 181898 253404 182134
rect 252804 146454 253404 181898
rect 252804 146218 252986 146454
rect 253222 146218 253404 146454
rect 252804 146134 253404 146218
rect 252804 145898 252986 146134
rect 253222 145898 253404 146134
rect 252804 110454 253404 145898
rect 252804 110218 252986 110454
rect 253222 110218 253404 110454
rect 252804 110134 253404 110218
rect 252804 109898 252986 110134
rect 253222 109898 253404 110134
rect 252804 74454 253404 109898
rect 252804 74218 252986 74454
rect 253222 74218 253404 74454
rect 252804 74134 253404 74218
rect 252804 73898 252986 74134
rect 253222 73898 253404 74134
rect 252804 38454 253404 73898
rect 252804 38218 252986 38454
rect 253222 38218 253404 38454
rect 252804 38134 253404 38218
rect 252804 37898 252986 38134
rect 253222 37898 253404 38134
rect 252804 2454 253404 37898
rect 252804 2218 252986 2454
rect 253222 2218 253404 2454
rect 252804 2134 253404 2218
rect 252804 1898 252986 2134
rect 253222 1898 253404 2134
rect 252804 -346 253404 1898
rect 252804 -582 252986 -346
rect 253222 -582 253404 -346
rect 252804 -666 253404 -582
rect 252804 -902 252986 -666
rect 253222 -902 253404 -666
rect 252804 -1844 253404 -902
rect 256404 510054 257004 545498
rect 256404 509818 256586 510054
rect 256822 509818 257004 510054
rect 256404 509734 257004 509818
rect 256404 509498 256586 509734
rect 256822 509498 257004 509734
rect 256404 474054 257004 509498
rect 256404 473818 256586 474054
rect 256822 473818 257004 474054
rect 256404 473734 257004 473818
rect 256404 473498 256586 473734
rect 256822 473498 257004 473734
rect 256404 438054 257004 473498
rect 256404 437818 256586 438054
rect 256822 437818 257004 438054
rect 256404 437734 257004 437818
rect 256404 437498 256586 437734
rect 256822 437498 257004 437734
rect 256404 402054 257004 437498
rect 256404 401818 256586 402054
rect 256822 401818 257004 402054
rect 256404 401734 257004 401818
rect 256404 401498 256586 401734
rect 256822 401498 257004 401734
rect 256404 366054 257004 401498
rect 256404 365818 256586 366054
rect 256822 365818 257004 366054
rect 256404 365734 257004 365818
rect 256404 365498 256586 365734
rect 256822 365498 257004 365734
rect 256404 330054 257004 365498
rect 256404 329818 256586 330054
rect 256822 329818 257004 330054
rect 256404 329734 257004 329818
rect 256404 329498 256586 329734
rect 256822 329498 257004 329734
rect 256404 294054 257004 329498
rect 256404 293818 256586 294054
rect 256822 293818 257004 294054
rect 256404 293734 257004 293818
rect 256404 293498 256586 293734
rect 256822 293498 257004 293734
rect 256404 258054 257004 293498
rect 256404 257818 256586 258054
rect 256822 257818 257004 258054
rect 256404 257734 257004 257818
rect 256404 257498 256586 257734
rect 256822 257498 257004 257734
rect 256404 222054 257004 257498
rect 256404 221818 256586 222054
rect 256822 221818 257004 222054
rect 256404 221734 257004 221818
rect 256404 221498 256586 221734
rect 256822 221498 257004 221734
rect 256404 186054 257004 221498
rect 256404 185818 256586 186054
rect 256822 185818 257004 186054
rect 256404 185734 257004 185818
rect 256404 185498 256586 185734
rect 256822 185498 257004 185734
rect 256404 150054 257004 185498
rect 256404 149818 256586 150054
rect 256822 149818 257004 150054
rect 256404 149734 257004 149818
rect 256404 149498 256586 149734
rect 256822 149498 257004 149734
rect 256404 114054 257004 149498
rect 256404 113818 256586 114054
rect 256822 113818 257004 114054
rect 256404 113734 257004 113818
rect 256404 113498 256586 113734
rect 256822 113498 257004 113734
rect 256404 78054 257004 113498
rect 256404 77818 256586 78054
rect 256822 77818 257004 78054
rect 256404 77734 257004 77818
rect 256404 77498 256586 77734
rect 256822 77498 257004 77734
rect 256404 42054 257004 77498
rect 256404 41818 256586 42054
rect 256822 41818 257004 42054
rect 256404 41734 257004 41818
rect 256404 41498 256586 41734
rect 256822 41498 257004 41734
rect 256404 6054 257004 41498
rect 256404 5818 256586 6054
rect 256822 5818 257004 6054
rect 256404 5734 257004 5818
rect 256404 5498 256586 5734
rect 256822 5498 257004 5734
rect 256404 -2186 257004 5498
rect 256404 -2422 256586 -2186
rect 256822 -2422 257004 -2186
rect 256404 -2506 257004 -2422
rect 256404 -2742 256586 -2506
rect 256822 -2742 257004 -2506
rect 256404 -3684 257004 -2742
rect 260004 693654 260604 707962
rect 260004 693418 260186 693654
rect 260422 693418 260604 693654
rect 260004 693334 260604 693418
rect 260004 693098 260186 693334
rect 260422 693098 260604 693334
rect 260004 657654 260604 693098
rect 260004 657418 260186 657654
rect 260422 657418 260604 657654
rect 260004 657334 260604 657418
rect 260004 657098 260186 657334
rect 260422 657098 260604 657334
rect 260004 621654 260604 657098
rect 260004 621418 260186 621654
rect 260422 621418 260604 621654
rect 260004 621334 260604 621418
rect 260004 621098 260186 621334
rect 260422 621098 260604 621334
rect 260004 585654 260604 621098
rect 260004 585418 260186 585654
rect 260422 585418 260604 585654
rect 260004 585334 260604 585418
rect 260004 585098 260186 585334
rect 260422 585098 260604 585334
rect 260004 549654 260604 585098
rect 260004 549418 260186 549654
rect 260422 549418 260604 549654
rect 260004 549334 260604 549418
rect 260004 549098 260186 549334
rect 260422 549098 260604 549334
rect 260004 513654 260604 549098
rect 263604 697254 264204 709802
rect 281604 711278 282204 711300
rect 281604 711042 281786 711278
rect 282022 711042 282204 711278
rect 281604 710958 282204 711042
rect 281604 710722 281786 710958
rect 282022 710722 282204 710958
rect 278004 709438 278604 709460
rect 278004 709202 278186 709438
rect 278422 709202 278604 709438
rect 278004 709118 278604 709202
rect 278004 708882 278186 709118
rect 278422 708882 278604 709118
rect 274404 707598 275004 707620
rect 274404 707362 274586 707598
rect 274822 707362 275004 707598
rect 274404 707278 275004 707362
rect 274404 707042 274586 707278
rect 274822 707042 275004 707278
rect 263604 697018 263786 697254
rect 264022 697018 264204 697254
rect 263604 696934 264204 697018
rect 263604 696698 263786 696934
rect 264022 696698 264204 696934
rect 263604 661254 264204 696698
rect 263604 661018 263786 661254
rect 264022 661018 264204 661254
rect 263604 660934 264204 661018
rect 263604 660698 263786 660934
rect 264022 660698 264204 660934
rect 263604 625254 264204 660698
rect 270804 705758 271404 705780
rect 270804 705522 270986 705758
rect 271222 705522 271404 705758
rect 270804 705438 271404 705522
rect 270804 705202 270986 705438
rect 271222 705202 271404 705438
rect 270804 668454 271404 705202
rect 270804 668218 270986 668454
rect 271222 668218 271404 668454
rect 270804 668134 271404 668218
rect 270804 667898 270986 668134
rect 271222 667898 271404 668134
rect 267411 645828 267477 645829
rect 267411 645764 267412 645828
rect 267476 645764 267477 645828
rect 267411 645763 267477 645764
rect 267414 640253 267474 645763
rect 267411 640252 267477 640253
rect 267411 640188 267412 640252
rect 267476 640188 267477 640252
rect 267411 640187 267477 640188
rect 263604 625018 263786 625254
rect 264022 625018 264204 625254
rect 263604 624934 264204 625018
rect 263604 624698 263786 624934
rect 264022 624698 264204 624934
rect 263604 589254 264204 624698
rect 263604 589018 263786 589254
rect 264022 589018 264204 589254
rect 263604 588934 264204 589018
rect 263604 588698 263786 588934
rect 264022 588698 264204 588934
rect 263604 553254 264204 588698
rect 263604 553018 263786 553254
rect 264022 553018 264204 553254
rect 263604 552934 264204 553018
rect 263604 552698 263786 552934
rect 264022 552698 264204 552934
rect 263179 519212 263245 519213
rect 263179 519148 263180 519212
rect 263244 519148 263245 519212
rect 263179 519147 263245 519148
rect 263182 518669 263242 519147
rect 263363 519076 263429 519077
rect 263363 519012 263364 519076
rect 263428 519012 263429 519076
rect 263363 519011 263429 519012
rect 263366 518805 263426 519011
rect 263363 518804 263429 518805
rect 263363 518740 263364 518804
rect 263428 518740 263429 518804
rect 263363 518739 263429 518740
rect 263179 518668 263245 518669
rect 263179 518604 263180 518668
rect 263244 518604 263245 518668
rect 263179 518603 263245 518604
rect 260004 513418 260186 513654
rect 260422 513418 260604 513654
rect 260004 513334 260604 513418
rect 260004 513098 260186 513334
rect 260422 513098 260604 513334
rect 260004 477654 260604 513098
rect 260004 477418 260186 477654
rect 260422 477418 260604 477654
rect 260004 477334 260604 477418
rect 260004 477098 260186 477334
rect 260422 477098 260604 477334
rect 260004 441654 260604 477098
rect 260004 441418 260186 441654
rect 260422 441418 260604 441654
rect 260004 441334 260604 441418
rect 260004 441098 260186 441334
rect 260422 441098 260604 441334
rect 260004 405654 260604 441098
rect 260004 405418 260186 405654
rect 260422 405418 260604 405654
rect 260004 405334 260604 405418
rect 260004 405098 260186 405334
rect 260422 405098 260604 405334
rect 260004 369654 260604 405098
rect 260004 369418 260186 369654
rect 260422 369418 260604 369654
rect 260004 369334 260604 369418
rect 260004 369098 260186 369334
rect 260422 369098 260604 369334
rect 260004 333654 260604 369098
rect 260004 333418 260186 333654
rect 260422 333418 260604 333654
rect 260004 333334 260604 333418
rect 260004 333098 260186 333334
rect 260422 333098 260604 333334
rect 260004 297654 260604 333098
rect 260004 297418 260186 297654
rect 260422 297418 260604 297654
rect 260004 297334 260604 297418
rect 260004 297098 260186 297334
rect 260422 297098 260604 297334
rect 260004 261654 260604 297098
rect 260004 261418 260186 261654
rect 260422 261418 260604 261654
rect 260004 261334 260604 261418
rect 260004 261098 260186 261334
rect 260422 261098 260604 261334
rect 260004 225654 260604 261098
rect 260004 225418 260186 225654
rect 260422 225418 260604 225654
rect 260004 225334 260604 225418
rect 260004 225098 260186 225334
rect 260422 225098 260604 225334
rect 260004 189654 260604 225098
rect 260004 189418 260186 189654
rect 260422 189418 260604 189654
rect 260004 189334 260604 189418
rect 260004 189098 260186 189334
rect 260422 189098 260604 189334
rect 260004 153654 260604 189098
rect 260004 153418 260186 153654
rect 260422 153418 260604 153654
rect 260004 153334 260604 153418
rect 260004 153098 260186 153334
rect 260422 153098 260604 153334
rect 260004 117654 260604 153098
rect 260004 117418 260186 117654
rect 260422 117418 260604 117654
rect 260004 117334 260604 117418
rect 260004 117098 260186 117334
rect 260422 117098 260604 117334
rect 260004 81654 260604 117098
rect 260004 81418 260186 81654
rect 260422 81418 260604 81654
rect 260004 81334 260604 81418
rect 260004 81098 260186 81334
rect 260422 81098 260604 81334
rect 260004 45654 260604 81098
rect 260004 45418 260186 45654
rect 260422 45418 260604 45654
rect 260004 45334 260604 45418
rect 260004 45098 260186 45334
rect 260422 45098 260604 45334
rect 260004 9654 260604 45098
rect 260004 9418 260186 9654
rect 260422 9418 260604 9654
rect 260004 9334 260604 9418
rect 260004 9098 260186 9334
rect 260422 9098 260604 9334
rect 260004 -4026 260604 9098
rect 260004 -4262 260186 -4026
rect 260422 -4262 260604 -4026
rect 260004 -4346 260604 -4262
rect 260004 -4582 260186 -4346
rect 260422 -4582 260604 -4346
rect 260004 -5524 260604 -4582
rect 263604 517254 264204 552698
rect 270804 632454 271404 667898
rect 270804 632218 270986 632454
rect 271222 632218 271404 632454
rect 270804 632134 271404 632218
rect 270804 631898 270986 632134
rect 271222 631898 271404 632134
rect 270804 596454 271404 631898
rect 270804 596218 270986 596454
rect 271222 596218 271404 596454
rect 270804 596134 271404 596218
rect 270804 595898 270986 596134
rect 271222 595898 271404 596134
rect 270804 560454 271404 595898
rect 270804 560218 270986 560454
rect 271222 560218 271404 560454
rect 270804 560134 271404 560218
rect 270804 559898 270986 560134
rect 271222 559898 271404 560134
rect 270804 524454 271404 559898
rect 270804 524218 270986 524454
rect 271222 524218 271404 524454
rect 270804 524134 271404 524218
rect 270804 523898 270986 524134
rect 271222 523898 271404 524134
rect 265571 519212 265637 519213
rect 265571 519148 265572 519212
rect 265636 519148 265637 519212
rect 265571 519147 265637 519148
rect 265574 517989 265634 519147
rect 264467 517988 264533 517989
rect 264467 517938 264468 517988
rect 264532 517938 264533 517988
rect 265571 517988 265637 517989
rect 265571 517924 265572 517988
rect 265636 517924 265637 517988
rect 265571 517923 265637 517924
rect 263604 517018 263786 517254
rect 264022 517018 264204 517254
rect 263604 516934 264204 517018
rect 263604 516698 263786 516934
rect 264022 516698 264204 516934
rect 263604 481254 264204 516698
rect 263604 481018 263786 481254
rect 264022 481018 264204 481254
rect 263604 480934 264204 481018
rect 263604 480698 263786 480934
rect 264022 480698 264204 480934
rect 263604 445254 264204 480698
rect 263604 445018 263786 445254
rect 264022 445018 264204 445254
rect 263604 444934 264204 445018
rect 263604 444698 263786 444934
rect 264022 444698 264204 444934
rect 263604 409254 264204 444698
rect 263604 409018 263786 409254
rect 264022 409018 264204 409254
rect 263604 408934 264204 409018
rect 263604 408698 263786 408934
rect 264022 408698 264204 408934
rect 263604 373254 264204 408698
rect 263604 373018 263786 373254
rect 264022 373018 264204 373254
rect 263604 372934 264204 373018
rect 263604 372698 263786 372934
rect 264022 372698 264204 372934
rect 263604 337254 264204 372698
rect 263604 337018 263786 337254
rect 264022 337018 264204 337254
rect 263604 336934 264204 337018
rect 263604 336698 263786 336934
rect 264022 336698 264204 336934
rect 263604 301254 264204 336698
rect 263604 301018 263786 301254
rect 264022 301018 264204 301254
rect 263604 300934 264204 301018
rect 263604 300698 263786 300934
rect 264022 300698 264204 300934
rect 263604 265254 264204 300698
rect 263604 265018 263786 265254
rect 264022 265018 264204 265254
rect 263604 264934 264204 265018
rect 263604 264698 263786 264934
rect 264022 264698 264204 264934
rect 263604 229254 264204 264698
rect 263604 229018 263786 229254
rect 264022 229018 264204 229254
rect 263604 228934 264204 229018
rect 263604 228698 263786 228934
rect 264022 228698 264204 228934
rect 263604 193254 264204 228698
rect 263604 193018 263786 193254
rect 264022 193018 264204 193254
rect 263604 192934 264204 193018
rect 263604 192698 263786 192934
rect 264022 192698 264204 192934
rect 263604 157254 264204 192698
rect 263604 157018 263786 157254
rect 264022 157018 264204 157254
rect 263604 156934 264204 157018
rect 263604 156698 263786 156934
rect 264022 156698 264204 156934
rect 263604 121254 264204 156698
rect 263604 121018 263786 121254
rect 264022 121018 264204 121254
rect 263604 120934 264204 121018
rect 263604 120698 263786 120934
rect 264022 120698 264204 120934
rect 263604 85254 264204 120698
rect 263604 85018 263786 85254
rect 264022 85018 264204 85254
rect 263604 84934 264204 85018
rect 263604 84698 263786 84934
rect 264022 84698 264204 84934
rect 263604 49254 264204 84698
rect 263604 49018 263786 49254
rect 264022 49018 264204 49254
rect 263604 48934 264204 49018
rect 263604 48698 263786 48934
rect 264022 48698 264204 48934
rect 263604 13254 264204 48698
rect 263604 13018 263786 13254
rect 264022 13018 264204 13254
rect 263604 12934 264204 13018
rect 263604 12698 263786 12934
rect 264022 12698 264204 12934
rect 245604 -7022 245786 -6786
rect 246022 -7022 246204 -6786
rect 245604 -7106 246204 -7022
rect 245604 -7342 245786 -7106
rect 246022 -7342 246204 -7106
rect 245604 -7364 246204 -7342
rect 263604 -5866 264204 12698
rect 270804 488454 271404 523898
rect 274404 672054 275004 707042
rect 274404 671818 274586 672054
rect 274822 671818 275004 672054
rect 274404 671734 275004 671818
rect 274404 671498 274586 671734
rect 274822 671498 275004 671734
rect 274404 636054 275004 671498
rect 274404 635818 274586 636054
rect 274822 635818 275004 636054
rect 274404 635734 275004 635818
rect 274404 635498 274586 635734
rect 274822 635498 275004 635734
rect 274404 600054 275004 635498
rect 274404 599818 274586 600054
rect 274822 599818 275004 600054
rect 274404 599734 275004 599818
rect 274404 599498 274586 599734
rect 274822 599498 275004 599734
rect 274404 564054 275004 599498
rect 274404 563818 274586 564054
rect 274822 563818 275004 564054
rect 274404 563734 275004 563818
rect 274404 563498 274586 563734
rect 274822 563498 275004 563734
rect 274404 528054 275004 563498
rect 274404 527818 274586 528054
rect 274822 527818 275004 528054
rect 274404 527734 275004 527818
rect 274404 527498 274586 527734
rect 274822 527498 275004 527734
rect 272931 519076 272997 519077
rect 272931 519012 272932 519076
rect 272996 519012 272997 519076
rect 272931 519011 272997 519012
rect 272934 518669 272994 519011
rect 272931 518668 272997 518669
rect 272931 518604 272932 518668
rect 272996 518604 272997 518668
rect 272931 518603 272997 518604
rect 273115 518668 273181 518669
rect 273115 518604 273116 518668
rect 273180 518604 273181 518668
rect 273115 518603 273181 518604
rect 273118 517989 273178 518603
rect 273115 517988 273181 517989
rect 273115 517924 273116 517988
rect 273180 517924 273181 517988
rect 273483 517988 273549 517989
rect 273483 517938 273484 517988
rect 273548 517938 273549 517988
rect 273115 517923 273181 517924
rect 270804 488218 270986 488454
rect 271222 488218 271404 488454
rect 270804 488134 271404 488218
rect 270804 487898 270986 488134
rect 271222 487898 271404 488134
rect 270804 452454 271404 487898
rect 270804 452218 270986 452454
rect 271222 452218 271404 452454
rect 270804 452134 271404 452218
rect 270804 451898 270986 452134
rect 271222 451898 271404 452134
rect 270804 416454 271404 451898
rect 270804 416218 270986 416454
rect 271222 416218 271404 416454
rect 270804 416134 271404 416218
rect 270804 415898 270986 416134
rect 271222 415898 271404 416134
rect 270804 380454 271404 415898
rect 270804 380218 270986 380454
rect 271222 380218 271404 380454
rect 270804 380134 271404 380218
rect 270804 379898 270986 380134
rect 271222 379898 271404 380134
rect 270804 344454 271404 379898
rect 270804 344218 270986 344454
rect 271222 344218 271404 344454
rect 270804 344134 271404 344218
rect 270804 343898 270986 344134
rect 271222 343898 271404 344134
rect 270804 308454 271404 343898
rect 270804 308218 270986 308454
rect 271222 308218 271404 308454
rect 270804 308134 271404 308218
rect 270804 307898 270986 308134
rect 271222 307898 271404 308134
rect 270804 272454 271404 307898
rect 270804 272218 270986 272454
rect 271222 272218 271404 272454
rect 270804 272134 271404 272218
rect 270804 271898 270986 272134
rect 271222 271898 271404 272134
rect 270804 236454 271404 271898
rect 270804 236218 270986 236454
rect 271222 236218 271404 236454
rect 270804 236134 271404 236218
rect 270804 235898 270986 236134
rect 271222 235898 271404 236134
rect 270804 200454 271404 235898
rect 270804 200218 270986 200454
rect 271222 200218 271404 200454
rect 270804 200134 271404 200218
rect 270804 199898 270986 200134
rect 271222 199898 271404 200134
rect 270804 164454 271404 199898
rect 270804 164218 270986 164454
rect 271222 164218 271404 164454
rect 270804 164134 271404 164218
rect 270804 163898 270986 164134
rect 271222 163898 271404 164134
rect 270804 128454 271404 163898
rect 270804 128218 270986 128454
rect 271222 128218 271404 128454
rect 270804 128134 271404 128218
rect 270804 127898 270986 128134
rect 271222 127898 271404 128134
rect 270804 92454 271404 127898
rect 270804 92218 270986 92454
rect 271222 92218 271404 92454
rect 270804 92134 271404 92218
rect 270804 91898 270986 92134
rect 271222 91898 271404 92134
rect 270804 56454 271404 91898
rect 270804 56218 270986 56454
rect 271222 56218 271404 56454
rect 270804 56134 271404 56218
rect 270804 55898 270986 56134
rect 271222 55898 271404 56134
rect 270804 20454 271404 55898
rect 270804 20218 270986 20454
rect 271222 20218 271404 20454
rect 270804 20134 271404 20218
rect 270804 19898 270986 20134
rect 271222 19898 271404 20134
rect 270804 -1266 271404 19898
rect 270804 -1502 270986 -1266
rect 271222 -1502 271404 -1266
rect 270804 -1586 271404 -1502
rect 270804 -1822 270986 -1586
rect 271222 -1822 271404 -1586
rect 270804 -1844 271404 -1822
rect 274404 492054 275004 527498
rect 274404 491818 274586 492054
rect 274822 491818 275004 492054
rect 274404 491734 275004 491818
rect 274404 491498 274586 491734
rect 274822 491498 275004 491734
rect 274404 456054 275004 491498
rect 274404 455818 274586 456054
rect 274822 455818 275004 456054
rect 274404 455734 275004 455818
rect 274404 455498 274586 455734
rect 274822 455498 275004 455734
rect 274404 420054 275004 455498
rect 274404 419818 274586 420054
rect 274822 419818 275004 420054
rect 274404 419734 275004 419818
rect 274404 419498 274586 419734
rect 274822 419498 275004 419734
rect 274404 384054 275004 419498
rect 274404 383818 274586 384054
rect 274822 383818 275004 384054
rect 274404 383734 275004 383818
rect 274404 383498 274586 383734
rect 274822 383498 275004 383734
rect 274404 348054 275004 383498
rect 274404 347818 274586 348054
rect 274822 347818 275004 348054
rect 274404 347734 275004 347818
rect 274404 347498 274586 347734
rect 274822 347498 275004 347734
rect 274404 312054 275004 347498
rect 274404 311818 274586 312054
rect 274822 311818 275004 312054
rect 274404 311734 275004 311818
rect 274404 311498 274586 311734
rect 274822 311498 275004 311734
rect 274404 276054 275004 311498
rect 274404 275818 274586 276054
rect 274822 275818 275004 276054
rect 274404 275734 275004 275818
rect 274404 275498 274586 275734
rect 274822 275498 275004 275734
rect 274404 240054 275004 275498
rect 274404 239818 274586 240054
rect 274822 239818 275004 240054
rect 274404 239734 275004 239818
rect 274404 239498 274586 239734
rect 274822 239498 275004 239734
rect 274404 204054 275004 239498
rect 278004 675654 278604 708882
rect 278004 675418 278186 675654
rect 278422 675418 278604 675654
rect 278004 675334 278604 675418
rect 278004 675098 278186 675334
rect 278422 675098 278604 675334
rect 278004 639654 278604 675098
rect 278004 639418 278186 639654
rect 278422 639418 278604 639654
rect 278004 639334 278604 639418
rect 278004 639098 278186 639334
rect 278422 639098 278604 639334
rect 278004 603654 278604 639098
rect 278004 603418 278186 603654
rect 278422 603418 278604 603654
rect 278004 603334 278604 603418
rect 278004 603098 278186 603334
rect 278422 603098 278604 603334
rect 278004 567654 278604 603098
rect 278004 567418 278186 567654
rect 278422 567418 278604 567654
rect 278004 567334 278604 567418
rect 278004 567098 278186 567334
rect 278422 567098 278604 567334
rect 278004 531654 278604 567098
rect 278004 531418 278186 531654
rect 278422 531418 278604 531654
rect 278004 531334 278604 531418
rect 278004 531098 278186 531334
rect 278422 531098 278604 531334
rect 278004 495654 278604 531098
rect 281604 679254 282204 710722
rect 299604 710358 300204 711300
rect 299604 710122 299786 710358
rect 300022 710122 300204 710358
rect 299604 710038 300204 710122
rect 299604 709802 299786 710038
rect 300022 709802 300204 710038
rect 296004 708518 296604 709460
rect 296004 708282 296186 708518
rect 296422 708282 296604 708518
rect 296004 708198 296604 708282
rect 296004 707962 296186 708198
rect 296422 707962 296604 708198
rect 292404 706678 293004 707620
rect 292404 706442 292586 706678
rect 292822 706442 293004 706678
rect 292404 706358 293004 706442
rect 292404 706122 292586 706358
rect 292822 706122 293004 706358
rect 281604 679018 281786 679254
rect 282022 679018 282204 679254
rect 281604 678934 282204 679018
rect 281604 678698 281786 678934
rect 282022 678698 282204 678934
rect 281604 643254 282204 678698
rect 281604 643018 281786 643254
rect 282022 643018 282204 643254
rect 281604 642934 282204 643018
rect 281604 642698 281786 642934
rect 282022 642698 282204 642934
rect 281604 607254 282204 642698
rect 281604 607018 281786 607254
rect 282022 607018 282204 607254
rect 281604 606934 282204 607018
rect 281604 606698 281786 606934
rect 282022 606698 282204 606934
rect 281604 571254 282204 606698
rect 281604 571018 281786 571254
rect 282022 571018 282204 571254
rect 281604 570934 282204 571018
rect 281604 570698 281786 570934
rect 282022 570698 282204 570934
rect 281604 535254 282204 570698
rect 281604 535018 281786 535254
rect 282022 535018 282204 535254
rect 281604 534934 282204 535018
rect 281604 534698 281786 534934
rect 282022 534698 282204 534934
rect 280107 519348 280173 519349
rect 280107 519284 280108 519348
rect 280172 519284 280173 519348
rect 280107 519283 280173 519284
rect 280110 519077 280170 519283
rect 280107 519076 280173 519077
rect 280107 519012 280108 519076
rect 280172 519012 280173 519076
rect 280107 519011 280173 519012
rect 278004 495418 278186 495654
rect 278422 495418 278604 495654
rect 278004 495334 278604 495418
rect 278004 495098 278186 495334
rect 278422 495098 278604 495334
rect 278004 459654 278604 495098
rect 278004 459418 278186 459654
rect 278422 459418 278604 459654
rect 278004 459334 278604 459418
rect 278004 459098 278186 459334
rect 278422 459098 278604 459334
rect 278004 423654 278604 459098
rect 278004 423418 278186 423654
rect 278422 423418 278604 423654
rect 278004 423334 278604 423418
rect 278004 423098 278186 423334
rect 278422 423098 278604 423334
rect 278004 387654 278604 423098
rect 278004 387418 278186 387654
rect 278422 387418 278604 387654
rect 278004 387334 278604 387418
rect 278004 387098 278186 387334
rect 278422 387098 278604 387334
rect 278004 351654 278604 387098
rect 278004 351418 278186 351654
rect 278422 351418 278604 351654
rect 278004 351334 278604 351418
rect 278004 351098 278186 351334
rect 278422 351098 278604 351334
rect 278004 315654 278604 351098
rect 278004 315418 278186 315654
rect 278422 315418 278604 315654
rect 278004 315334 278604 315418
rect 278004 315098 278186 315334
rect 278422 315098 278604 315334
rect 278004 279654 278604 315098
rect 278004 279418 278186 279654
rect 278422 279418 278604 279654
rect 278004 279334 278604 279418
rect 278004 279098 278186 279334
rect 278422 279098 278604 279334
rect 278004 243654 278604 279098
rect 278004 243418 278186 243654
rect 278422 243418 278604 243654
rect 278004 243334 278604 243418
rect 278004 243098 278186 243334
rect 278422 243098 278604 243334
rect 275875 217972 275941 217973
rect 275875 217908 275876 217972
rect 275940 217908 275941 217972
rect 275875 217907 275941 217908
rect 275878 217701 275938 217907
rect 275875 217700 275941 217701
rect 275875 217636 275876 217700
rect 275940 217636 275941 217700
rect 275875 217635 275941 217636
rect 274404 203818 274586 204054
rect 274822 203818 275004 204054
rect 274404 203734 275004 203818
rect 274404 203498 274586 203734
rect 274822 203498 275004 203734
rect 274404 168054 275004 203498
rect 274404 167818 274586 168054
rect 274822 167818 275004 168054
rect 274404 167734 275004 167818
rect 274404 167498 274586 167734
rect 274822 167498 275004 167734
rect 274404 132054 275004 167498
rect 278004 207654 278604 243098
rect 278004 207418 278186 207654
rect 278422 207418 278604 207654
rect 278004 207334 278604 207418
rect 278004 207098 278186 207334
rect 278422 207098 278604 207334
rect 278004 171654 278604 207098
rect 278004 171418 278186 171654
rect 278422 171418 278604 171654
rect 278004 171334 278604 171418
rect 278004 171098 278186 171334
rect 278422 171098 278604 171334
rect 277163 162756 277229 162757
rect 277163 162692 277164 162756
rect 277228 162692 277229 162756
rect 277163 162691 277229 162692
rect 277166 153237 277226 162691
rect 277163 153236 277229 153237
rect 277163 153172 277164 153236
rect 277228 153172 277229 153236
rect 277163 153171 277229 153172
rect 274404 131818 274586 132054
rect 274822 131818 275004 132054
rect 274404 131734 275004 131818
rect 274404 131498 274586 131734
rect 274822 131498 275004 131734
rect 274404 96054 275004 131498
rect 274404 95818 274586 96054
rect 274822 95818 275004 96054
rect 274404 95734 275004 95818
rect 274404 95498 274586 95734
rect 274822 95498 275004 95734
rect 274404 60054 275004 95498
rect 274404 59818 274586 60054
rect 274822 59818 275004 60054
rect 274404 59734 275004 59818
rect 274404 59498 274586 59734
rect 274822 59498 275004 59734
rect 274404 24054 275004 59498
rect 274404 23818 274586 24054
rect 274822 23818 275004 24054
rect 274404 23734 275004 23818
rect 274404 23498 274586 23734
rect 274822 23498 275004 23734
rect 274404 -3106 275004 23498
rect 274404 -3342 274586 -3106
rect 274822 -3342 275004 -3106
rect 274404 -3426 275004 -3342
rect 274404 -3662 274586 -3426
rect 274822 -3662 275004 -3426
rect 274404 -3684 275004 -3662
rect 278004 135654 278604 171098
rect 278004 135418 278186 135654
rect 278422 135418 278604 135654
rect 278004 135334 278604 135418
rect 278004 135098 278186 135334
rect 278422 135098 278604 135334
rect 278004 99654 278604 135098
rect 278004 99418 278186 99654
rect 278422 99418 278604 99654
rect 278004 99334 278604 99418
rect 278004 99098 278186 99334
rect 278422 99098 278604 99334
rect 278004 63654 278604 99098
rect 278004 63418 278186 63654
rect 278422 63418 278604 63654
rect 278004 63334 278604 63418
rect 278004 63098 278186 63334
rect 278422 63098 278604 63334
rect 278004 27654 278604 63098
rect 278004 27418 278186 27654
rect 278422 27418 278604 27654
rect 278004 27334 278604 27418
rect 278004 27098 278186 27334
rect 278422 27098 278604 27334
rect 278004 -4946 278604 27098
rect 278004 -5182 278186 -4946
rect 278422 -5182 278604 -4946
rect 278004 -5266 278604 -5182
rect 278004 -5502 278186 -5266
rect 278422 -5502 278604 -5266
rect 278004 -5524 278604 -5502
rect 281604 499254 282204 534698
rect 288804 704838 289404 705780
rect 288804 704602 288986 704838
rect 289222 704602 289404 704838
rect 288804 704518 289404 704602
rect 288804 704282 288986 704518
rect 289222 704282 289404 704518
rect 288804 686454 289404 704282
rect 288804 686218 288986 686454
rect 289222 686218 289404 686454
rect 288804 686134 289404 686218
rect 288804 685898 288986 686134
rect 289222 685898 289404 686134
rect 288804 650454 289404 685898
rect 288804 650218 288986 650454
rect 289222 650218 289404 650454
rect 288804 650134 289404 650218
rect 288804 649898 288986 650134
rect 289222 649898 289404 650134
rect 288804 614454 289404 649898
rect 288804 614218 288986 614454
rect 289222 614218 289404 614454
rect 288804 614134 289404 614218
rect 288804 613898 288986 614134
rect 289222 613898 289404 614134
rect 288804 578454 289404 613898
rect 288804 578218 288986 578454
rect 289222 578218 289404 578454
rect 288804 578134 289404 578218
rect 288804 577898 288986 578134
rect 289222 577898 289404 578134
rect 288804 542454 289404 577898
rect 288804 542218 288986 542454
rect 289222 542218 289404 542454
rect 288804 542134 289404 542218
rect 288804 541898 288986 542134
rect 289222 541898 289404 542134
rect 284891 519348 284957 519349
rect 284891 519284 284892 519348
rect 284956 519284 284957 519348
rect 284891 519283 284957 519284
rect 284894 518669 284954 519283
rect 283051 518668 283117 518669
rect 283051 518604 283052 518668
rect 283116 518604 283117 518668
rect 283051 518603 283117 518604
rect 284891 518668 284957 518669
rect 284891 518604 284892 518668
rect 284956 518604 284957 518668
rect 284891 518603 284957 518604
rect 283054 517989 283114 518603
rect 282867 517988 282933 517989
rect 282867 517924 282868 517988
rect 282932 517924 282933 517988
rect 282867 517923 282933 517924
rect 283051 517988 283117 517989
rect 283051 517924 283052 517988
rect 283116 517924 283117 517988
rect 283051 517923 283117 517924
rect 282870 517850 282930 517923
rect 282870 517790 283334 517850
rect 281604 499018 281786 499254
rect 282022 499018 282204 499254
rect 281604 498934 282204 499018
rect 281604 498698 281786 498934
rect 282022 498698 282204 498934
rect 281604 463254 282204 498698
rect 281604 463018 281786 463254
rect 282022 463018 282204 463254
rect 281604 462934 282204 463018
rect 281604 462698 281786 462934
rect 282022 462698 282204 462934
rect 281604 427254 282204 462698
rect 281604 427018 281786 427254
rect 282022 427018 282204 427254
rect 281604 426934 282204 427018
rect 281604 426698 281786 426934
rect 282022 426698 282204 426934
rect 281604 391254 282204 426698
rect 281604 391018 281786 391254
rect 282022 391018 282204 391254
rect 281604 390934 282204 391018
rect 281604 390698 281786 390934
rect 282022 390698 282204 390934
rect 281604 355254 282204 390698
rect 281604 355018 281786 355254
rect 282022 355018 282204 355254
rect 281604 354934 282204 355018
rect 281604 354698 281786 354934
rect 282022 354698 282204 354934
rect 281604 319254 282204 354698
rect 281604 319018 281786 319254
rect 282022 319018 282204 319254
rect 281604 318934 282204 319018
rect 281604 318698 281786 318934
rect 282022 318698 282204 318934
rect 281604 283254 282204 318698
rect 281604 283018 281786 283254
rect 282022 283018 282204 283254
rect 281604 282934 282204 283018
rect 281604 282698 281786 282934
rect 282022 282698 282204 282934
rect 281604 247254 282204 282698
rect 281604 247018 281786 247254
rect 282022 247018 282204 247254
rect 281604 246934 282204 247018
rect 281604 246698 281786 246934
rect 282022 246698 282204 246934
rect 281604 211254 282204 246698
rect 281604 211018 281786 211254
rect 282022 211018 282204 211254
rect 281604 210934 282204 211018
rect 281604 210698 281786 210934
rect 282022 210698 282204 210934
rect 281604 175254 282204 210698
rect 281604 175018 281786 175254
rect 282022 175018 282204 175254
rect 281604 174934 282204 175018
rect 281604 174698 281786 174934
rect 282022 174698 282204 174934
rect 281604 139254 282204 174698
rect 281604 139018 281786 139254
rect 282022 139018 282204 139254
rect 281604 138934 282204 139018
rect 281604 138698 281786 138934
rect 282022 138698 282204 138934
rect 281604 103254 282204 138698
rect 288804 506454 289404 541898
rect 288804 506218 288986 506454
rect 289222 506218 289404 506454
rect 288804 506134 289404 506218
rect 288804 505898 288986 506134
rect 289222 505898 289404 506134
rect 288804 470454 289404 505898
rect 288804 470218 288986 470454
rect 289222 470218 289404 470454
rect 288804 470134 289404 470218
rect 288804 469898 288986 470134
rect 289222 469898 289404 470134
rect 288804 434454 289404 469898
rect 288804 434218 288986 434454
rect 289222 434218 289404 434454
rect 288804 434134 289404 434218
rect 288804 433898 288986 434134
rect 289222 433898 289404 434134
rect 288804 398454 289404 433898
rect 288804 398218 288986 398454
rect 289222 398218 289404 398454
rect 288804 398134 289404 398218
rect 288804 397898 288986 398134
rect 289222 397898 289404 398134
rect 288804 362454 289404 397898
rect 288804 362218 288986 362454
rect 289222 362218 289404 362454
rect 288804 362134 289404 362218
rect 288804 361898 288986 362134
rect 289222 361898 289404 362134
rect 288804 326454 289404 361898
rect 288804 326218 288986 326454
rect 289222 326218 289404 326454
rect 288804 326134 289404 326218
rect 288804 325898 288986 326134
rect 289222 325898 289404 326134
rect 288804 290454 289404 325898
rect 288804 290218 288986 290454
rect 289222 290218 289404 290454
rect 288804 290134 289404 290218
rect 288804 289898 288986 290134
rect 289222 289898 289404 290134
rect 288804 254454 289404 289898
rect 288804 254218 288986 254454
rect 289222 254218 289404 254454
rect 288804 254134 289404 254218
rect 288804 253898 288986 254134
rect 289222 253898 289404 254134
rect 288804 218454 289404 253898
rect 288804 218218 288986 218454
rect 289222 218218 289404 218454
rect 288804 218134 289404 218218
rect 288804 217898 288986 218134
rect 289222 217898 289404 218134
rect 288804 182454 289404 217898
rect 288804 182218 288986 182454
rect 289222 182218 289404 182454
rect 288804 182134 289404 182218
rect 288804 181898 288986 182134
rect 289222 181898 289404 182134
rect 288804 146454 289404 181898
rect 288804 146218 288986 146454
rect 289222 146218 289404 146454
rect 288804 146134 289404 146218
rect 288804 145898 288986 146134
rect 289222 145898 289404 146134
rect 283971 123996 284037 123997
rect 283971 123932 283972 123996
rect 284036 123932 284037 123996
rect 283971 123931 284037 123932
rect 283974 106317 284034 123931
rect 288804 110454 289404 145898
rect 288804 110218 288986 110454
rect 289222 110218 289404 110454
rect 288804 110134 289404 110218
rect 288804 109898 288986 110134
rect 289222 109898 289404 110134
rect 283971 106316 284037 106317
rect 283971 106252 283972 106316
rect 284036 106252 284037 106316
rect 283971 106251 284037 106252
rect 281604 103018 281786 103254
rect 282022 103018 282204 103254
rect 281604 102934 282204 103018
rect 281604 102698 281786 102934
rect 282022 102698 282204 102934
rect 281604 67254 282204 102698
rect 281604 67018 281786 67254
rect 282022 67018 282204 67254
rect 281604 66934 282204 67018
rect 281604 66698 281786 66934
rect 282022 66698 282204 66934
rect 281604 31254 282204 66698
rect 281604 31018 281786 31254
rect 282022 31018 282204 31254
rect 281604 30934 282204 31018
rect 281604 30698 281786 30934
rect 282022 30698 282204 30934
rect 263604 -6102 263786 -5866
rect 264022 -6102 264204 -5866
rect 263604 -6186 264204 -6102
rect 263604 -6422 263786 -6186
rect 264022 -6422 264204 -6186
rect 263604 -7364 264204 -6422
rect 281604 -6786 282204 30698
rect 288804 74454 289404 109898
rect 288804 74218 288986 74454
rect 289222 74218 289404 74454
rect 288804 74134 289404 74218
rect 288804 73898 288986 74134
rect 289222 73898 289404 74134
rect 288804 38454 289404 73898
rect 288804 38218 288986 38454
rect 289222 38218 289404 38454
rect 288804 38134 289404 38218
rect 288804 37898 288986 38134
rect 289222 37898 289404 38134
rect 288804 2454 289404 37898
rect 288804 2218 288986 2454
rect 289222 2218 289404 2454
rect 288804 2134 289404 2218
rect 288804 1898 288986 2134
rect 289222 1898 289404 2134
rect 288804 -346 289404 1898
rect 288804 -582 288986 -346
rect 289222 -582 289404 -346
rect 288804 -666 289404 -582
rect 288804 -902 288986 -666
rect 289222 -902 289404 -666
rect 288804 -1844 289404 -902
rect 292404 690054 293004 706122
rect 292404 689818 292586 690054
rect 292822 689818 293004 690054
rect 292404 689734 293004 689818
rect 292404 689498 292586 689734
rect 292822 689498 293004 689734
rect 292404 654054 293004 689498
rect 292404 653818 292586 654054
rect 292822 653818 293004 654054
rect 292404 653734 293004 653818
rect 292404 653498 292586 653734
rect 292822 653498 293004 653734
rect 292404 618054 293004 653498
rect 292404 617818 292586 618054
rect 292822 617818 293004 618054
rect 292404 617734 293004 617818
rect 292404 617498 292586 617734
rect 292822 617498 293004 617734
rect 292404 582054 293004 617498
rect 292404 581818 292586 582054
rect 292822 581818 293004 582054
rect 292404 581734 293004 581818
rect 292404 581498 292586 581734
rect 292822 581498 293004 581734
rect 292404 546054 293004 581498
rect 292404 545818 292586 546054
rect 292822 545818 293004 546054
rect 292404 545734 293004 545818
rect 292404 545498 292586 545734
rect 292822 545498 293004 545734
rect 292404 510054 293004 545498
rect 296004 693654 296604 707962
rect 296004 693418 296186 693654
rect 296422 693418 296604 693654
rect 296004 693334 296604 693418
rect 296004 693098 296186 693334
rect 296422 693098 296604 693334
rect 296004 657654 296604 693098
rect 296004 657418 296186 657654
rect 296422 657418 296604 657654
rect 296004 657334 296604 657418
rect 296004 657098 296186 657334
rect 296422 657098 296604 657334
rect 296004 621654 296604 657098
rect 296004 621418 296186 621654
rect 296422 621418 296604 621654
rect 296004 621334 296604 621418
rect 296004 621098 296186 621334
rect 296422 621098 296604 621334
rect 296004 585654 296604 621098
rect 296004 585418 296186 585654
rect 296422 585418 296604 585654
rect 296004 585334 296604 585418
rect 296004 585098 296186 585334
rect 296422 585098 296604 585334
rect 296004 549654 296604 585098
rect 296004 549418 296186 549654
rect 296422 549418 296604 549654
rect 296004 549334 296604 549418
rect 296004 549098 296186 549334
rect 296422 549098 296604 549334
rect 294459 519212 294525 519213
rect 294459 519148 294460 519212
rect 294524 519148 294525 519212
rect 294459 519147 294525 519148
rect 294275 518940 294341 518941
rect 294275 518876 294276 518940
rect 294340 518876 294341 518940
rect 294275 518875 294341 518876
rect 294278 518669 294338 518875
rect 294275 518668 294341 518669
rect 294275 518604 294276 518668
rect 294340 518604 294341 518668
rect 294275 518603 294341 518604
rect 294462 518261 294522 519147
rect 294643 518668 294709 518669
rect 294643 518604 294644 518668
rect 294708 518604 294709 518668
rect 294643 518603 294709 518604
rect 294459 518260 294525 518261
rect 294459 518196 294460 518260
rect 294524 518196 294525 518260
rect 294459 518195 294525 518196
rect 294646 517989 294706 518603
rect 294643 517988 294709 517989
rect 294643 517924 294644 517988
rect 294708 517924 294709 517988
rect 294643 517923 294709 517924
rect 292404 509818 292586 510054
rect 292822 509818 293004 510054
rect 292404 509734 293004 509818
rect 292404 509498 292586 509734
rect 292822 509498 293004 509734
rect 292404 474054 293004 509498
rect 292404 473818 292586 474054
rect 292822 473818 293004 474054
rect 292404 473734 293004 473818
rect 292404 473498 292586 473734
rect 292822 473498 293004 473734
rect 292404 438054 293004 473498
rect 292404 437818 292586 438054
rect 292822 437818 293004 438054
rect 292404 437734 293004 437818
rect 292404 437498 292586 437734
rect 292822 437498 293004 437734
rect 292404 402054 293004 437498
rect 292404 401818 292586 402054
rect 292822 401818 293004 402054
rect 292404 401734 293004 401818
rect 292404 401498 292586 401734
rect 292822 401498 293004 401734
rect 292404 366054 293004 401498
rect 292404 365818 292586 366054
rect 292822 365818 293004 366054
rect 292404 365734 293004 365818
rect 292404 365498 292586 365734
rect 292822 365498 293004 365734
rect 292404 330054 293004 365498
rect 292404 329818 292586 330054
rect 292822 329818 293004 330054
rect 292404 329734 293004 329818
rect 292404 329498 292586 329734
rect 292822 329498 293004 329734
rect 292404 294054 293004 329498
rect 292404 293818 292586 294054
rect 292822 293818 293004 294054
rect 292404 293734 293004 293818
rect 292404 293498 292586 293734
rect 292822 293498 293004 293734
rect 292404 258054 293004 293498
rect 292404 257818 292586 258054
rect 292822 257818 293004 258054
rect 292404 257734 293004 257818
rect 292404 257498 292586 257734
rect 292822 257498 293004 257734
rect 292404 222054 293004 257498
rect 292404 221818 292586 222054
rect 292822 221818 293004 222054
rect 292404 221734 293004 221818
rect 292404 221498 292586 221734
rect 292822 221498 293004 221734
rect 292404 186054 293004 221498
rect 292404 185818 292586 186054
rect 292822 185818 293004 186054
rect 292404 185734 293004 185818
rect 292404 185498 292586 185734
rect 292822 185498 293004 185734
rect 292404 150054 293004 185498
rect 292404 149818 292586 150054
rect 292822 149818 293004 150054
rect 292404 149734 293004 149818
rect 292404 149498 292586 149734
rect 292822 149498 293004 149734
rect 292404 114054 293004 149498
rect 292404 113818 292586 114054
rect 292822 113818 293004 114054
rect 292404 113734 293004 113818
rect 292404 113498 292586 113734
rect 292822 113498 293004 113734
rect 292404 78054 293004 113498
rect 292404 77818 292586 78054
rect 292822 77818 293004 78054
rect 292404 77734 293004 77818
rect 292404 77498 292586 77734
rect 292822 77498 293004 77734
rect 292404 42054 293004 77498
rect 292404 41818 292586 42054
rect 292822 41818 293004 42054
rect 292404 41734 293004 41818
rect 292404 41498 292586 41734
rect 292822 41498 293004 41734
rect 292404 6054 293004 41498
rect 292404 5818 292586 6054
rect 292822 5818 293004 6054
rect 292404 5734 293004 5818
rect 292404 5498 292586 5734
rect 292822 5498 293004 5734
rect 292404 -2186 293004 5498
rect 292404 -2422 292586 -2186
rect 292822 -2422 293004 -2186
rect 292404 -2506 293004 -2422
rect 292404 -2742 292586 -2506
rect 292822 -2742 293004 -2506
rect 292404 -3684 293004 -2742
rect 296004 513654 296604 549098
rect 299604 697254 300204 709802
rect 317604 711278 318204 711300
rect 317604 711042 317786 711278
rect 318022 711042 318204 711278
rect 317604 710958 318204 711042
rect 317604 710722 317786 710958
rect 318022 710722 318204 710958
rect 314004 709438 314604 709460
rect 314004 709202 314186 709438
rect 314422 709202 314604 709438
rect 314004 709118 314604 709202
rect 314004 708882 314186 709118
rect 314422 708882 314604 709118
rect 310404 707598 311004 707620
rect 310404 707362 310586 707598
rect 310822 707362 311004 707598
rect 310404 707278 311004 707362
rect 310404 707042 310586 707278
rect 310822 707042 311004 707278
rect 299604 697018 299786 697254
rect 300022 697018 300204 697254
rect 299604 696934 300204 697018
rect 299604 696698 299786 696934
rect 300022 696698 300204 696934
rect 299604 661254 300204 696698
rect 299604 661018 299786 661254
rect 300022 661018 300204 661254
rect 299604 660934 300204 661018
rect 299604 660698 299786 660934
rect 300022 660698 300204 660934
rect 299604 625254 300204 660698
rect 299604 625018 299786 625254
rect 300022 625018 300204 625254
rect 299604 624934 300204 625018
rect 299604 624698 299786 624934
rect 300022 624698 300204 624934
rect 299604 589254 300204 624698
rect 299604 589018 299786 589254
rect 300022 589018 300204 589254
rect 299604 588934 300204 589018
rect 299604 588698 299786 588934
rect 300022 588698 300204 588934
rect 299604 553254 300204 588698
rect 299604 553018 299786 553254
rect 300022 553018 300204 553254
rect 299604 552934 300204 553018
rect 299604 552698 299786 552934
rect 300022 552698 300204 552934
rect 299243 519212 299309 519213
rect 299243 519148 299244 519212
rect 299308 519148 299309 519212
rect 299243 519147 299309 519148
rect 298875 518940 298941 518941
rect 298875 518876 298876 518940
rect 298940 518876 298941 518940
rect 298875 518875 298941 518876
rect 298878 518669 298938 518875
rect 298691 518668 298757 518669
rect 298691 518604 298692 518668
rect 298756 518604 298757 518668
rect 298691 518603 298757 518604
rect 298875 518668 298941 518669
rect 298875 518604 298876 518668
rect 298940 518604 298941 518668
rect 298875 518603 298941 518604
rect 298694 518530 298754 518603
rect 298694 518470 298938 518530
rect 298878 517989 298938 518470
rect 299246 518261 299306 519147
rect 299059 518260 299125 518261
rect 299059 518196 299060 518260
rect 299124 518196 299125 518260
rect 299059 518195 299125 518196
rect 299243 518260 299309 518261
rect 299243 518196 299244 518260
rect 299308 518196 299309 518260
rect 299243 518195 299309 518196
rect 298875 517988 298941 517989
rect 298875 517924 298876 517988
rect 298940 517924 298941 517988
rect 298875 517923 298941 517924
rect 298507 517852 298573 517853
rect 298507 517788 298508 517852
rect 298572 517850 298573 517852
rect 298875 517852 298941 517853
rect 298875 517850 298876 517852
rect 298572 517790 298876 517850
rect 298572 517788 298573 517790
rect 298507 517787 298573 517788
rect 298875 517788 298876 517790
rect 298940 517788 298941 517852
rect 299062 517850 299122 518195
rect 299243 518124 299309 518125
rect 299243 518060 299244 518124
rect 299308 518060 299309 518124
rect 299243 518059 299309 518060
rect 299246 517850 299306 518059
rect 299062 517790 299306 517850
rect 298875 517787 298941 517788
rect 296004 513418 296186 513654
rect 296422 513418 296604 513654
rect 296004 513334 296604 513418
rect 296004 513098 296186 513334
rect 296422 513098 296604 513334
rect 296004 477654 296604 513098
rect 296004 477418 296186 477654
rect 296422 477418 296604 477654
rect 296004 477334 296604 477418
rect 296004 477098 296186 477334
rect 296422 477098 296604 477334
rect 296004 441654 296604 477098
rect 296004 441418 296186 441654
rect 296422 441418 296604 441654
rect 296004 441334 296604 441418
rect 296004 441098 296186 441334
rect 296422 441098 296604 441334
rect 296004 405654 296604 441098
rect 296004 405418 296186 405654
rect 296422 405418 296604 405654
rect 296004 405334 296604 405418
rect 296004 405098 296186 405334
rect 296422 405098 296604 405334
rect 296004 369654 296604 405098
rect 296004 369418 296186 369654
rect 296422 369418 296604 369654
rect 296004 369334 296604 369418
rect 296004 369098 296186 369334
rect 296422 369098 296604 369334
rect 296004 333654 296604 369098
rect 296004 333418 296186 333654
rect 296422 333418 296604 333654
rect 296004 333334 296604 333418
rect 296004 333098 296186 333334
rect 296422 333098 296604 333334
rect 296004 297654 296604 333098
rect 296004 297418 296186 297654
rect 296422 297418 296604 297654
rect 296004 297334 296604 297418
rect 296004 297098 296186 297334
rect 296422 297098 296604 297334
rect 296004 261654 296604 297098
rect 296004 261418 296186 261654
rect 296422 261418 296604 261654
rect 296004 261334 296604 261418
rect 296004 261098 296186 261334
rect 296422 261098 296604 261334
rect 296004 225654 296604 261098
rect 296004 225418 296186 225654
rect 296422 225418 296604 225654
rect 296004 225334 296604 225418
rect 296004 225098 296186 225334
rect 296422 225098 296604 225334
rect 296004 189654 296604 225098
rect 296004 189418 296186 189654
rect 296422 189418 296604 189654
rect 296004 189334 296604 189418
rect 296004 189098 296186 189334
rect 296422 189098 296604 189334
rect 296004 153654 296604 189098
rect 296004 153418 296186 153654
rect 296422 153418 296604 153654
rect 296004 153334 296604 153418
rect 296004 153098 296186 153334
rect 296422 153098 296604 153334
rect 296004 117654 296604 153098
rect 296004 117418 296186 117654
rect 296422 117418 296604 117654
rect 296004 117334 296604 117418
rect 296004 117098 296186 117334
rect 296422 117098 296604 117334
rect 296004 81654 296604 117098
rect 296004 81418 296186 81654
rect 296422 81418 296604 81654
rect 296004 81334 296604 81418
rect 296004 81098 296186 81334
rect 296422 81098 296604 81334
rect 296004 45654 296604 81098
rect 296004 45418 296186 45654
rect 296422 45418 296604 45654
rect 296004 45334 296604 45418
rect 296004 45098 296186 45334
rect 296422 45098 296604 45334
rect 296004 9654 296604 45098
rect 296004 9418 296186 9654
rect 296422 9418 296604 9654
rect 296004 9334 296604 9418
rect 296004 9098 296186 9334
rect 296422 9098 296604 9334
rect 296004 -4026 296604 9098
rect 296004 -4262 296186 -4026
rect 296422 -4262 296604 -4026
rect 296004 -4346 296604 -4262
rect 296004 -4582 296186 -4346
rect 296422 -4582 296604 -4346
rect 296004 -5524 296604 -4582
rect 299604 517254 300204 552698
rect 306804 705758 307404 705780
rect 306804 705522 306986 705758
rect 307222 705522 307404 705758
rect 306804 705438 307404 705522
rect 306804 705202 306986 705438
rect 307222 705202 307404 705438
rect 306804 668454 307404 705202
rect 306804 668218 306986 668454
rect 307222 668218 307404 668454
rect 306804 668134 307404 668218
rect 306804 667898 306986 668134
rect 307222 667898 307404 668134
rect 306804 632454 307404 667898
rect 306804 632218 306986 632454
rect 307222 632218 307404 632454
rect 306804 632134 307404 632218
rect 306804 631898 306986 632134
rect 307222 631898 307404 632134
rect 306804 596454 307404 631898
rect 306804 596218 306986 596454
rect 307222 596218 307404 596454
rect 306804 596134 307404 596218
rect 306804 595898 306986 596134
rect 307222 595898 307404 596134
rect 306804 560454 307404 595898
rect 306804 560218 306986 560454
rect 307222 560218 307404 560454
rect 306804 560134 307404 560218
rect 306804 559898 306986 560134
rect 307222 559898 307404 560134
rect 306804 524454 307404 559898
rect 306804 524218 306986 524454
rect 307222 524218 307404 524454
rect 306804 524134 307404 524218
rect 306804 523898 306986 524134
rect 307222 523898 307404 524134
rect 302739 518940 302805 518941
rect 302739 518876 302740 518940
rect 302804 518876 302805 518940
rect 302739 518875 302805 518876
rect 301819 518668 301885 518669
rect 301819 518604 301820 518668
rect 301884 518604 301885 518668
rect 301819 518603 301885 518604
rect 302003 518668 302069 518669
rect 302003 518604 302004 518668
rect 302068 518604 302069 518668
rect 302003 518603 302069 518604
rect 301822 517850 301882 518603
rect 302006 517989 302066 518603
rect 302003 517988 302069 517989
rect 302003 517924 302004 517988
rect 302068 517924 302069 517988
rect 302003 517923 302069 517924
rect 302187 517988 302253 517989
rect 302187 517924 302188 517988
rect 302252 517924 302253 517988
rect 302742 517938 302802 518875
rect 302187 517923 302253 517924
rect 302190 517850 302250 517923
rect 301822 517790 302250 517850
rect 299604 517018 299786 517254
rect 300022 517018 300204 517254
rect 299604 516934 300204 517018
rect 299604 516698 299786 516934
rect 300022 516698 300204 516934
rect 299604 481254 300204 516698
rect 299604 481018 299786 481254
rect 300022 481018 300204 481254
rect 299604 480934 300204 481018
rect 299604 480698 299786 480934
rect 300022 480698 300204 480934
rect 299604 445254 300204 480698
rect 299604 445018 299786 445254
rect 300022 445018 300204 445254
rect 299604 444934 300204 445018
rect 299604 444698 299786 444934
rect 300022 444698 300204 444934
rect 299604 409254 300204 444698
rect 299604 409018 299786 409254
rect 300022 409018 300204 409254
rect 299604 408934 300204 409018
rect 299604 408698 299786 408934
rect 300022 408698 300204 408934
rect 299604 373254 300204 408698
rect 299604 373018 299786 373254
rect 300022 373018 300204 373254
rect 299604 372934 300204 373018
rect 299604 372698 299786 372934
rect 300022 372698 300204 372934
rect 299604 337254 300204 372698
rect 299604 337018 299786 337254
rect 300022 337018 300204 337254
rect 299604 336934 300204 337018
rect 299604 336698 299786 336934
rect 300022 336698 300204 336934
rect 299604 301254 300204 336698
rect 299604 301018 299786 301254
rect 300022 301018 300204 301254
rect 299604 300934 300204 301018
rect 299604 300698 299786 300934
rect 300022 300698 300204 300934
rect 299604 265254 300204 300698
rect 299604 265018 299786 265254
rect 300022 265018 300204 265254
rect 299604 264934 300204 265018
rect 299604 264698 299786 264934
rect 300022 264698 300204 264934
rect 299604 229254 300204 264698
rect 299604 229018 299786 229254
rect 300022 229018 300204 229254
rect 299604 228934 300204 229018
rect 299604 228698 299786 228934
rect 300022 228698 300204 228934
rect 299604 193254 300204 228698
rect 299604 193018 299786 193254
rect 300022 193018 300204 193254
rect 299604 192934 300204 193018
rect 299604 192698 299786 192934
rect 300022 192698 300204 192934
rect 299604 157254 300204 192698
rect 299604 157018 299786 157254
rect 300022 157018 300204 157254
rect 299604 156934 300204 157018
rect 299604 156698 299786 156934
rect 300022 156698 300204 156934
rect 299604 121254 300204 156698
rect 299604 121018 299786 121254
rect 300022 121018 300204 121254
rect 299604 120934 300204 121018
rect 299604 120698 299786 120934
rect 300022 120698 300204 120934
rect 299604 85254 300204 120698
rect 299604 85018 299786 85254
rect 300022 85018 300204 85254
rect 299604 84934 300204 85018
rect 299604 84698 299786 84934
rect 300022 84698 300204 84934
rect 299604 49254 300204 84698
rect 299604 49018 299786 49254
rect 300022 49018 300204 49254
rect 299604 48934 300204 49018
rect 299604 48698 299786 48934
rect 300022 48698 300204 48934
rect 299604 13254 300204 48698
rect 299604 13018 299786 13254
rect 300022 13018 300204 13254
rect 299604 12934 300204 13018
rect 299604 12698 299786 12934
rect 300022 12698 300204 12934
rect 281604 -7022 281786 -6786
rect 282022 -7022 282204 -6786
rect 281604 -7106 282204 -7022
rect 281604 -7342 281786 -7106
rect 282022 -7342 282204 -7106
rect 281604 -7364 282204 -7342
rect 299604 -5866 300204 12698
rect 306804 488454 307404 523898
rect 310404 672054 311004 707042
rect 310404 671818 310586 672054
rect 310822 671818 311004 672054
rect 310404 671734 311004 671818
rect 310404 671498 310586 671734
rect 310822 671498 311004 671734
rect 310404 636054 311004 671498
rect 310404 635818 310586 636054
rect 310822 635818 311004 636054
rect 310404 635734 311004 635818
rect 310404 635498 310586 635734
rect 310822 635498 311004 635734
rect 310404 600054 311004 635498
rect 310404 599818 310586 600054
rect 310822 599818 311004 600054
rect 310404 599734 311004 599818
rect 310404 599498 310586 599734
rect 310822 599498 311004 599734
rect 310404 564054 311004 599498
rect 310404 563818 310586 564054
rect 310822 563818 311004 564054
rect 310404 563734 311004 563818
rect 310404 563498 310586 563734
rect 310822 563498 311004 563734
rect 310404 528054 311004 563498
rect 310404 527818 310586 528054
rect 310822 527818 311004 528054
rect 310404 527734 311004 527818
rect 310404 527498 310586 527734
rect 310822 527498 311004 527734
rect 309363 519484 309429 519485
rect 309363 519420 309364 519484
rect 309428 519420 309429 519484
rect 309363 519419 309429 519420
rect 309179 518668 309245 518669
rect 309179 518604 309180 518668
rect 309244 518604 309245 518668
rect 309179 518603 309245 518604
rect 309182 518530 309242 518603
rect 309366 518530 309426 519419
rect 309182 518470 309426 518530
rect 306804 488218 306986 488454
rect 307222 488218 307404 488454
rect 306804 488134 307404 488218
rect 306804 487898 306986 488134
rect 307222 487898 307404 488134
rect 306804 452454 307404 487898
rect 306804 452218 306986 452454
rect 307222 452218 307404 452454
rect 306804 452134 307404 452218
rect 306804 451898 306986 452134
rect 307222 451898 307404 452134
rect 306804 416454 307404 451898
rect 306804 416218 306986 416454
rect 307222 416218 307404 416454
rect 306804 416134 307404 416218
rect 306804 415898 306986 416134
rect 307222 415898 307404 416134
rect 306804 380454 307404 415898
rect 306804 380218 306986 380454
rect 307222 380218 307404 380454
rect 306804 380134 307404 380218
rect 306804 379898 306986 380134
rect 307222 379898 307404 380134
rect 306804 344454 307404 379898
rect 306804 344218 306986 344454
rect 307222 344218 307404 344454
rect 306804 344134 307404 344218
rect 306804 343898 306986 344134
rect 307222 343898 307404 344134
rect 306804 308454 307404 343898
rect 306804 308218 306986 308454
rect 307222 308218 307404 308454
rect 306804 308134 307404 308218
rect 306804 307898 306986 308134
rect 307222 307898 307404 308134
rect 306804 272454 307404 307898
rect 306804 272218 306986 272454
rect 307222 272218 307404 272454
rect 306804 272134 307404 272218
rect 306804 271898 306986 272134
rect 307222 271898 307404 272134
rect 306804 236454 307404 271898
rect 306804 236218 306986 236454
rect 307222 236218 307404 236454
rect 306804 236134 307404 236218
rect 306804 235898 306986 236134
rect 307222 235898 307404 236134
rect 306804 200454 307404 235898
rect 306804 200218 306986 200454
rect 307222 200218 307404 200454
rect 306804 200134 307404 200218
rect 306804 199898 306986 200134
rect 307222 199898 307404 200134
rect 306804 164454 307404 199898
rect 306804 164218 306986 164454
rect 307222 164218 307404 164454
rect 306804 164134 307404 164218
rect 306804 163898 306986 164134
rect 307222 163898 307404 164134
rect 306804 128454 307404 163898
rect 306804 128218 306986 128454
rect 307222 128218 307404 128454
rect 306804 128134 307404 128218
rect 306804 127898 306986 128134
rect 307222 127898 307404 128134
rect 306804 92454 307404 127898
rect 306804 92218 306986 92454
rect 307222 92218 307404 92454
rect 306804 92134 307404 92218
rect 306804 91898 306986 92134
rect 307222 91898 307404 92134
rect 306804 56454 307404 91898
rect 306804 56218 306986 56454
rect 307222 56218 307404 56454
rect 306804 56134 307404 56218
rect 306804 55898 306986 56134
rect 307222 55898 307404 56134
rect 306804 20454 307404 55898
rect 310404 492054 311004 527498
rect 314004 675654 314604 708882
rect 314004 675418 314186 675654
rect 314422 675418 314604 675654
rect 314004 675334 314604 675418
rect 314004 675098 314186 675334
rect 314422 675098 314604 675334
rect 314004 639654 314604 675098
rect 314004 639418 314186 639654
rect 314422 639418 314604 639654
rect 314004 639334 314604 639418
rect 314004 639098 314186 639334
rect 314422 639098 314604 639334
rect 314004 603654 314604 639098
rect 314004 603418 314186 603654
rect 314422 603418 314604 603654
rect 314004 603334 314604 603418
rect 314004 603098 314186 603334
rect 314422 603098 314604 603334
rect 314004 567654 314604 603098
rect 314004 567418 314186 567654
rect 314422 567418 314604 567654
rect 314004 567334 314604 567418
rect 314004 567098 314186 567334
rect 314422 567098 314604 567334
rect 314004 531654 314604 567098
rect 314004 531418 314186 531654
rect 314422 531418 314604 531654
rect 314004 531334 314604 531418
rect 314004 531098 314186 531334
rect 314422 531098 314604 531334
rect 313227 519484 313293 519485
rect 313227 519420 313228 519484
rect 313292 519420 313293 519484
rect 313227 519419 313293 519420
rect 312675 519348 312741 519349
rect 312675 519284 312676 519348
rect 312740 519284 312741 519348
rect 312675 519283 312741 519284
rect 312678 518941 312738 519283
rect 313230 519213 313290 519419
rect 313227 519212 313293 519213
rect 313227 519148 313228 519212
rect 313292 519148 313293 519212
rect 313227 519147 313293 519148
rect 312675 518940 312741 518941
rect 312675 518876 312676 518940
rect 312740 518876 312741 518940
rect 312675 518875 312741 518876
rect 310404 491818 310586 492054
rect 310822 491818 311004 492054
rect 310404 491734 311004 491818
rect 310404 491498 310586 491734
rect 310822 491498 311004 491734
rect 310404 456054 311004 491498
rect 310404 455818 310586 456054
rect 310822 455818 311004 456054
rect 310404 455734 311004 455818
rect 310404 455498 310586 455734
rect 310822 455498 311004 455734
rect 310404 420054 311004 455498
rect 310404 419818 310586 420054
rect 310822 419818 311004 420054
rect 310404 419734 311004 419818
rect 310404 419498 310586 419734
rect 310822 419498 311004 419734
rect 310404 384054 311004 419498
rect 310404 383818 310586 384054
rect 310822 383818 311004 384054
rect 310404 383734 311004 383818
rect 310404 383498 310586 383734
rect 310822 383498 311004 383734
rect 310404 348054 311004 383498
rect 310404 347818 310586 348054
rect 310822 347818 311004 348054
rect 310404 347734 311004 347818
rect 310404 347498 310586 347734
rect 310822 347498 311004 347734
rect 310404 312054 311004 347498
rect 310404 311818 310586 312054
rect 310822 311818 311004 312054
rect 310404 311734 311004 311818
rect 310404 311498 310586 311734
rect 310822 311498 311004 311734
rect 310404 276054 311004 311498
rect 310404 275818 310586 276054
rect 310822 275818 311004 276054
rect 310404 275734 311004 275818
rect 310404 275498 310586 275734
rect 310822 275498 311004 275734
rect 310404 240054 311004 275498
rect 310404 239818 310586 240054
rect 310822 239818 311004 240054
rect 310404 239734 311004 239818
rect 310404 239498 310586 239734
rect 310822 239498 311004 239734
rect 310404 204054 311004 239498
rect 310404 203818 310586 204054
rect 310822 203818 311004 204054
rect 310404 203734 311004 203818
rect 310404 203498 310586 203734
rect 310822 203498 311004 203734
rect 310404 168054 311004 203498
rect 310404 167818 310586 168054
rect 310822 167818 311004 168054
rect 310404 167734 311004 167818
rect 310404 167498 310586 167734
rect 310822 167498 311004 167734
rect 310404 132054 311004 167498
rect 310404 131818 310586 132054
rect 310822 131818 311004 132054
rect 310404 131734 311004 131818
rect 310404 131498 310586 131734
rect 310822 131498 311004 131734
rect 310404 96054 311004 131498
rect 310404 95818 310586 96054
rect 310822 95818 311004 96054
rect 310404 95734 311004 95818
rect 310404 95498 310586 95734
rect 310822 95498 311004 95734
rect 310404 60054 311004 95498
rect 310404 59818 310586 60054
rect 310822 59818 311004 60054
rect 310404 59734 311004 59818
rect 310404 59498 310586 59734
rect 310822 59498 311004 59734
rect 307707 40492 307773 40493
rect 307707 40428 307708 40492
rect 307772 40428 307773 40492
rect 307707 40427 307773 40428
rect 307710 40221 307770 40427
rect 307707 40220 307773 40221
rect 307707 40156 307708 40220
rect 307772 40156 307773 40220
rect 307707 40155 307773 40156
rect 306804 20218 306986 20454
rect 307222 20218 307404 20454
rect 306804 20134 307404 20218
rect 306804 19898 306986 20134
rect 307222 19898 307404 20134
rect 306804 -1266 307404 19898
rect 306804 -1502 306986 -1266
rect 307222 -1502 307404 -1266
rect 306804 -1586 307404 -1502
rect 306804 -1822 306986 -1586
rect 307222 -1822 307404 -1586
rect 306804 -1844 307404 -1822
rect 310404 24054 311004 59498
rect 310404 23818 310586 24054
rect 310822 23818 311004 24054
rect 310404 23734 311004 23818
rect 310404 23498 310586 23734
rect 310822 23498 311004 23734
rect 310404 -3106 311004 23498
rect 310404 -3342 310586 -3106
rect 310822 -3342 311004 -3106
rect 310404 -3426 311004 -3342
rect 310404 -3662 310586 -3426
rect 310822 -3662 311004 -3426
rect 310404 -3684 311004 -3662
rect 314004 495654 314604 531098
rect 314004 495418 314186 495654
rect 314422 495418 314604 495654
rect 314004 495334 314604 495418
rect 314004 495098 314186 495334
rect 314422 495098 314604 495334
rect 314004 459654 314604 495098
rect 314004 459418 314186 459654
rect 314422 459418 314604 459654
rect 314004 459334 314604 459418
rect 314004 459098 314186 459334
rect 314422 459098 314604 459334
rect 314004 423654 314604 459098
rect 314004 423418 314186 423654
rect 314422 423418 314604 423654
rect 314004 423334 314604 423418
rect 314004 423098 314186 423334
rect 314422 423098 314604 423334
rect 314004 387654 314604 423098
rect 314004 387418 314186 387654
rect 314422 387418 314604 387654
rect 314004 387334 314604 387418
rect 314004 387098 314186 387334
rect 314422 387098 314604 387334
rect 314004 351654 314604 387098
rect 314004 351418 314186 351654
rect 314422 351418 314604 351654
rect 314004 351334 314604 351418
rect 314004 351098 314186 351334
rect 314422 351098 314604 351334
rect 314004 315654 314604 351098
rect 314004 315418 314186 315654
rect 314422 315418 314604 315654
rect 314004 315334 314604 315418
rect 314004 315098 314186 315334
rect 314422 315098 314604 315334
rect 314004 279654 314604 315098
rect 314004 279418 314186 279654
rect 314422 279418 314604 279654
rect 314004 279334 314604 279418
rect 314004 279098 314186 279334
rect 314422 279098 314604 279334
rect 314004 243654 314604 279098
rect 314004 243418 314186 243654
rect 314422 243418 314604 243654
rect 314004 243334 314604 243418
rect 314004 243098 314186 243334
rect 314422 243098 314604 243334
rect 314004 207654 314604 243098
rect 314004 207418 314186 207654
rect 314422 207418 314604 207654
rect 314004 207334 314604 207418
rect 314004 207098 314186 207334
rect 314422 207098 314604 207334
rect 314004 171654 314604 207098
rect 314004 171418 314186 171654
rect 314422 171418 314604 171654
rect 314004 171334 314604 171418
rect 314004 171098 314186 171334
rect 314422 171098 314604 171334
rect 314004 135654 314604 171098
rect 314004 135418 314186 135654
rect 314422 135418 314604 135654
rect 314004 135334 314604 135418
rect 314004 135098 314186 135334
rect 314422 135098 314604 135334
rect 314004 99654 314604 135098
rect 314004 99418 314186 99654
rect 314422 99418 314604 99654
rect 314004 99334 314604 99418
rect 314004 99098 314186 99334
rect 314422 99098 314604 99334
rect 314004 63654 314604 99098
rect 314004 63418 314186 63654
rect 314422 63418 314604 63654
rect 314004 63334 314604 63418
rect 314004 63098 314186 63334
rect 314422 63098 314604 63334
rect 314004 27654 314604 63098
rect 314004 27418 314186 27654
rect 314422 27418 314604 27654
rect 314004 27334 314604 27418
rect 314004 27098 314186 27334
rect 314422 27098 314604 27334
rect 314004 -4946 314604 27098
rect 314004 -5182 314186 -4946
rect 314422 -5182 314604 -4946
rect 314004 -5266 314604 -5182
rect 314004 -5502 314186 -5266
rect 314422 -5502 314604 -5266
rect 314004 -5524 314604 -5502
rect 317604 679254 318204 710722
rect 335604 710358 336204 711300
rect 335604 710122 335786 710358
rect 336022 710122 336204 710358
rect 335604 710038 336204 710122
rect 335604 709802 335786 710038
rect 336022 709802 336204 710038
rect 332004 708518 332604 709460
rect 332004 708282 332186 708518
rect 332422 708282 332604 708518
rect 332004 708198 332604 708282
rect 332004 707962 332186 708198
rect 332422 707962 332604 708198
rect 328404 706678 329004 707620
rect 328404 706442 328586 706678
rect 328822 706442 329004 706678
rect 328404 706358 329004 706442
rect 328404 706122 328586 706358
rect 328822 706122 329004 706358
rect 317604 679018 317786 679254
rect 318022 679018 318204 679254
rect 317604 678934 318204 679018
rect 317604 678698 317786 678934
rect 318022 678698 318204 678934
rect 317604 643254 318204 678698
rect 317604 643018 317786 643254
rect 318022 643018 318204 643254
rect 317604 642934 318204 643018
rect 317604 642698 317786 642934
rect 318022 642698 318204 642934
rect 317604 607254 318204 642698
rect 317604 607018 317786 607254
rect 318022 607018 318204 607254
rect 317604 606934 318204 607018
rect 317604 606698 317786 606934
rect 318022 606698 318204 606934
rect 317604 571254 318204 606698
rect 317604 571018 317786 571254
rect 318022 571018 318204 571254
rect 317604 570934 318204 571018
rect 317604 570698 317786 570934
rect 318022 570698 318204 570934
rect 317604 535254 318204 570698
rect 317604 535018 317786 535254
rect 318022 535018 318204 535254
rect 317604 534934 318204 535018
rect 317604 534698 317786 534934
rect 318022 534698 318204 534934
rect 317604 499254 318204 534698
rect 324804 704838 325404 705780
rect 324804 704602 324986 704838
rect 325222 704602 325404 704838
rect 324804 704518 325404 704602
rect 324804 704282 324986 704518
rect 325222 704282 325404 704518
rect 324804 686454 325404 704282
rect 324804 686218 324986 686454
rect 325222 686218 325404 686454
rect 324804 686134 325404 686218
rect 324804 685898 324986 686134
rect 325222 685898 325404 686134
rect 324804 650454 325404 685898
rect 324804 650218 324986 650454
rect 325222 650218 325404 650454
rect 324804 650134 325404 650218
rect 324804 649898 324986 650134
rect 325222 649898 325404 650134
rect 324804 614454 325404 649898
rect 324804 614218 324986 614454
rect 325222 614218 325404 614454
rect 324804 614134 325404 614218
rect 324804 613898 324986 614134
rect 325222 613898 325404 614134
rect 324804 578454 325404 613898
rect 324804 578218 324986 578454
rect 325222 578218 325404 578454
rect 324804 578134 325404 578218
rect 324804 577898 324986 578134
rect 325222 577898 325404 578134
rect 324804 542454 325404 577898
rect 324804 542218 324986 542454
rect 325222 542218 325404 542454
rect 324804 542134 325404 542218
rect 324804 541898 324986 542134
rect 325222 541898 325404 542134
rect 322795 519212 322861 519213
rect 322795 519148 322796 519212
rect 322860 519148 322861 519212
rect 322795 519147 322861 519148
rect 321691 518804 321757 518805
rect 321691 518740 321692 518804
rect 321756 518740 321757 518804
rect 321691 518739 321757 518740
rect 321507 518668 321573 518669
rect 321507 518604 321508 518668
rect 321572 518604 321573 518668
rect 321507 518603 321573 518604
rect 321510 518530 321570 518603
rect 321694 518530 321754 518739
rect 322798 518669 322858 519147
rect 322795 518668 322861 518669
rect 322795 518604 322796 518668
rect 322860 518604 322861 518668
rect 322795 518603 322861 518604
rect 321510 518470 321754 518530
rect 317604 499018 317786 499254
rect 318022 499018 318204 499254
rect 317604 498934 318204 499018
rect 317604 498698 317786 498934
rect 318022 498698 318204 498934
rect 317604 463254 318204 498698
rect 317604 463018 317786 463254
rect 318022 463018 318204 463254
rect 317604 462934 318204 463018
rect 317604 462698 317786 462934
rect 318022 462698 318204 462934
rect 317604 427254 318204 462698
rect 317604 427018 317786 427254
rect 318022 427018 318204 427254
rect 317604 426934 318204 427018
rect 317604 426698 317786 426934
rect 318022 426698 318204 426934
rect 317604 391254 318204 426698
rect 317604 391018 317786 391254
rect 318022 391018 318204 391254
rect 317604 390934 318204 391018
rect 317604 390698 317786 390934
rect 318022 390698 318204 390934
rect 317604 355254 318204 390698
rect 317604 355018 317786 355254
rect 318022 355018 318204 355254
rect 317604 354934 318204 355018
rect 317604 354698 317786 354934
rect 318022 354698 318204 354934
rect 317604 319254 318204 354698
rect 317604 319018 317786 319254
rect 318022 319018 318204 319254
rect 317604 318934 318204 319018
rect 317604 318698 317786 318934
rect 318022 318698 318204 318934
rect 317604 283254 318204 318698
rect 317604 283018 317786 283254
rect 318022 283018 318204 283254
rect 317604 282934 318204 283018
rect 317604 282698 317786 282934
rect 318022 282698 318204 282934
rect 317604 247254 318204 282698
rect 317604 247018 317786 247254
rect 318022 247018 318204 247254
rect 317604 246934 318204 247018
rect 317604 246698 317786 246934
rect 318022 246698 318204 246934
rect 317604 211254 318204 246698
rect 317604 211018 317786 211254
rect 318022 211018 318204 211254
rect 317604 210934 318204 211018
rect 317604 210698 317786 210934
rect 318022 210698 318204 210934
rect 317604 175254 318204 210698
rect 317604 175018 317786 175254
rect 318022 175018 318204 175254
rect 317604 174934 318204 175018
rect 317604 174698 317786 174934
rect 318022 174698 318204 174934
rect 317604 139254 318204 174698
rect 324804 506454 325404 541898
rect 324804 506218 324986 506454
rect 325222 506218 325404 506454
rect 324804 506134 325404 506218
rect 324804 505898 324986 506134
rect 325222 505898 325404 506134
rect 324804 470454 325404 505898
rect 324804 470218 324986 470454
rect 325222 470218 325404 470454
rect 324804 470134 325404 470218
rect 324804 469898 324986 470134
rect 325222 469898 325404 470134
rect 324804 434454 325404 469898
rect 324804 434218 324986 434454
rect 325222 434218 325404 434454
rect 324804 434134 325404 434218
rect 324804 433898 324986 434134
rect 325222 433898 325404 434134
rect 324804 398454 325404 433898
rect 324804 398218 324986 398454
rect 325222 398218 325404 398454
rect 324804 398134 325404 398218
rect 324804 397898 324986 398134
rect 325222 397898 325404 398134
rect 324804 362454 325404 397898
rect 324804 362218 324986 362454
rect 325222 362218 325404 362454
rect 324804 362134 325404 362218
rect 324804 361898 324986 362134
rect 325222 361898 325404 362134
rect 324804 326454 325404 361898
rect 324804 326218 324986 326454
rect 325222 326218 325404 326454
rect 324804 326134 325404 326218
rect 324804 325898 324986 326134
rect 325222 325898 325404 326134
rect 324804 290454 325404 325898
rect 324804 290218 324986 290454
rect 325222 290218 325404 290454
rect 324804 290134 325404 290218
rect 324804 289898 324986 290134
rect 325222 289898 325404 290134
rect 324804 254454 325404 289898
rect 324804 254218 324986 254454
rect 325222 254218 325404 254454
rect 324804 254134 325404 254218
rect 324804 253898 324986 254134
rect 325222 253898 325404 254134
rect 324804 218454 325404 253898
rect 324804 218218 324986 218454
rect 325222 218218 325404 218454
rect 324804 218134 325404 218218
rect 324804 217898 324986 218134
rect 325222 217898 325404 218134
rect 324804 182454 325404 217898
rect 324804 182218 324986 182454
rect 325222 182218 325404 182454
rect 324804 182134 325404 182218
rect 324804 181898 324986 182134
rect 325222 181898 325404 182134
rect 318563 147796 318629 147797
rect 318563 147732 318564 147796
rect 318628 147732 318629 147796
rect 318563 147731 318629 147732
rect 318566 143581 318626 147731
rect 324804 146454 325404 181898
rect 324804 146218 324986 146454
rect 325222 146218 325404 146454
rect 324804 146134 325404 146218
rect 324804 145898 324986 146134
rect 325222 145898 325404 146134
rect 318563 143580 318629 143581
rect 318563 143516 318564 143580
rect 318628 143516 318629 143580
rect 318563 143515 318629 143516
rect 317604 139018 317786 139254
rect 318022 139018 318204 139254
rect 317604 138934 318204 139018
rect 317604 138698 317786 138934
rect 318022 138698 318204 138934
rect 317604 103254 318204 138698
rect 317604 103018 317786 103254
rect 318022 103018 318204 103254
rect 317604 102934 318204 103018
rect 317604 102698 317786 102934
rect 318022 102698 318204 102934
rect 317604 67254 318204 102698
rect 317604 67018 317786 67254
rect 318022 67018 318204 67254
rect 317604 66934 318204 67018
rect 317604 66698 317786 66934
rect 318022 66698 318204 66934
rect 317604 31254 318204 66698
rect 317604 31018 317786 31254
rect 318022 31018 318204 31254
rect 317604 30934 318204 31018
rect 317604 30698 317786 30934
rect 318022 30698 318204 30934
rect 299604 -6102 299786 -5866
rect 300022 -6102 300204 -5866
rect 299604 -6186 300204 -6102
rect 299604 -6422 299786 -6186
rect 300022 -6422 300204 -6186
rect 299604 -7364 300204 -6422
rect 317604 -6786 318204 30698
rect 324804 110454 325404 145898
rect 324804 110218 324986 110454
rect 325222 110218 325404 110454
rect 324804 110134 325404 110218
rect 324804 109898 324986 110134
rect 325222 109898 325404 110134
rect 324804 74454 325404 109898
rect 324804 74218 324986 74454
rect 325222 74218 325404 74454
rect 324804 74134 325404 74218
rect 324804 73898 324986 74134
rect 325222 73898 325404 74134
rect 324804 38454 325404 73898
rect 328404 690054 329004 706122
rect 328404 689818 328586 690054
rect 328822 689818 329004 690054
rect 328404 689734 329004 689818
rect 328404 689498 328586 689734
rect 328822 689498 329004 689734
rect 328404 654054 329004 689498
rect 328404 653818 328586 654054
rect 328822 653818 329004 654054
rect 328404 653734 329004 653818
rect 328404 653498 328586 653734
rect 328822 653498 329004 653734
rect 328404 618054 329004 653498
rect 328404 617818 328586 618054
rect 328822 617818 329004 618054
rect 328404 617734 329004 617818
rect 328404 617498 328586 617734
rect 328822 617498 329004 617734
rect 328404 582054 329004 617498
rect 328404 581818 328586 582054
rect 328822 581818 329004 582054
rect 328404 581734 329004 581818
rect 328404 581498 328586 581734
rect 328822 581498 329004 581734
rect 328404 546054 329004 581498
rect 328404 545818 328586 546054
rect 328822 545818 329004 546054
rect 328404 545734 329004 545818
rect 328404 545498 328586 545734
rect 328822 545498 329004 545734
rect 328404 510054 329004 545498
rect 328404 509818 328586 510054
rect 328822 509818 329004 510054
rect 328404 509734 329004 509818
rect 328404 509498 328586 509734
rect 328822 509498 329004 509734
rect 328404 474054 329004 509498
rect 328404 473818 328586 474054
rect 328822 473818 329004 474054
rect 328404 473734 329004 473818
rect 328404 473498 328586 473734
rect 328822 473498 329004 473734
rect 328404 438054 329004 473498
rect 328404 437818 328586 438054
rect 328822 437818 329004 438054
rect 328404 437734 329004 437818
rect 328404 437498 328586 437734
rect 328822 437498 329004 437734
rect 328404 402054 329004 437498
rect 328404 401818 328586 402054
rect 328822 401818 329004 402054
rect 328404 401734 329004 401818
rect 328404 401498 328586 401734
rect 328822 401498 329004 401734
rect 328404 366054 329004 401498
rect 328404 365818 328586 366054
rect 328822 365818 329004 366054
rect 328404 365734 329004 365818
rect 328404 365498 328586 365734
rect 328822 365498 329004 365734
rect 328404 330054 329004 365498
rect 328404 329818 328586 330054
rect 328822 329818 329004 330054
rect 328404 329734 329004 329818
rect 328404 329498 328586 329734
rect 328822 329498 329004 329734
rect 328404 294054 329004 329498
rect 328404 293818 328586 294054
rect 328822 293818 329004 294054
rect 328404 293734 329004 293818
rect 328404 293498 328586 293734
rect 328822 293498 329004 293734
rect 328404 258054 329004 293498
rect 328404 257818 328586 258054
rect 328822 257818 329004 258054
rect 328404 257734 329004 257818
rect 328404 257498 328586 257734
rect 328822 257498 329004 257734
rect 328404 222054 329004 257498
rect 328404 221818 328586 222054
rect 328822 221818 329004 222054
rect 328404 221734 329004 221818
rect 328404 221498 328586 221734
rect 328822 221498 329004 221734
rect 328404 186054 329004 221498
rect 328404 185818 328586 186054
rect 328822 185818 329004 186054
rect 328404 185734 329004 185818
rect 328404 185498 328586 185734
rect 328822 185498 329004 185734
rect 328404 150054 329004 185498
rect 328404 149818 328586 150054
rect 328822 149818 329004 150054
rect 328404 149734 329004 149818
rect 328404 149498 328586 149734
rect 328822 149498 329004 149734
rect 328404 114054 329004 149498
rect 332004 693654 332604 707962
rect 332004 693418 332186 693654
rect 332422 693418 332604 693654
rect 332004 693334 332604 693418
rect 332004 693098 332186 693334
rect 332422 693098 332604 693334
rect 332004 657654 332604 693098
rect 332004 657418 332186 657654
rect 332422 657418 332604 657654
rect 332004 657334 332604 657418
rect 332004 657098 332186 657334
rect 332422 657098 332604 657334
rect 332004 621654 332604 657098
rect 332004 621418 332186 621654
rect 332422 621418 332604 621654
rect 332004 621334 332604 621418
rect 332004 621098 332186 621334
rect 332422 621098 332604 621334
rect 332004 585654 332604 621098
rect 332004 585418 332186 585654
rect 332422 585418 332604 585654
rect 332004 585334 332604 585418
rect 332004 585098 332186 585334
rect 332422 585098 332604 585334
rect 332004 549654 332604 585098
rect 332004 549418 332186 549654
rect 332422 549418 332604 549654
rect 332004 549334 332604 549418
rect 332004 549098 332186 549334
rect 332422 549098 332604 549334
rect 332004 513654 332604 549098
rect 335604 697254 336204 709802
rect 353604 711278 354204 711300
rect 353604 711042 353786 711278
rect 354022 711042 354204 711278
rect 353604 710958 354204 711042
rect 353604 710722 353786 710958
rect 354022 710722 354204 710958
rect 350004 709438 350604 709460
rect 350004 709202 350186 709438
rect 350422 709202 350604 709438
rect 350004 709118 350604 709202
rect 350004 708882 350186 709118
rect 350422 708882 350604 709118
rect 346404 707598 347004 707620
rect 346404 707362 346586 707598
rect 346822 707362 347004 707598
rect 346404 707278 347004 707362
rect 346404 707042 346586 707278
rect 346822 707042 347004 707278
rect 335604 697018 335786 697254
rect 336022 697018 336204 697254
rect 335604 696934 336204 697018
rect 335604 696698 335786 696934
rect 336022 696698 336204 696934
rect 335604 661254 336204 696698
rect 335604 661018 335786 661254
rect 336022 661018 336204 661254
rect 335604 660934 336204 661018
rect 335604 660698 335786 660934
rect 336022 660698 336204 660934
rect 335604 625254 336204 660698
rect 335604 625018 335786 625254
rect 336022 625018 336204 625254
rect 335604 624934 336204 625018
rect 335604 624698 335786 624934
rect 336022 624698 336204 624934
rect 335604 589254 336204 624698
rect 335604 589018 335786 589254
rect 336022 589018 336204 589254
rect 335604 588934 336204 589018
rect 335604 588698 335786 588934
rect 336022 588698 336204 588934
rect 335604 553254 336204 588698
rect 335604 553018 335786 553254
rect 336022 553018 336204 553254
rect 335604 552934 336204 553018
rect 335604 552698 335786 552934
rect 336022 552698 336204 552934
rect 335307 518804 335373 518805
rect 335307 518740 335308 518804
rect 335372 518740 335373 518804
rect 335307 518739 335373 518740
rect 335310 517938 335370 518739
rect 332004 513418 332186 513654
rect 332422 513418 332604 513654
rect 332004 513334 332604 513418
rect 332004 513098 332186 513334
rect 332422 513098 332604 513334
rect 332004 477654 332604 513098
rect 332004 477418 332186 477654
rect 332422 477418 332604 477654
rect 332004 477334 332604 477418
rect 332004 477098 332186 477334
rect 332422 477098 332604 477334
rect 332004 441654 332604 477098
rect 332004 441418 332186 441654
rect 332422 441418 332604 441654
rect 332004 441334 332604 441418
rect 332004 441098 332186 441334
rect 332422 441098 332604 441334
rect 332004 405654 332604 441098
rect 332004 405418 332186 405654
rect 332422 405418 332604 405654
rect 332004 405334 332604 405418
rect 332004 405098 332186 405334
rect 332422 405098 332604 405334
rect 332004 369654 332604 405098
rect 332004 369418 332186 369654
rect 332422 369418 332604 369654
rect 332004 369334 332604 369418
rect 332004 369098 332186 369334
rect 332422 369098 332604 369334
rect 332004 333654 332604 369098
rect 332004 333418 332186 333654
rect 332422 333418 332604 333654
rect 332004 333334 332604 333418
rect 332004 333098 332186 333334
rect 332422 333098 332604 333334
rect 332004 297654 332604 333098
rect 332004 297418 332186 297654
rect 332422 297418 332604 297654
rect 332004 297334 332604 297418
rect 332004 297098 332186 297334
rect 332422 297098 332604 297334
rect 332004 261654 332604 297098
rect 332004 261418 332186 261654
rect 332422 261418 332604 261654
rect 332004 261334 332604 261418
rect 332004 261098 332186 261334
rect 332422 261098 332604 261334
rect 332004 225654 332604 261098
rect 332004 225418 332186 225654
rect 332422 225418 332604 225654
rect 332004 225334 332604 225418
rect 332004 225098 332186 225334
rect 332422 225098 332604 225334
rect 332004 189654 332604 225098
rect 332004 189418 332186 189654
rect 332422 189418 332604 189654
rect 332004 189334 332604 189418
rect 332004 189098 332186 189334
rect 332422 189098 332604 189334
rect 332004 153654 332604 189098
rect 332004 153418 332186 153654
rect 332422 153418 332604 153654
rect 332004 153334 332604 153418
rect 332004 153098 332186 153334
rect 332422 153098 332604 153334
rect 329603 147796 329669 147797
rect 329603 147732 329604 147796
rect 329668 147732 329669 147796
rect 329603 147731 329669 147732
rect 329606 144941 329666 147731
rect 329603 144940 329669 144941
rect 329603 144876 329604 144940
rect 329668 144876 329669 144940
rect 329603 144875 329669 144876
rect 329603 128484 329669 128485
rect 329603 128420 329604 128484
rect 329668 128420 329669 128484
rect 329603 128419 329669 128420
rect 329606 125629 329666 128419
rect 329603 125628 329669 125629
rect 329603 125564 329604 125628
rect 329668 125564 329669 125628
rect 329603 125563 329669 125564
rect 328404 113818 328586 114054
rect 328822 113818 329004 114054
rect 328404 113734 329004 113818
rect 328404 113498 328586 113734
rect 328822 113498 329004 113734
rect 328404 78054 329004 113498
rect 332004 117654 332604 153098
rect 332004 117418 332186 117654
rect 332422 117418 332604 117654
rect 332004 117334 332604 117418
rect 332004 117098 332186 117334
rect 332422 117098 332604 117334
rect 329603 109172 329669 109173
rect 329603 109108 329604 109172
rect 329668 109108 329669 109172
rect 329603 109107 329669 109108
rect 329606 106317 329666 109107
rect 329603 106316 329669 106317
rect 329603 106252 329604 106316
rect 329668 106252 329669 106316
rect 329603 106251 329669 106252
rect 328404 77818 328586 78054
rect 328822 77818 329004 78054
rect 328404 77734 329004 77818
rect 328404 77498 328586 77734
rect 328822 77498 329004 77734
rect 328404 42054 329004 77498
rect 332004 81654 332604 117098
rect 332004 81418 332186 81654
rect 332422 81418 332604 81654
rect 332004 81334 332604 81418
rect 332004 81098 332186 81334
rect 332422 81098 332604 81334
rect 329419 51236 329485 51237
rect 329419 51172 329420 51236
rect 329484 51172 329485 51236
rect 329419 51171 329485 51172
rect 329422 48381 329482 51171
rect 329419 48380 329485 48381
rect 329419 48316 329420 48380
rect 329484 48316 329485 48380
rect 329419 48315 329485 48316
rect 328404 41818 328586 42054
rect 328822 41818 329004 42054
rect 328404 41734 329004 41818
rect 328404 41498 328586 41734
rect 328822 41498 329004 41734
rect 327027 40628 327093 40629
rect 327027 40564 327028 40628
rect 327092 40564 327093 40628
rect 327027 40563 327093 40564
rect 327030 40357 327090 40563
rect 327027 40356 327093 40357
rect 327027 40292 327028 40356
rect 327092 40292 327093 40356
rect 327027 40291 327093 40292
rect 324804 38218 324986 38454
rect 325222 38218 325404 38454
rect 324804 38134 325404 38218
rect 324804 37898 324986 38134
rect 325222 37898 325404 38134
rect 324804 2454 325404 37898
rect 324804 2218 324986 2454
rect 325222 2218 325404 2454
rect 324804 2134 325404 2218
rect 324804 1898 324986 2134
rect 325222 1898 325404 2134
rect 324804 -346 325404 1898
rect 324804 -582 324986 -346
rect 325222 -582 325404 -346
rect 324804 -666 325404 -582
rect 324804 -902 324986 -666
rect 325222 -902 325404 -666
rect 324804 -1844 325404 -902
rect 328404 6054 329004 41498
rect 328404 5818 328586 6054
rect 328822 5818 329004 6054
rect 328404 5734 329004 5818
rect 328404 5498 328586 5734
rect 328822 5498 329004 5734
rect 328404 -2186 329004 5498
rect 328404 -2422 328586 -2186
rect 328822 -2422 329004 -2186
rect 328404 -2506 329004 -2422
rect 328404 -2742 328586 -2506
rect 328822 -2742 329004 -2506
rect 328404 -3684 329004 -2742
rect 332004 45654 332604 81098
rect 332004 45418 332186 45654
rect 332422 45418 332604 45654
rect 332004 45334 332604 45418
rect 332004 45098 332186 45334
rect 332422 45098 332604 45334
rect 332004 9654 332604 45098
rect 332004 9418 332186 9654
rect 332422 9418 332604 9654
rect 332004 9334 332604 9418
rect 332004 9098 332186 9334
rect 332422 9098 332604 9334
rect 332004 -4026 332604 9098
rect 332004 -4262 332186 -4026
rect 332422 -4262 332604 -4026
rect 332004 -4346 332604 -4262
rect 332004 -4582 332186 -4346
rect 332422 -4582 332604 -4346
rect 332004 -5524 332604 -4582
rect 335604 517254 336204 552698
rect 342804 705758 343404 705780
rect 342804 705522 342986 705758
rect 343222 705522 343404 705758
rect 342804 705438 343404 705522
rect 342804 705202 342986 705438
rect 343222 705202 343404 705438
rect 342804 668454 343404 705202
rect 342804 668218 342986 668454
rect 343222 668218 343404 668454
rect 342804 668134 343404 668218
rect 342804 667898 342986 668134
rect 343222 667898 343404 668134
rect 342804 632454 343404 667898
rect 342804 632218 342986 632454
rect 343222 632218 343404 632454
rect 342804 632134 343404 632218
rect 342804 631898 342986 632134
rect 343222 631898 343404 632134
rect 342804 596454 343404 631898
rect 342804 596218 342986 596454
rect 343222 596218 343404 596454
rect 342804 596134 343404 596218
rect 342804 595898 342986 596134
rect 343222 595898 343404 596134
rect 342804 560454 343404 595898
rect 342804 560218 342986 560454
rect 343222 560218 343404 560454
rect 342804 560134 343404 560218
rect 342804 559898 342986 560134
rect 343222 559898 343404 560134
rect 342804 524454 343404 559898
rect 342804 524218 342986 524454
rect 343222 524218 343404 524454
rect 342804 524134 343404 524218
rect 342804 523898 342986 524134
rect 343222 523898 343404 524134
rect 336411 518804 336477 518805
rect 336411 518740 336412 518804
rect 336476 518740 336477 518804
rect 336411 518739 336477 518740
rect 336414 517938 336474 518739
rect 335604 517018 335786 517254
rect 336022 517018 336204 517254
rect 335604 516934 336204 517018
rect 335604 516698 335786 516934
rect 336022 516698 336204 516934
rect 335604 481254 336204 516698
rect 335604 481018 335786 481254
rect 336022 481018 336204 481254
rect 335604 480934 336204 481018
rect 335604 480698 335786 480934
rect 336022 480698 336204 480934
rect 335604 445254 336204 480698
rect 335604 445018 335786 445254
rect 336022 445018 336204 445254
rect 335604 444934 336204 445018
rect 335604 444698 335786 444934
rect 336022 444698 336204 444934
rect 335604 409254 336204 444698
rect 335604 409018 335786 409254
rect 336022 409018 336204 409254
rect 335604 408934 336204 409018
rect 335604 408698 335786 408934
rect 336022 408698 336204 408934
rect 335604 373254 336204 408698
rect 335604 373018 335786 373254
rect 336022 373018 336204 373254
rect 335604 372934 336204 373018
rect 335604 372698 335786 372934
rect 336022 372698 336204 372934
rect 335604 337254 336204 372698
rect 335604 337018 335786 337254
rect 336022 337018 336204 337254
rect 335604 336934 336204 337018
rect 335604 336698 335786 336934
rect 336022 336698 336204 336934
rect 335604 301254 336204 336698
rect 335604 301018 335786 301254
rect 336022 301018 336204 301254
rect 335604 300934 336204 301018
rect 335604 300698 335786 300934
rect 336022 300698 336204 300934
rect 335604 265254 336204 300698
rect 335604 265018 335786 265254
rect 336022 265018 336204 265254
rect 335604 264934 336204 265018
rect 335604 264698 335786 264934
rect 336022 264698 336204 264934
rect 335604 229254 336204 264698
rect 335604 229018 335786 229254
rect 336022 229018 336204 229254
rect 335604 228934 336204 229018
rect 335604 228698 335786 228934
rect 336022 228698 336204 228934
rect 335604 193254 336204 228698
rect 335604 193018 335786 193254
rect 336022 193018 336204 193254
rect 335604 192934 336204 193018
rect 335604 192698 335786 192934
rect 336022 192698 336204 192934
rect 335604 157254 336204 192698
rect 335604 157018 335786 157254
rect 336022 157018 336204 157254
rect 335604 156934 336204 157018
rect 335604 156698 335786 156934
rect 336022 156698 336204 156934
rect 335604 121254 336204 156698
rect 335604 121018 335786 121254
rect 336022 121018 336204 121254
rect 335604 120934 336204 121018
rect 335604 120698 335786 120934
rect 336022 120698 336204 120934
rect 335604 85254 336204 120698
rect 335604 85018 335786 85254
rect 336022 85018 336204 85254
rect 335604 84934 336204 85018
rect 335604 84698 335786 84934
rect 336022 84698 336204 84934
rect 335604 49254 336204 84698
rect 335604 49018 335786 49254
rect 336022 49018 336204 49254
rect 335604 48934 336204 49018
rect 335604 48698 335786 48934
rect 336022 48698 336204 48934
rect 335604 13254 336204 48698
rect 342804 488454 343404 523898
rect 342804 488218 342986 488454
rect 343222 488218 343404 488454
rect 342804 488134 343404 488218
rect 342804 487898 342986 488134
rect 343222 487898 343404 488134
rect 342804 452454 343404 487898
rect 342804 452218 342986 452454
rect 343222 452218 343404 452454
rect 342804 452134 343404 452218
rect 342804 451898 342986 452134
rect 343222 451898 343404 452134
rect 342804 416454 343404 451898
rect 342804 416218 342986 416454
rect 343222 416218 343404 416454
rect 342804 416134 343404 416218
rect 342804 415898 342986 416134
rect 343222 415898 343404 416134
rect 342804 380454 343404 415898
rect 342804 380218 342986 380454
rect 343222 380218 343404 380454
rect 342804 380134 343404 380218
rect 342804 379898 342986 380134
rect 343222 379898 343404 380134
rect 342804 344454 343404 379898
rect 342804 344218 342986 344454
rect 343222 344218 343404 344454
rect 342804 344134 343404 344218
rect 342804 343898 342986 344134
rect 343222 343898 343404 344134
rect 342804 308454 343404 343898
rect 342804 308218 342986 308454
rect 343222 308218 343404 308454
rect 342804 308134 343404 308218
rect 342804 307898 342986 308134
rect 343222 307898 343404 308134
rect 342804 272454 343404 307898
rect 342804 272218 342986 272454
rect 343222 272218 343404 272454
rect 342804 272134 343404 272218
rect 342804 271898 342986 272134
rect 343222 271898 343404 272134
rect 342804 236454 343404 271898
rect 342804 236218 342986 236454
rect 343222 236218 343404 236454
rect 342804 236134 343404 236218
rect 342804 235898 342986 236134
rect 343222 235898 343404 236134
rect 342804 200454 343404 235898
rect 342804 200218 342986 200454
rect 343222 200218 343404 200454
rect 342804 200134 343404 200218
rect 342804 199898 342986 200134
rect 343222 199898 343404 200134
rect 342804 164454 343404 199898
rect 342804 164218 342986 164454
rect 343222 164218 343404 164454
rect 342804 164134 343404 164218
rect 342804 163898 342986 164134
rect 343222 163898 343404 164134
rect 342804 128454 343404 163898
rect 342804 128218 342986 128454
rect 343222 128218 343404 128454
rect 342804 128134 343404 128218
rect 342804 127898 342986 128134
rect 343222 127898 343404 128134
rect 342804 92454 343404 127898
rect 342804 92218 342986 92454
rect 343222 92218 343404 92454
rect 342804 92134 343404 92218
rect 342804 91898 342986 92134
rect 343222 91898 343404 92134
rect 342804 56454 343404 91898
rect 342804 56218 342986 56454
rect 343222 56218 343404 56454
rect 342804 56134 343404 56218
rect 342804 55898 342986 56134
rect 343222 55898 343404 56134
rect 336779 40628 336845 40629
rect 336779 40564 336780 40628
rect 336844 40564 336845 40628
rect 336779 40563 336845 40564
rect 336595 40492 336661 40493
rect 336595 40428 336596 40492
rect 336660 40490 336661 40492
rect 336782 40490 336842 40563
rect 336660 40430 336842 40490
rect 336660 40428 336661 40430
rect 336595 40427 336661 40428
rect 335604 13018 335786 13254
rect 336022 13018 336204 13254
rect 335604 12934 336204 13018
rect 335604 12698 335786 12934
rect 336022 12698 336204 12934
rect 317604 -7022 317786 -6786
rect 318022 -7022 318204 -6786
rect 317604 -7106 318204 -7022
rect 317604 -7342 317786 -7106
rect 318022 -7342 318204 -7106
rect 317604 -7364 318204 -7342
rect 335604 -5866 336204 12698
rect 342804 20454 343404 55898
rect 342804 20218 342986 20454
rect 343222 20218 343404 20454
rect 342804 20134 343404 20218
rect 342804 19898 342986 20134
rect 343222 19898 343404 20134
rect 342804 -1266 343404 19898
rect 342804 -1502 342986 -1266
rect 343222 -1502 343404 -1266
rect 342804 -1586 343404 -1502
rect 342804 -1822 342986 -1586
rect 343222 -1822 343404 -1586
rect 342804 -1844 343404 -1822
rect 346404 672054 347004 707042
rect 346404 671818 346586 672054
rect 346822 671818 347004 672054
rect 346404 671734 347004 671818
rect 346404 671498 346586 671734
rect 346822 671498 347004 671734
rect 346404 636054 347004 671498
rect 346404 635818 346586 636054
rect 346822 635818 347004 636054
rect 346404 635734 347004 635818
rect 346404 635498 346586 635734
rect 346822 635498 347004 635734
rect 346404 600054 347004 635498
rect 346404 599818 346586 600054
rect 346822 599818 347004 600054
rect 346404 599734 347004 599818
rect 346404 599498 346586 599734
rect 346822 599498 347004 599734
rect 346404 564054 347004 599498
rect 346404 563818 346586 564054
rect 346822 563818 347004 564054
rect 346404 563734 347004 563818
rect 346404 563498 346586 563734
rect 346822 563498 347004 563734
rect 346404 528054 347004 563498
rect 346404 527818 346586 528054
rect 346822 527818 347004 528054
rect 346404 527734 347004 527818
rect 346404 527498 346586 527734
rect 346822 527498 347004 527734
rect 346404 492054 347004 527498
rect 346404 491818 346586 492054
rect 346822 491818 347004 492054
rect 346404 491734 347004 491818
rect 346404 491498 346586 491734
rect 346822 491498 347004 491734
rect 346404 456054 347004 491498
rect 346404 455818 346586 456054
rect 346822 455818 347004 456054
rect 346404 455734 347004 455818
rect 346404 455498 346586 455734
rect 346822 455498 347004 455734
rect 346404 420054 347004 455498
rect 346404 419818 346586 420054
rect 346822 419818 347004 420054
rect 346404 419734 347004 419818
rect 346404 419498 346586 419734
rect 346822 419498 347004 419734
rect 346404 384054 347004 419498
rect 346404 383818 346586 384054
rect 346822 383818 347004 384054
rect 346404 383734 347004 383818
rect 346404 383498 346586 383734
rect 346822 383498 347004 383734
rect 346404 348054 347004 383498
rect 346404 347818 346586 348054
rect 346822 347818 347004 348054
rect 346404 347734 347004 347818
rect 346404 347498 346586 347734
rect 346822 347498 347004 347734
rect 346404 312054 347004 347498
rect 346404 311818 346586 312054
rect 346822 311818 347004 312054
rect 346404 311734 347004 311818
rect 346404 311498 346586 311734
rect 346822 311498 347004 311734
rect 346404 276054 347004 311498
rect 346404 275818 346586 276054
rect 346822 275818 347004 276054
rect 346404 275734 347004 275818
rect 346404 275498 346586 275734
rect 346822 275498 347004 275734
rect 346404 240054 347004 275498
rect 346404 239818 346586 240054
rect 346822 239818 347004 240054
rect 346404 239734 347004 239818
rect 346404 239498 346586 239734
rect 346822 239498 347004 239734
rect 346404 204054 347004 239498
rect 346404 203818 346586 204054
rect 346822 203818 347004 204054
rect 346404 203734 347004 203818
rect 346404 203498 346586 203734
rect 346822 203498 347004 203734
rect 346404 168054 347004 203498
rect 346404 167818 346586 168054
rect 346822 167818 347004 168054
rect 346404 167734 347004 167818
rect 346404 167498 346586 167734
rect 346822 167498 347004 167734
rect 346404 132054 347004 167498
rect 346404 131818 346586 132054
rect 346822 131818 347004 132054
rect 346404 131734 347004 131818
rect 346404 131498 346586 131734
rect 346822 131498 347004 131734
rect 346404 96054 347004 131498
rect 346404 95818 346586 96054
rect 346822 95818 347004 96054
rect 346404 95734 347004 95818
rect 346404 95498 346586 95734
rect 346822 95498 347004 95734
rect 346404 60054 347004 95498
rect 346404 59818 346586 60054
rect 346822 59818 347004 60054
rect 346404 59734 347004 59818
rect 346404 59498 346586 59734
rect 346822 59498 347004 59734
rect 346404 24054 347004 59498
rect 346404 23818 346586 24054
rect 346822 23818 347004 24054
rect 346404 23734 347004 23818
rect 346404 23498 346586 23734
rect 346822 23498 347004 23734
rect 346404 -3106 347004 23498
rect 346404 -3342 346586 -3106
rect 346822 -3342 347004 -3106
rect 346404 -3426 347004 -3342
rect 346404 -3662 346586 -3426
rect 346822 -3662 347004 -3426
rect 346404 -3684 347004 -3662
rect 350004 675654 350604 708882
rect 350004 675418 350186 675654
rect 350422 675418 350604 675654
rect 350004 675334 350604 675418
rect 350004 675098 350186 675334
rect 350422 675098 350604 675334
rect 350004 639654 350604 675098
rect 350004 639418 350186 639654
rect 350422 639418 350604 639654
rect 350004 639334 350604 639418
rect 350004 639098 350186 639334
rect 350422 639098 350604 639334
rect 350004 603654 350604 639098
rect 350004 603418 350186 603654
rect 350422 603418 350604 603654
rect 350004 603334 350604 603418
rect 350004 603098 350186 603334
rect 350422 603098 350604 603334
rect 350004 567654 350604 603098
rect 350004 567418 350186 567654
rect 350422 567418 350604 567654
rect 350004 567334 350604 567418
rect 350004 567098 350186 567334
rect 350422 567098 350604 567334
rect 350004 531654 350604 567098
rect 350004 531418 350186 531654
rect 350422 531418 350604 531654
rect 350004 531334 350604 531418
rect 350004 531098 350186 531334
rect 350422 531098 350604 531334
rect 350004 495654 350604 531098
rect 350004 495418 350186 495654
rect 350422 495418 350604 495654
rect 350004 495334 350604 495418
rect 350004 495098 350186 495334
rect 350422 495098 350604 495334
rect 350004 459654 350604 495098
rect 350004 459418 350186 459654
rect 350422 459418 350604 459654
rect 350004 459334 350604 459418
rect 350004 459098 350186 459334
rect 350422 459098 350604 459334
rect 350004 423654 350604 459098
rect 350004 423418 350186 423654
rect 350422 423418 350604 423654
rect 350004 423334 350604 423418
rect 350004 423098 350186 423334
rect 350422 423098 350604 423334
rect 350004 387654 350604 423098
rect 350004 387418 350186 387654
rect 350422 387418 350604 387654
rect 350004 387334 350604 387418
rect 350004 387098 350186 387334
rect 350422 387098 350604 387334
rect 350004 351654 350604 387098
rect 350004 351418 350186 351654
rect 350422 351418 350604 351654
rect 350004 351334 350604 351418
rect 350004 351098 350186 351334
rect 350422 351098 350604 351334
rect 350004 315654 350604 351098
rect 350004 315418 350186 315654
rect 350422 315418 350604 315654
rect 350004 315334 350604 315418
rect 350004 315098 350186 315334
rect 350422 315098 350604 315334
rect 350004 279654 350604 315098
rect 350004 279418 350186 279654
rect 350422 279418 350604 279654
rect 350004 279334 350604 279418
rect 350004 279098 350186 279334
rect 350422 279098 350604 279334
rect 350004 243654 350604 279098
rect 350004 243418 350186 243654
rect 350422 243418 350604 243654
rect 350004 243334 350604 243418
rect 350004 243098 350186 243334
rect 350422 243098 350604 243334
rect 350004 207654 350604 243098
rect 350004 207418 350186 207654
rect 350422 207418 350604 207654
rect 350004 207334 350604 207418
rect 350004 207098 350186 207334
rect 350422 207098 350604 207334
rect 350004 171654 350604 207098
rect 350004 171418 350186 171654
rect 350422 171418 350604 171654
rect 350004 171334 350604 171418
rect 350004 171098 350186 171334
rect 350422 171098 350604 171334
rect 350004 135654 350604 171098
rect 350004 135418 350186 135654
rect 350422 135418 350604 135654
rect 350004 135334 350604 135418
rect 350004 135098 350186 135334
rect 350422 135098 350604 135334
rect 350004 99654 350604 135098
rect 350004 99418 350186 99654
rect 350422 99418 350604 99654
rect 350004 99334 350604 99418
rect 350004 99098 350186 99334
rect 350422 99098 350604 99334
rect 350004 63654 350604 99098
rect 350004 63418 350186 63654
rect 350422 63418 350604 63654
rect 350004 63334 350604 63418
rect 350004 63098 350186 63334
rect 350422 63098 350604 63334
rect 350004 27654 350604 63098
rect 350004 27418 350186 27654
rect 350422 27418 350604 27654
rect 350004 27334 350604 27418
rect 350004 27098 350186 27334
rect 350422 27098 350604 27334
rect 350004 -4946 350604 27098
rect 350004 -5182 350186 -4946
rect 350422 -5182 350604 -4946
rect 350004 -5266 350604 -5182
rect 350004 -5502 350186 -5266
rect 350422 -5502 350604 -5266
rect 350004 -5524 350604 -5502
rect 353604 679254 354204 710722
rect 371604 710358 372204 711300
rect 371604 710122 371786 710358
rect 372022 710122 372204 710358
rect 371604 710038 372204 710122
rect 371604 709802 371786 710038
rect 372022 709802 372204 710038
rect 368004 708518 368604 709460
rect 368004 708282 368186 708518
rect 368422 708282 368604 708518
rect 368004 708198 368604 708282
rect 368004 707962 368186 708198
rect 368422 707962 368604 708198
rect 364404 706678 365004 707620
rect 364404 706442 364586 706678
rect 364822 706442 365004 706678
rect 364404 706358 365004 706442
rect 364404 706122 364586 706358
rect 364822 706122 365004 706358
rect 353604 679018 353786 679254
rect 354022 679018 354204 679254
rect 353604 678934 354204 679018
rect 353604 678698 353786 678934
rect 354022 678698 354204 678934
rect 353604 643254 354204 678698
rect 353604 643018 353786 643254
rect 354022 643018 354204 643254
rect 353604 642934 354204 643018
rect 353604 642698 353786 642934
rect 354022 642698 354204 642934
rect 353604 607254 354204 642698
rect 353604 607018 353786 607254
rect 354022 607018 354204 607254
rect 353604 606934 354204 607018
rect 353604 606698 353786 606934
rect 354022 606698 354204 606934
rect 353604 571254 354204 606698
rect 353604 571018 353786 571254
rect 354022 571018 354204 571254
rect 353604 570934 354204 571018
rect 353604 570698 353786 570934
rect 354022 570698 354204 570934
rect 353604 535254 354204 570698
rect 353604 535018 353786 535254
rect 354022 535018 354204 535254
rect 353604 534934 354204 535018
rect 353604 534698 353786 534934
rect 354022 534698 354204 534934
rect 353604 499254 354204 534698
rect 360804 704838 361404 705780
rect 360804 704602 360986 704838
rect 361222 704602 361404 704838
rect 360804 704518 361404 704602
rect 360804 704282 360986 704518
rect 361222 704282 361404 704518
rect 360804 686454 361404 704282
rect 360804 686218 360986 686454
rect 361222 686218 361404 686454
rect 360804 686134 361404 686218
rect 360804 685898 360986 686134
rect 361222 685898 361404 686134
rect 360804 650454 361404 685898
rect 360804 650218 360986 650454
rect 361222 650218 361404 650454
rect 360804 650134 361404 650218
rect 360804 649898 360986 650134
rect 361222 649898 361404 650134
rect 360804 614454 361404 649898
rect 360804 614218 360986 614454
rect 361222 614218 361404 614454
rect 360804 614134 361404 614218
rect 360804 613898 360986 614134
rect 361222 613898 361404 614134
rect 360804 578454 361404 613898
rect 360804 578218 360986 578454
rect 361222 578218 361404 578454
rect 360804 578134 361404 578218
rect 360804 577898 360986 578134
rect 361222 577898 361404 578134
rect 360804 542454 361404 577898
rect 360804 542218 360986 542454
rect 361222 542218 361404 542454
rect 360804 542134 361404 542218
rect 360804 541898 360986 542134
rect 361222 541898 361404 542134
rect 359779 523020 359845 523021
rect 359779 522956 359780 523020
rect 359844 522956 359845 523020
rect 359779 522955 359845 522956
rect 359595 522884 359661 522885
rect 359595 522820 359596 522884
rect 359660 522820 359661 522884
rect 359595 522819 359661 522820
rect 359411 522748 359477 522749
rect 359411 522684 359412 522748
rect 359476 522684 359477 522748
rect 359411 522683 359477 522684
rect 359043 519348 359109 519349
rect 359043 519284 359044 519348
rect 359108 519284 359109 519348
rect 359043 519283 359109 519284
rect 353604 499018 353786 499254
rect 354022 499018 354204 499254
rect 353604 498934 354204 499018
rect 353604 498698 353786 498934
rect 354022 498698 354204 498934
rect 353604 463254 354204 498698
rect 353604 463018 353786 463254
rect 354022 463018 354204 463254
rect 353604 462934 354204 463018
rect 353604 462698 353786 462934
rect 354022 462698 354204 462934
rect 353604 427254 354204 462698
rect 353604 427018 353786 427254
rect 354022 427018 354204 427254
rect 353604 426934 354204 427018
rect 353604 426698 353786 426934
rect 354022 426698 354204 426934
rect 353604 391254 354204 426698
rect 353604 391018 353786 391254
rect 354022 391018 354204 391254
rect 353604 390934 354204 391018
rect 353604 390698 353786 390934
rect 354022 390698 354204 390934
rect 353604 355254 354204 390698
rect 353604 355018 353786 355254
rect 354022 355018 354204 355254
rect 353604 354934 354204 355018
rect 353604 354698 353786 354934
rect 354022 354698 354204 354934
rect 353604 319254 354204 354698
rect 353604 319018 353786 319254
rect 354022 319018 354204 319254
rect 353604 318934 354204 319018
rect 353604 318698 353786 318934
rect 354022 318698 354204 318934
rect 353604 283254 354204 318698
rect 353604 283018 353786 283254
rect 354022 283018 354204 283254
rect 353604 282934 354204 283018
rect 353604 282698 353786 282934
rect 354022 282698 354204 282934
rect 353604 247254 354204 282698
rect 353604 247018 353786 247254
rect 354022 247018 354204 247254
rect 353604 246934 354204 247018
rect 353604 246698 353786 246934
rect 354022 246698 354204 246934
rect 353604 211254 354204 246698
rect 353604 211018 353786 211254
rect 354022 211018 354204 211254
rect 353604 210934 354204 211018
rect 353604 210698 353786 210934
rect 354022 210698 354204 210934
rect 353604 175254 354204 210698
rect 353604 175018 353786 175254
rect 354022 175018 354204 175254
rect 353604 174934 354204 175018
rect 353604 174698 353786 174934
rect 354022 174698 354204 174934
rect 353604 139254 354204 174698
rect 353604 139018 353786 139254
rect 354022 139018 354204 139254
rect 353604 138934 354204 139018
rect 353604 138698 353786 138934
rect 354022 138698 354204 138934
rect 353604 103254 354204 138698
rect 353604 103018 353786 103254
rect 354022 103018 354204 103254
rect 353604 102934 354204 103018
rect 353604 102698 353786 102934
rect 354022 102698 354204 102934
rect 353604 67254 354204 102698
rect 353604 67018 353786 67254
rect 354022 67018 354204 67254
rect 353604 66934 354204 67018
rect 353604 66698 353786 66934
rect 354022 66698 354204 66934
rect 353604 31254 354204 66698
rect 359046 64837 359106 519283
rect 359414 251293 359474 522683
rect 359598 298213 359658 522819
rect 359782 485893 359842 522955
rect 360804 506454 361404 541898
rect 364404 690054 365004 706122
rect 364404 689818 364586 690054
rect 364822 689818 365004 690054
rect 364404 689734 365004 689818
rect 364404 689498 364586 689734
rect 364822 689498 365004 689734
rect 364404 654054 365004 689498
rect 364404 653818 364586 654054
rect 364822 653818 365004 654054
rect 364404 653734 365004 653818
rect 364404 653498 364586 653734
rect 364822 653498 365004 653734
rect 364404 618054 365004 653498
rect 364404 617818 364586 618054
rect 364822 617818 365004 618054
rect 364404 617734 365004 617818
rect 364404 617498 364586 617734
rect 364822 617498 365004 617734
rect 364404 582054 365004 617498
rect 364404 581818 364586 582054
rect 364822 581818 365004 582054
rect 364404 581734 365004 581818
rect 364404 581498 364586 581734
rect 364822 581498 365004 581734
rect 364404 546054 365004 581498
rect 364404 545818 364586 546054
rect 364822 545818 365004 546054
rect 364404 545734 365004 545818
rect 364404 545498 364586 545734
rect 364822 545498 365004 545734
rect 361619 519348 361685 519349
rect 361619 519284 361620 519348
rect 361684 519284 361685 519348
rect 361619 519283 361685 519284
rect 362907 519348 362973 519349
rect 362907 519284 362908 519348
rect 362972 519284 362973 519348
rect 362907 519283 362973 519284
rect 360804 506218 360986 506454
rect 361222 506218 361404 506454
rect 360804 506134 361404 506218
rect 360804 505898 360986 506134
rect 361222 505898 361404 506134
rect 359779 485892 359845 485893
rect 359779 485828 359780 485892
rect 359844 485828 359845 485892
rect 359779 485827 359845 485828
rect 360804 470454 361404 505898
rect 360804 470218 360986 470454
rect 361222 470218 361404 470454
rect 360804 470134 361404 470218
rect 360804 469898 360986 470134
rect 361222 469898 361404 470134
rect 360804 434454 361404 469898
rect 360804 434218 360986 434454
rect 361222 434218 361404 434454
rect 360804 434134 361404 434218
rect 360804 433898 360986 434134
rect 361222 433898 361404 434134
rect 360804 398454 361404 433898
rect 360804 398218 360986 398454
rect 361222 398218 361404 398454
rect 360804 398134 361404 398218
rect 360804 397898 360986 398134
rect 361222 397898 361404 398134
rect 360804 362454 361404 397898
rect 360804 362218 360986 362454
rect 361222 362218 361404 362454
rect 360804 362134 361404 362218
rect 360804 361898 360986 362134
rect 361222 361898 361404 362134
rect 360804 326454 361404 361898
rect 360804 326218 360986 326454
rect 361222 326218 361404 326454
rect 360804 326134 361404 326218
rect 360804 325898 360986 326134
rect 361222 325898 361404 326134
rect 359595 298212 359661 298213
rect 359595 298148 359596 298212
rect 359660 298148 359661 298212
rect 359595 298147 359661 298148
rect 360804 290454 361404 325898
rect 360804 290218 360986 290454
rect 361222 290218 361404 290454
rect 360804 290134 361404 290218
rect 360804 289898 360986 290134
rect 361222 289898 361404 290134
rect 360804 254454 361404 289898
rect 360804 254218 360986 254454
rect 361222 254218 361404 254454
rect 360804 254134 361404 254218
rect 360804 253898 360986 254134
rect 361222 253898 361404 254134
rect 359411 251292 359477 251293
rect 359411 251228 359412 251292
rect 359476 251228 359477 251292
rect 359411 251227 359477 251228
rect 360804 218454 361404 253898
rect 360804 218218 360986 218454
rect 361222 218218 361404 218454
rect 360804 218134 361404 218218
rect 360804 217898 360986 218134
rect 361222 217898 361404 218134
rect 360804 182454 361404 217898
rect 360804 182218 360986 182454
rect 361222 182218 361404 182454
rect 360804 182134 361404 182218
rect 360804 181898 360986 182134
rect 361222 181898 361404 182134
rect 360804 146454 361404 181898
rect 360804 146218 360986 146454
rect 361222 146218 361404 146454
rect 360804 146134 361404 146218
rect 360804 145898 360986 146134
rect 361222 145898 361404 146134
rect 360804 110454 361404 145898
rect 360804 110218 360986 110454
rect 361222 110218 361404 110454
rect 360804 110134 361404 110218
rect 360804 109898 360986 110134
rect 361222 109898 361404 110134
rect 360804 74454 361404 109898
rect 360804 74218 360986 74454
rect 361222 74218 361404 74454
rect 360804 74134 361404 74218
rect 360804 73898 360986 74134
rect 361222 73898 361404 74134
rect 359043 64836 359109 64837
rect 359043 64772 359044 64836
rect 359108 64772 359109 64836
rect 359043 64771 359109 64772
rect 353604 31018 353786 31254
rect 354022 31018 354204 31254
rect 353604 30934 354204 31018
rect 353604 30698 353786 30934
rect 354022 30698 354204 30934
rect 335604 -6102 335786 -5866
rect 336022 -6102 336204 -5866
rect 335604 -6186 336204 -6102
rect 335604 -6422 335786 -6186
rect 336022 -6422 336204 -6186
rect 335604 -7364 336204 -6422
rect 353604 -6786 354204 30698
rect 360804 38454 361404 73898
rect 360804 38218 360986 38454
rect 361222 38218 361404 38454
rect 360804 38134 361404 38218
rect 360804 37898 360986 38134
rect 361222 37898 361404 38134
rect 360804 2454 361404 37898
rect 361622 10301 361682 519283
rect 362910 21997 362970 519283
rect 364404 510054 365004 545498
rect 368004 693654 368604 707962
rect 368004 693418 368186 693654
rect 368422 693418 368604 693654
rect 368004 693334 368604 693418
rect 368004 693098 368186 693334
rect 368422 693098 368604 693334
rect 368004 657654 368604 693098
rect 368004 657418 368186 657654
rect 368422 657418 368604 657654
rect 368004 657334 368604 657418
rect 368004 657098 368186 657334
rect 368422 657098 368604 657334
rect 368004 621654 368604 657098
rect 368004 621418 368186 621654
rect 368422 621418 368604 621654
rect 368004 621334 368604 621418
rect 368004 621098 368186 621334
rect 368422 621098 368604 621334
rect 368004 585654 368604 621098
rect 368004 585418 368186 585654
rect 368422 585418 368604 585654
rect 368004 585334 368604 585418
rect 368004 585098 368186 585334
rect 368422 585098 368604 585334
rect 368004 549654 368604 585098
rect 368004 549418 368186 549654
rect 368422 549418 368604 549654
rect 368004 549334 368604 549418
rect 368004 549098 368186 549334
rect 368422 549098 368604 549334
rect 366219 520300 366285 520301
rect 366219 520236 366220 520300
rect 366284 520236 366285 520300
rect 366219 520235 366285 520236
rect 364404 509818 364586 510054
rect 364822 509818 365004 510054
rect 364404 509734 365004 509818
rect 364404 509498 364586 509734
rect 364822 509498 365004 509734
rect 364404 474054 365004 509498
rect 364404 473818 364586 474054
rect 364822 473818 365004 474054
rect 364404 473734 365004 473818
rect 364404 473498 364586 473734
rect 364822 473498 365004 473734
rect 364404 438054 365004 473498
rect 364404 437818 364586 438054
rect 364822 437818 365004 438054
rect 364404 437734 365004 437818
rect 364404 437498 364586 437734
rect 364822 437498 365004 437734
rect 364404 402054 365004 437498
rect 364404 401818 364586 402054
rect 364822 401818 365004 402054
rect 364404 401734 365004 401818
rect 364404 401498 364586 401734
rect 364822 401498 365004 401734
rect 364404 366054 365004 401498
rect 364404 365818 364586 366054
rect 364822 365818 365004 366054
rect 364404 365734 365004 365818
rect 364404 365498 364586 365734
rect 364822 365498 365004 365734
rect 364404 330054 365004 365498
rect 364404 329818 364586 330054
rect 364822 329818 365004 330054
rect 364404 329734 365004 329818
rect 364404 329498 364586 329734
rect 364822 329498 365004 329734
rect 364404 294054 365004 329498
rect 364404 293818 364586 294054
rect 364822 293818 365004 294054
rect 364404 293734 365004 293818
rect 364404 293498 364586 293734
rect 364822 293498 365004 293734
rect 364404 258054 365004 293498
rect 364404 257818 364586 258054
rect 364822 257818 365004 258054
rect 364404 257734 365004 257818
rect 364404 257498 364586 257734
rect 364822 257498 365004 257734
rect 364404 222054 365004 257498
rect 364404 221818 364586 222054
rect 364822 221818 365004 222054
rect 364404 221734 365004 221818
rect 364404 221498 364586 221734
rect 364822 221498 365004 221734
rect 364404 186054 365004 221498
rect 366222 204645 366282 520235
rect 367323 518940 367389 518941
rect 367323 518876 367324 518940
rect 367388 518876 367389 518940
rect 367323 518875 367389 518876
rect 367326 518530 367386 518875
rect 367142 518470 367386 518530
rect 367142 518125 367202 518470
rect 367323 518396 367389 518397
rect 367323 518332 367324 518396
rect 367388 518332 367389 518396
rect 367323 518331 367389 518332
rect 367326 518125 367386 518331
rect 367139 518124 367205 518125
rect 367139 518060 367140 518124
rect 367204 518060 367205 518124
rect 367139 518059 367205 518060
rect 367323 518124 367389 518125
rect 367323 518060 367324 518124
rect 367388 518060 367389 518124
rect 367323 518059 367389 518060
rect 367323 517852 367389 517853
rect 367323 517788 367324 517852
rect 367388 517788 367389 517852
rect 367323 517787 367389 517788
rect 367326 517717 367386 517787
rect 367323 517716 367389 517717
rect 367323 517652 367324 517716
rect 367388 517652 367389 517716
rect 367323 517651 367389 517652
rect 368004 513654 368604 549098
rect 371604 697254 372204 709802
rect 389604 711278 390204 711300
rect 389604 711042 389786 711278
rect 390022 711042 390204 711278
rect 389604 710958 390204 711042
rect 389604 710722 389786 710958
rect 390022 710722 390204 710958
rect 386004 709438 386604 709460
rect 386004 709202 386186 709438
rect 386422 709202 386604 709438
rect 386004 709118 386604 709202
rect 386004 708882 386186 709118
rect 386422 708882 386604 709118
rect 382404 707598 383004 707620
rect 382404 707362 382586 707598
rect 382822 707362 383004 707598
rect 382404 707278 383004 707362
rect 382404 707042 382586 707278
rect 382822 707042 383004 707278
rect 371604 697018 371786 697254
rect 372022 697018 372204 697254
rect 371604 696934 372204 697018
rect 371604 696698 371786 696934
rect 372022 696698 372204 696934
rect 371604 661254 372204 696698
rect 371604 661018 371786 661254
rect 372022 661018 372204 661254
rect 371604 660934 372204 661018
rect 371604 660698 371786 660934
rect 372022 660698 372204 660934
rect 371604 625254 372204 660698
rect 371604 625018 371786 625254
rect 372022 625018 372204 625254
rect 371604 624934 372204 625018
rect 371604 624698 371786 624934
rect 372022 624698 372204 624934
rect 371604 589254 372204 624698
rect 371604 589018 371786 589254
rect 372022 589018 372204 589254
rect 371604 588934 372204 589018
rect 371604 588698 371786 588934
rect 372022 588698 372204 588934
rect 371604 553254 372204 588698
rect 371604 553018 371786 553254
rect 372022 553018 372204 553254
rect 371604 552934 372204 553018
rect 371604 552698 371786 552934
rect 372022 552698 372204 552934
rect 368979 517716 369045 517717
rect 368979 517652 368980 517716
rect 369044 517652 369045 517716
rect 368979 517651 369045 517652
rect 368004 513418 368186 513654
rect 368422 513418 368604 513654
rect 368004 513334 368604 513418
rect 368004 513098 368186 513334
rect 368422 513098 368604 513334
rect 367139 486436 367205 486437
rect 367139 486372 367140 486436
rect 367204 486372 367205 486436
rect 367139 486371 367205 486372
rect 367142 486165 367202 486371
rect 367139 486164 367205 486165
rect 367139 486100 367140 486164
rect 367204 486100 367205 486164
rect 367139 486099 367205 486100
rect 368004 477654 368604 513098
rect 368004 477418 368186 477654
rect 368422 477418 368604 477654
rect 368004 477334 368604 477418
rect 368004 477098 368186 477334
rect 368422 477098 368604 477334
rect 368004 441654 368604 477098
rect 368004 441418 368186 441654
rect 368422 441418 368604 441654
rect 368004 441334 368604 441418
rect 368004 441098 368186 441334
rect 368422 441098 368604 441334
rect 368004 405654 368604 441098
rect 368004 405418 368186 405654
rect 368422 405418 368604 405654
rect 368004 405334 368604 405418
rect 368004 405098 368186 405334
rect 368422 405098 368604 405334
rect 368004 369654 368604 405098
rect 368004 369418 368186 369654
rect 368422 369418 368604 369654
rect 368004 369334 368604 369418
rect 368004 369098 368186 369334
rect 368422 369098 368604 369334
rect 368004 333654 368604 369098
rect 368004 333418 368186 333654
rect 368422 333418 368604 333654
rect 368004 333334 368604 333418
rect 368004 333098 368186 333334
rect 368422 333098 368604 333334
rect 368004 297654 368604 333098
rect 368982 310861 369042 517651
rect 371604 517254 372204 552698
rect 371604 517018 371786 517254
rect 372022 517018 372204 517254
rect 371604 516934 372204 517018
rect 371604 516698 371786 516934
rect 372022 516698 372204 516934
rect 371604 481254 372204 516698
rect 371604 481018 371786 481254
rect 372022 481018 372204 481254
rect 371604 480934 372204 481018
rect 371604 480698 371786 480934
rect 372022 480698 372204 480934
rect 371604 445254 372204 480698
rect 371604 445018 371786 445254
rect 372022 445018 372204 445254
rect 371604 444934 372204 445018
rect 371604 444698 371786 444934
rect 372022 444698 372204 444934
rect 371604 409254 372204 444698
rect 371604 409018 371786 409254
rect 372022 409018 372204 409254
rect 371604 408934 372204 409018
rect 371604 408698 371786 408934
rect 372022 408698 372204 408934
rect 371604 373254 372204 408698
rect 371604 373018 371786 373254
rect 372022 373018 372204 373254
rect 371604 372934 372204 373018
rect 371604 372698 371786 372934
rect 372022 372698 372204 372934
rect 371604 337254 372204 372698
rect 371604 337018 371786 337254
rect 372022 337018 372204 337254
rect 371604 336934 372204 337018
rect 371604 336698 371786 336934
rect 372022 336698 372204 336934
rect 368979 310860 369045 310861
rect 368979 310796 368980 310860
rect 369044 310796 369045 310860
rect 368979 310795 369045 310796
rect 368004 297418 368186 297654
rect 368422 297418 368604 297654
rect 368004 297334 368604 297418
rect 368004 297098 368186 297334
rect 368422 297098 368604 297334
rect 368004 261654 368604 297098
rect 368004 261418 368186 261654
rect 368422 261418 368604 261654
rect 368004 261334 368604 261418
rect 368004 261098 368186 261334
rect 368422 261098 368604 261334
rect 368004 225654 368604 261098
rect 368004 225418 368186 225654
rect 368422 225418 368604 225654
rect 368004 225334 368604 225418
rect 368004 225098 368186 225334
rect 368422 225098 368604 225334
rect 366219 204644 366285 204645
rect 366219 204580 366220 204644
rect 366284 204580 366285 204644
rect 366219 204579 366285 204580
rect 364404 185818 364586 186054
rect 364822 185818 365004 186054
rect 364404 185734 365004 185818
rect 364404 185498 364586 185734
rect 364822 185498 365004 185734
rect 364404 150054 365004 185498
rect 364404 149818 364586 150054
rect 364822 149818 365004 150054
rect 364404 149734 365004 149818
rect 364404 149498 364586 149734
rect 364822 149498 365004 149734
rect 364404 114054 365004 149498
rect 364404 113818 364586 114054
rect 364822 113818 365004 114054
rect 364404 113734 365004 113818
rect 364404 113498 364586 113734
rect 364822 113498 365004 113734
rect 364404 78054 365004 113498
rect 364404 77818 364586 78054
rect 364822 77818 365004 78054
rect 364404 77734 365004 77818
rect 364404 77498 364586 77734
rect 364822 77498 365004 77734
rect 364404 42054 365004 77498
rect 364404 41818 364586 42054
rect 364822 41818 365004 42054
rect 364404 41734 365004 41818
rect 364404 41498 364586 41734
rect 364822 41498 365004 41734
rect 362907 21996 362973 21997
rect 362907 21932 362908 21996
rect 362972 21932 362973 21996
rect 362907 21931 362973 21932
rect 361619 10300 361685 10301
rect 361619 10236 361620 10300
rect 361684 10236 361685 10300
rect 361619 10235 361685 10236
rect 360804 2218 360986 2454
rect 361222 2218 361404 2454
rect 360804 2134 361404 2218
rect 360804 1898 360986 2134
rect 361222 1898 361404 2134
rect 360804 -346 361404 1898
rect 360804 -582 360986 -346
rect 361222 -582 361404 -346
rect 360804 -666 361404 -582
rect 360804 -902 360986 -666
rect 361222 -902 361404 -666
rect 360804 -1844 361404 -902
rect 364404 6054 365004 41498
rect 364404 5818 364586 6054
rect 364822 5818 365004 6054
rect 364404 5734 365004 5818
rect 364404 5498 364586 5734
rect 364822 5498 365004 5734
rect 364404 -2186 365004 5498
rect 364404 -2422 364586 -2186
rect 364822 -2422 365004 -2186
rect 364404 -2506 365004 -2422
rect 364404 -2742 364586 -2506
rect 364822 -2742 365004 -2506
rect 364404 -3684 365004 -2742
rect 368004 189654 368604 225098
rect 368004 189418 368186 189654
rect 368422 189418 368604 189654
rect 368004 189334 368604 189418
rect 368004 189098 368186 189334
rect 368422 189098 368604 189334
rect 368004 153654 368604 189098
rect 368004 153418 368186 153654
rect 368422 153418 368604 153654
rect 368004 153334 368604 153418
rect 368004 153098 368186 153334
rect 368422 153098 368604 153334
rect 368004 117654 368604 153098
rect 368004 117418 368186 117654
rect 368422 117418 368604 117654
rect 368004 117334 368604 117418
rect 368004 117098 368186 117334
rect 368422 117098 368604 117334
rect 368004 81654 368604 117098
rect 368004 81418 368186 81654
rect 368422 81418 368604 81654
rect 368004 81334 368604 81418
rect 368004 81098 368186 81334
rect 368422 81098 368604 81334
rect 368004 45654 368604 81098
rect 368004 45418 368186 45654
rect 368422 45418 368604 45654
rect 368004 45334 368604 45418
rect 368004 45098 368186 45334
rect 368422 45098 368604 45334
rect 368004 9654 368604 45098
rect 368004 9418 368186 9654
rect 368422 9418 368604 9654
rect 368004 9334 368604 9418
rect 368004 9098 368186 9334
rect 368422 9098 368604 9334
rect 368004 -4026 368604 9098
rect 368004 -4262 368186 -4026
rect 368422 -4262 368604 -4026
rect 368004 -4346 368604 -4262
rect 368004 -4582 368186 -4346
rect 368422 -4582 368604 -4346
rect 368004 -5524 368604 -4582
rect 371604 301254 372204 336698
rect 371604 301018 371786 301254
rect 372022 301018 372204 301254
rect 371604 300934 372204 301018
rect 371604 300698 371786 300934
rect 372022 300698 372204 300934
rect 371604 265254 372204 300698
rect 371604 265018 371786 265254
rect 372022 265018 372204 265254
rect 371604 264934 372204 265018
rect 371604 264698 371786 264934
rect 372022 264698 372204 264934
rect 371604 229254 372204 264698
rect 371604 229018 371786 229254
rect 372022 229018 372204 229254
rect 371604 228934 372204 229018
rect 371604 228698 371786 228934
rect 372022 228698 372204 228934
rect 371604 193254 372204 228698
rect 371604 193018 371786 193254
rect 372022 193018 372204 193254
rect 371604 192934 372204 193018
rect 371604 192698 371786 192934
rect 372022 192698 372204 192934
rect 371604 157254 372204 192698
rect 371604 157018 371786 157254
rect 372022 157018 372204 157254
rect 371604 156934 372204 157018
rect 371604 156698 371786 156934
rect 372022 156698 372204 156934
rect 371604 121254 372204 156698
rect 371604 121018 371786 121254
rect 372022 121018 372204 121254
rect 371604 120934 372204 121018
rect 371604 120698 371786 120934
rect 372022 120698 372204 120934
rect 371604 85254 372204 120698
rect 371604 85018 371786 85254
rect 372022 85018 372204 85254
rect 371604 84934 372204 85018
rect 371604 84698 371786 84934
rect 372022 84698 372204 84934
rect 371604 49254 372204 84698
rect 371604 49018 371786 49254
rect 372022 49018 372204 49254
rect 371604 48934 372204 49018
rect 371604 48698 371786 48934
rect 372022 48698 372204 48934
rect 371604 13254 372204 48698
rect 371604 13018 371786 13254
rect 372022 13018 372204 13254
rect 371604 12934 372204 13018
rect 371604 12698 371786 12934
rect 372022 12698 372204 12934
rect 353604 -7022 353786 -6786
rect 354022 -7022 354204 -6786
rect 353604 -7106 354204 -7022
rect 353604 -7342 353786 -7106
rect 354022 -7342 354204 -7106
rect 353604 -7364 354204 -7342
rect 371604 -5866 372204 12698
rect 378804 705758 379404 705780
rect 378804 705522 378986 705758
rect 379222 705522 379404 705758
rect 378804 705438 379404 705522
rect 378804 705202 378986 705438
rect 379222 705202 379404 705438
rect 378804 668454 379404 705202
rect 378804 668218 378986 668454
rect 379222 668218 379404 668454
rect 378804 668134 379404 668218
rect 378804 667898 378986 668134
rect 379222 667898 379404 668134
rect 378804 632454 379404 667898
rect 378804 632218 378986 632454
rect 379222 632218 379404 632454
rect 378804 632134 379404 632218
rect 378804 631898 378986 632134
rect 379222 631898 379404 632134
rect 378804 596454 379404 631898
rect 378804 596218 378986 596454
rect 379222 596218 379404 596454
rect 378804 596134 379404 596218
rect 378804 595898 378986 596134
rect 379222 595898 379404 596134
rect 378804 560454 379404 595898
rect 378804 560218 378986 560454
rect 379222 560218 379404 560454
rect 378804 560134 379404 560218
rect 378804 559898 378986 560134
rect 379222 559898 379404 560134
rect 378804 524454 379404 559898
rect 378804 524218 378986 524454
rect 379222 524218 379404 524454
rect 378804 524134 379404 524218
rect 378804 523898 378986 524134
rect 379222 523898 379404 524134
rect 378804 488454 379404 523898
rect 378804 488218 378986 488454
rect 379222 488218 379404 488454
rect 378804 488134 379404 488218
rect 378804 487898 378986 488134
rect 379222 487898 379404 488134
rect 378804 452454 379404 487898
rect 378804 452218 378986 452454
rect 379222 452218 379404 452454
rect 378804 452134 379404 452218
rect 378804 451898 378986 452134
rect 379222 451898 379404 452134
rect 378804 416454 379404 451898
rect 378804 416218 378986 416454
rect 379222 416218 379404 416454
rect 378804 416134 379404 416218
rect 378804 415898 378986 416134
rect 379222 415898 379404 416134
rect 378804 380454 379404 415898
rect 378804 380218 378986 380454
rect 379222 380218 379404 380454
rect 378804 380134 379404 380218
rect 378804 379898 378986 380134
rect 379222 379898 379404 380134
rect 378804 344454 379404 379898
rect 378804 344218 378986 344454
rect 379222 344218 379404 344454
rect 378804 344134 379404 344218
rect 378804 343898 378986 344134
rect 379222 343898 379404 344134
rect 378804 308454 379404 343898
rect 378804 308218 378986 308454
rect 379222 308218 379404 308454
rect 378804 308134 379404 308218
rect 378804 307898 378986 308134
rect 379222 307898 379404 308134
rect 378804 272454 379404 307898
rect 378804 272218 378986 272454
rect 379222 272218 379404 272454
rect 378804 272134 379404 272218
rect 378804 271898 378986 272134
rect 379222 271898 379404 272134
rect 378804 236454 379404 271898
rect 378804 236218 378986 236454
rect 379222 236218 379404 236454
rect 378804 236134 379404 236218
rect 378804 235898 378986 236134
rect 379222 235898 379404 236134
rect 378804 200454 379404 235898
rect 378804 200218 378986 200454
rect 379222 200218 379404 200454
rect 378804 200134 379404 200218
rect 378804 199898 378986 200134
rect 379222 199898 379404 200134
rect 378804 164454 379404 199898
rect 378804 164218 378986 164454
rect 379222 164218 379404 164454
rect 378804 164134 379404 164218
rect 378804 163898 378986 164134
rect 379222 163898 379404 164134
rect 378804 128454 379404 163898
rect 378804 128218 378986 128454
rect 379222 128218 379404 128454
rect 378804 128134 379404 128218
rect 378804 127898 378986 128134
rect 379222 127898 379404 128134
rect 378804 92454 379404 127898
rect 378804 92218 378986 92454
rect 379222 92218 379404 92454
rect 378804 92134 379404 92218
rect 378804 91898 378986 92134
rect 379222 91898 379404 92134
rect 378804 56454 379404 91898
rect 378804 56218 378986 56454
rect 379222 56218 379404 56454
rect 378804 56134 379404 56218
rect 378804 55898 378986 56134
rect 379222 55898 379404 56134
rect 378804 20454 379404 55898
rect 378804 20218 378986 20454
rect 379222 20218 379404 20454
rect 378804 20134 379404 20218
rect 378804 19898 378986 20134
rect 379222 19898 379404 20134
rect 378804 -1266 379404 19898
rect 378804 -1502 378986 -1266
rect 379222 -1502 379404 -1266
rect 378804 -1586 379404 -1502
rect 378804 -1822 378986 -1586
rect 379222 -1822 379404 -1586
rect 378804 -1844 379404 -1822
rect 382404 672054 383004 707042
rect 382404 671818 382586 672054
rect 382822 671818 383004 672054
rect 382404 671734 383004 671818
rect 382404 671498 382586 671734
rect 382822 671498 383004 671734
rect 382404 636054 383004 671498
rect 382404 635818 382586 636054
rect 382822 635818 383004 636054
rect 382404 635734 383004 635818
rect 382404 635498 382586 635734
rect 382822 635498 383004 635734
rect 382404 600054 383004 635498
rect 382404 599818 382586 600054
rect 382822 599818 383004 600054
rect 382404 599734 383004 599818
rect 382404 599498 382586 599734
rect 382822 599498 383004 599734
rect 382404 564054 383004 599498
rect 382404 563818 382586 564054
rect 382822 563818 383004 564054
rect 382404 563734 383004 563818
rect 382404 563498 382586 563734
rect 382822 563498 383004 563734
rect 382404 528054 383004 563498
rect 382404 527818 382586 528054
rect 382822 527818 383004 528054
rect 382404 527734 383004 527818
rect 382404 527498 382586 527734
rect 382822 527498 383004 527734
rect 382404 492054 383004 527498
rect 382404 491818 382586 492054
rect 382822 491818 383004 492054
rect 382404 491734 383004 491818
rect 382404 491498 382586 491734
rect 382822 491498 383004 491734
rect 382404 456054 383004 491498
rect 386004 675654 386604 708882
rect 386004 675418 386186 675654
rect 386422 675418 386604 675654
rect 386004 675334 386604 675418
rect 386004 675098 386186 675334
rect 386422 675098 386604 675334
rect 386004 639654 386604 675098
rect 386004 639418 386186 639654
rect 386422 639418 386604 639654
rect 386004 639334 386604 639418
rect 386004 639098 386186 639334
rect 386422 639098 386604 639334
rect 386004 603654 386604 639098
rect 386004 603418 386186 603654
rect 386422 603418 386604 603654
rect 386004 603334 386604 603418
rect 386004 603098 386186 603334
rect 386422 603098 386604 603334
rect 386004 567654 386604 603098
rect 386004 567418 386186 567654
rect 386422 567418 386604 567654
rect 386004 567334 386604 567418
rect 386004 567098 386186 567334
rect 386422 567098 386604 567334
rect 386004 531654 386604 567098
rect 386004 531418 386186 531654
rect 386422 531418 386604 531654
rect 386004 531334 386604 531418
rect 386004 531098 386186 531334
rect 386422 531098 386604 531334
rect 386004 495654 386604 531098
rect 386004 495418 386186 495654
rect 386422 495418 386604 495654
rect 386004 495334 386604 495418
rect 386004 495098 386186 495334
rect 386422 495098 386604 495334
rect 384987 486300 385053 486301
rect 384987 486236 384988 486300
rect 385052 486236 385053 486300
rect 384987 486235 385053 486236
rect 384990 486029 385050 486235
rect 384987 486028 385053 486029
rect 384987 485964 384988 486028
rect 385052 485964 385053 486028
rect 384987 485963 385053 485964
rect 382404 455818 382586 456054
rect 382822 455818 383004 456054
rect 382404 455734 383004 455818
rect 382404 455498 382586 455734
rect 382822 455498 383004 455734
rect 382404 420054 383004 455498
rect 382404 419818 382586 420054
rect 382822 419818 383004 420054
rect 382404 419734 383004 419818
rect 382404 419498 382586 419734
rect 382822 419498 383004 419734
rect 382404 384054 383004 419498
rect 382404 383818 382586 384054
rect 382822 383818 383004 384054
rect 382404 383734 383004 383818
rect 382404 383498 382586 383734
rect 382822 383498 383004 383734
rect 382404 348054 383004 383498
rect 382404 347818 382586 348054
rect 382822 347818 383004 348054
rect 382404 347734 383004 347818
rect 382404 347498 382586 347734
rect 382822 347498 383004 347734
rect 382404 312054 383004 347498
rect 382404 311818 382586 312054
rect 382822 311818 383004 312054
rect 382404 311734 383004 311818
rect 382404 311498 382586 311734
rect 382822 311498 383004 311734
rect 382404 276054 383004 311498
rect 382404 275818 382586 276054
rect 382822 275818 383004 276054
rect 382404 275734 383004 275818
rect 382404 275498 382586 275734
rect 382822 275498 383004 275734
rect 382404 240054 383004 275498
rect 382404 239818 382586 240054
rect 382822 239818 383004 240054
rect 382404 239734 383004 239818
rect 382404 239498 382586 239734
rect 382822 239498 383004 239734
rect 382404 204054 383004 239498
rect 382404 203818 382586 204054
rect 382822 203818 383004 204054
rect 382404 203734 383004 203818
rect 382404 203498 382586 203734
rect 382822 203498 383004 203734
rect 382404 168054 383004 203498
rect 382404 167818 382586 168054
rect 382822 167818 383004 168054
rect 382404 167734 383004 167818
rect 382404 167498 382586 167734
rect 382822 167498 383004 167734
rect 382404 132054 383004 167498
rect 382404 131818 382586 132054
rect 382822 131818 383004 132054
rect 382404 131734 383004 131818
rect 382404 131498 382586 131734
rect 382822 131498 383004 131734
rect 382404 96054 383004 131498
rect 382404 95818 382586 96054
rect 382822 95818 383004 96054
rect 382404 95734 383004 95818
rect 382404 95498 382586 95734
rect 382822 95498 383004 95734
rect 382404 60054 383004 95498
rect 382404 59818 382586 60054
rect 382822 59818 383004 60054
rect 382404 59734 383004 59818
rect 382404 59498 382586 59734
rect 382822 59498 383004 59734
rect 382404 24054 383004 59498
rect 386004 459654 386604 495098
rect 386004 459418 386186 459654
rect 386422 459418 386604 459654
rect 386004 459334 386604 459418
rect 386004 459098 386186 459334
rect 386422 459098 386604 459334
rect 386004 423654 386604 459098
rect 386004 423418 386186 423654
rect 386422 423418 386604 423654
rect 386004 423334 386604 423418
rect 386004 423098 386186 423334
rect 386422 423098 386604 423334
rect 386004 387654 386604 423098
rect 386004 387418 386186 387654
rect 386422 387418 386604 387654
rect 386004 387334 386604 387418
rect 386004 387098 386186 387334
rect 386422 387098 386604 387334
rect 386004 351654 386604 387098
rect 386004 351418 386186 351654
rect 386422 351418 386604 351654
rect 386004 351334 386604 351418
rect 386004 351098 386186 351334
rect 386422 351098 386604 351334
rect 386004 315654 386604 351098
rect 386004 315418 386186 315654
rect 386422 315418 386604 315654
rect 386004 315334 386604 315418
rect 386004 315098 386186 315334
rect 386422 315098 386604 315334
rect 386004 279654 386604 315098
rect 386004 279418 386186 279654
rect 386422 279418 386604 279654
rect 386004 279334 386604 279418
rect 386004 279098 386186 279334
rect 386422 279098 386604 279334
rect 386004 243654 386604 279098
rect 386004 243418 386186 243654
rect 386422 243418 386604 243654
rect 386004 243334 386604 243418
rect 386004 243098 386186 243334
rect 386422 243098 386604 243334
rect 386004 207654 386604 243098
rect 386004 207418 386186 207654
rect 386422 207418 386604 207654
rect 386004 207334 386604 207418
rect 386004 207098 386186 207334
rect 386422 207098 386604 207334
rect 386004 171654 386604 207098
rect 386004 171418 386186 171654
rect 386422 171418 386604 171654
rect 386004 171334 386604 171418
rect 386004 171098 386186 171334
rect 386422 171098 386604 171334
rect 386004 135654 386604 171098
rect 386004 135418 386186 135654
rect 386422 135418 386604 135654
rect 386004 135334 386604 135418
rect 386004 135098 386186 135334
rect 386422 135098 386604 135334
rect 386004 99654 386604 135098
rect 386004 99418 386186 99654
rect 386422 99418 386604 99654
rect 386004 99334 386604 99418
rect 386004 99098 386186 99334
rect 386422 99098 386604 99334
rect 386004 63654 386604 99098
rect 386004 63418 386186 63654
rect 386422 63418 386604 63654
rect 386004 63334 386604 63418
rect 386004 63098 386186 63334
rect 386422 63098 386604 63334
rect 384987 40492 385053 40493
rect 384987 40428 384988 40492
rect 385052 40428 385053 40492
rect 384987 40427 385053 40428
rect 384990 40221 385050 40427
rect 384987 40220 385053 40221
rect 384987 40156 384988 40220
rect 385052 40156 385053 40220
rect 384987 40155 385053 40156
rect 382404 23818 382586 24054
rect 382822 23818 383004 24054
rect 382404 23734 383004 23818
rect 382404 23498 382586 23734
rect 382822 23498 383004 23734
rect 382404 -3106 383004 23498
rect 382404 -3342 382586 -3106
rect 382822 -3342 383004 -3106
rect 382404 -3426 383004 -3342
rect 382404 -3662 382586 -3426
rect 382822 -3662 383004 -3426
rect 382404 -3684 383004 -3662
rect 386004 27654 386604 63098
rect 386004 27418 386186 27654
rect 386422 27418 386604 27654
rect 386004 27334 386604 27418
rect 386004 27098 386186 27334
rect 386422 27098 386604 27334
rect 386004 -4946 386604 27098
rect 386004 -5182 386186 -4946
rect 386422 -5182 386604 -4946
rect 386004 -5266 386604 -5182
rect 386004 -5502 386186 -5266
rect 386422 -5502 386604 -5266
rect 386004 -5524 386604 -5502
rect 389604 679254 390204 710722
rect 407604 710358 408204 711300
rect 407604 710122 407786 710358
rect 408022 710122 408204 710358
rect 407604 710038 408204 710122
rect 407604 709802 407786 710038
rect 408022 709802 408204 710038
rect 404004 708518 404604 709460
rect 404004 708282 404186 708518
rect 404422 708282 404604 708518
rect 404004 708198 404604 708282
rect 404004 707962 404186 708198
rect 404422 707962 404604 708198
rect 400404 706678 401004 707620
rect 400404 706442 400586 706678
rect 400822 706442 401004 706678
rect 400404 706358 401004 706442
rect 400404 706122 400586 706358
rect 400822 706122 401004 706358
rect 389604 679018 389786 679254
rect 390022 679018 390204 679254
rect 389604 678934 390204 679018
rect 389604 678698 389786 678934
rect 390022 678698 390204 678934
rect 389604 643254 390204 678698
rect 389604 643018 389786 643254
rect 390022 643018 390204 643254
rect 389604 642934 390204 643018
rect 389604 642698 389786 642934
rect 390022 642698 390204 642934
rect 389604 607254 390204 642698
rect 389604 607018 389786 607254
rect 390022 607018 390204 607254
rect 389604 606934 390204 607018
rect 389604 606698 389786 606934
rect 390022 606698 390204 606934
rect 389604 571254 390204 606698
rect 389604 571018 389786 571254
rect 390022 571018 390204 571254
rect 389604 570934 390204 571018
rect 389604 570698 389786 570934
rect 390022 570698 390204 570934
rect 389604 535254 390204 570698
rect 389604 535018 389786 535254
rect 390022 535018 390204 535254
rect 389604 534934 390204 535018
rect 389604 534698 389786 534934
rect 390022 534698 390204 534934
rect 389604 499254 390204 534698
rect 389604 499018 389786 499254
rect 390022 499018 390204 499254
rect 389604 498934 390204 499018
rect 389604 498698 389786 498934
rect 390022 498698 390204 498934
rect 389604 463254 390204 498698
rect 389604 463018 389786 463254
rect 390022 463018 390204 463254
rect 389604 462934 390204 463018
rect 389604 462698 389786 462934
rect 390022 462698 390204 462934
rect 389604 427254 390204 462698
rect 389604 427018 389786 427254
rect 390022 427018 390204 427254
rect 389604 426934 390204 427018
rect 389604 426698 389786 426934
rect 390022 426698 390204 426934
rect 389604 391254 390204 426698
rect 389604 391018 389786 391254
rect 390022 391018 390204 391254
rect 389604 390934 390204 391018
rect 389604 390698 389786 390934
rect 390022 390698 390204 390934
rect 389604 355254 390204 390698
rect 389604 355018 389786 355254
rect 390022 355018 390204 355254
rect 389604 354934 390204 355018
rect 389604 354698 389786 354934
rect 390022 354698 390204 354934
rect 389604 319254 390204 354698
rect 389604 319018 389786 319254
rect 390022 319018 390204 319254
rect 389604 318934 390204 319018
rect 389604 318698 389786 318934
rect 390022 318698 390204 318934
rect 389604 283254 390204 318698
rect 389604 283018 389786 283254
rect 390022 283018 390204 283254
rect 389604 282934 390204 283018
rect 389604 282698 389786 282934
rect 390022 282698 390204 282934
rect 389604 247254 390204 282698
rect 389604 247018 389786 247254
rect 390022 247018 390204 247254
rect 389604 246934 390204 247018
rect 389604 246698 389786 246934
rect 390022 246698 390204 246934
rect 389604 211254 390204 246698
rect 389604 211018 389786 211254
rect 390022 211018 390204 211254
rect 389604 210934 390204 211018
rect 389604 210698 389786 210934
rect 390022 210698 390204 210934
rect 389604 175254 390204 210698
rect 389604 175018 389786 175254
rect 390022 175018 390204 175254
rect 389604 174934 390204 175018
rect 389604 174698 389786 174934
rect 390022 174698 390204 174934
rect 389604 139254 390204 174698
rect 389604 139018 389786 139254
rect 390022 139018 390204 139254
rect 389604 138934 390204 139018
rect 389604 138698 389786 138934
rect 390022 138698 390204 138934
rect 389604 103254 390204 138698
rect 389604 103018 389786 103254
rect 390022 103018 390204 103254
rect 389604 102934 390204 103018
rect 389604 102698 389786 102934
rect 390022 102698 390204 102934
rect 389604 67254 390204 102698
rect 389604 67018 389786 67254
rect 390022 67018 390204 67254
rect 389604 66934 390204 67018
rect 389604 66698 389786 66934
rect 390022 66698 390204 66934
rect 389604 31254 390204 66698
rect 389604 31018 389786 31254
rect 390022 31018 390204 31254
rect 389604 30934 390204 31018
rect 389604 30698 389786 30934
rect 390022 30698 390204 30934
rect 371604 -6102 371786 -5866
rect 372022 -6102 372204 -5866
rect 371604 -6186 372204 -6102
rect 371604 -6422 371786 -6186
rect 372022 -6422 372204 -6186
rect 371604 -7364 372204 -6422
rect 389604 -6786 390204 30698
rect 396804 704838 397404 705780
rect 396804 704602 396986 704838
rect 397222 704602 397404 704838
rect 396804 704518 397404 704602
rect 396804 704282 396986 704518
rect 397222 704282 397404 704518
rect 396804 686454 397404 704282
rect 396804 686218 396986 686454
rect 397222 686218 397404 686454
rect 396804 686134 397404 686218
rect 396804 685898 396986 686134
rect 397222 685898 397404 686134
rect 396804 650454 397404 685898
rect 396804 650218 396986 650454
rect 397222 650218 397404 650454
rect 396804 650134 397404 650218
rect 396804 649898 396986 650134
rect 397222 649898 397404 650134
rect 396804 614454 397404 649898
rect 396804 614218 396986 614454
rect 397222 614218 397404 614454
rect 396804 614134 397404 614218
rect 396804 613898 396986 614134
rect 397222 613898 397404 614134
rect 396804 578454 397404 613898
rect 396804 578218 396986 578454
rect 397222 578218 397404 578454
rect 396804 578134 397404 578218
rect 396804 577898 396986 578134
rect 397222 577898 397404 578134
rect 396804 542454 397404 577898
rect 396804 542218 396986 542454
rect 397222 542218 397404 542454
rect 396804 542134 397404 542218
rect 396804 541898 396986 542134
rect 397222 541898 397404 542134
rect 396804 506454 397404 541898
rect 396804 506218 396986 506454
rect 397222 506218 397404 506454
rect 396804 506134 397404 506218
rect 396804 505898 396986 506134
rect 397222 505898 397404 506134
rect 396804 470454 397404 505898
rect 396804 470218 396986 470454
rect 397222 470218 397404 470454
rect 396804 470134 397404 470218
rect 396804 469898 396986 470134
rect 397222 469898 397404 470134
rect 396804 434454 397404 469898
rect 396804 434218 396986 434454
rect 397222 434218 397404 434454
rect 396804 434134 397404 434218
rect 396804 433898 396986 434134
rect 397222 433898 397404 434134
rect 396804 398454 397404 433898
rect 396804 398218 396986 398454
rect 397222 398218 397404 398454
rect 396804 398134 397404 398218
rect 396804 397898 396986 398134
rect 397222 397898 397404 398134
rect 396804 362454 397404 397898
rect 396804 362218 396986 362454
rect 397222 362218 397404 362454
rect 396804 362134 397404 362218
rect 396804 361898 396986 362134
rect 397222 361898 397404 362134
rect 396804 326454 397404 361898
rect 396804 326218 396986 326454
rect 397222 326218 397404 326454
rect 396804 326134 397404 326218
rect 396804 325898 396986 326134
rect 397222 325898 397404 326134
rect 396804 290454 397404 325898
rect 396804 290218 396986 290454
rect 397222 290218 397404 290454
rect 396804 290134 397404 290218
rect 396804 289898 396986 290134
rect 397222 289898 397404 290134
rect 396804 254454 397404 289898
rect 396804 254218 396986 254454
rect 397222 254218 397404 254454
rect 396804 254134 397404 254218
rect 396804 253898 396986 254134
rect 397222 253898 397404 254134
rect 396804 218454 397404 253898
rect 396804 218218 396986 218454
rect 397222 218218 397404 218454
rect 396804 218134 397404 218218
rect 396804 217898 396986 218134
rect 397222 217898 397404 218134
rect 396804 182454 397404 217898
rect 396804 182218 396986 182454
rect 397222 182218 397404 182454
rect 396804 182134 397404 182218
rect 396804 181898 396986 182134
rect 397222 181898 397404 182134
rect 396804 146454 397404 181898
rect 396804 146218 396986 146454
rect 397222 146218 397404 146454
rect 396804 146134 397404 146218
rect 396804 145898 396986 146134
rect 397222 145898 397404 146134
rect 396804 110454 397404 145898
rect 396804 110218 396986 110454
rect 397222 110218 397404 110454
rect 396804 110134 397404 110218
rect 396804 109898 396986 110134
rect 397222 109898 397404 110134
rect 396804 74454 397404 109898
rect 396804 74218 396986 74454
rect 397222 74218 397404 74454
rect 396804 74134 397404 74218
rect 396804 73898 396986 74134
rect 397222 73898 397404 74134
rect 396804 38454 397404 73898
rect 396804 38218 396986 38454
rect 397222 38218 397404 38454
rect 396804 38134 397404 38218
rect 396804 37898 396986 38134
rect 397222 37898 397404 38134
rect 396804 2454 397404 37898
rect 396804 2218 396986 2454
rect 397222 2218 397404 2454
rect 396804 2134 397404 2218
rect 396804 1898 396986 2134
rect 397222 1898 397404 2134
rect 396804 -346 397404 1898
rect 396804 -582 396986 -346
rect 397222 -582 397404 -346
rect 396804 -666 397404 -582
rect 396804 -902 396986 -666
rect 397222 -902 397404 -666
rect 396804 -1844 397404 -902
rect 400404 690054 401004 706122
rect 400404 689818 400586 690054
rect 400822 689818 401004 690054
rect 400404 689734 401004 689818
rect 400404 689498 400586 689734
rect 400822 689498 401004 689734
rect 400404 654054 401004 689498
rect 400404 653818 400586 654054
rect 400822 653818 401004 654054
rect 400404 653734 401004 653818
rect 400404 653498 400586 653734
rect 400822 653498 401004 653734
rect 400404 618054 401004 653498
rect 400404 617818 400586 618054
rect 400822 617818 401004 618054
rect 400404 617734 401004 617818
rect 400404 617498 400586 617734
rect 400822 617498 401004 617734
rect 400404 582054 401004 617498
rect 400404 581818 400586 582054
rect 400822 581818 401004 582054
rect 400404 581734 401004 581818
rect 400404 581498 400586 581734
rect 400822 581498 401004 581734
rect 400404 546054 401004 581498
rect 400404 545818 400586 546054
rect 400822 545818 401004 546054
rect 400404 545734 401004 545818
rect 400404 545498 400586 545734
rect 400822 545498 401004 545734
rect 400404 510054 401004 545498
rect 400404 509818 400586 510054
rect 400822 509818 401004 510054
rect 400404 509734 401004 509818
rect 400404 509498 400586 509734
rect 400822 509498 401004 509734
rect 400404 474054 401004 509498
rect 400404 473818 400586 474054
rect 400822 473818 401004 474054
rect 400404 473734 401004 473818
rect 400404 473498 400586 473734
rect 400822 473498 401004 473734
rect 400404 438054 401004 473498
rect 400404 437818 400586 438054
rect 400822 437818 401004 438054
rect 400404 437734 401004 437818
rect 400404 437498 400586 437734
rect 400822 437498 401004 437734
rect 400404 402054 401004 437498
rect 400404 401818 400586 402054
rect 400822 401818 401004 402054
rect 400404 401734 401004 401818
rect 400404 401498 400586 401734
rect 400822 401498 401004 401734
rect 400404 366054 401004 401498
rect 400404 365818 400586 366054
rect 400822 365818 401004 366054
rect 400404 365734 401004 365818
rect 400404 365498 400586 365734
rect 400822 365498 401004 365734
rect 400404 330054 401004 365498
rect 400404 329818 400586 330054
rect 400822 329818 401004 330054
rect 400404 329734 401004 329818
rect 400404 329498 400586 329734
rect 400822 329498 401004 329734
rect 400404 294054 401004 329498
rect 400404 293818 400586 294054
rect 400822 293818 401004 294054
rect 400404 293734 401004 293818
rect 400404 293498 400586 293734
rect 400822 293498 401004 293734
rect 400404 258054 401004 293498
rect 400404 257818 400586 258054
rect 400822 257818 401004 258054
rect 400404 257734 401004 257818
rect 400404 257498 400586 257734
rect 400822 257498 401004 257734
rect 400404 222054 401004 257498
rect 400404 221818 400586 222054
rect 400822 221818 401004 222054
rect 400404 221734 401004 221818
rect 400404 221498 400586 221734
rect 400822 221498 401004 221734
rect 400404 186054 401004 221498
rect 400404 185818 400586 186054
rect 400822 185818 401004 186054
rect 400404 185734 401004 185818
rect 400404 185498 400586 185734
rect 400822 185498 401004 185734
rect 400404 150054 401004 185498
rect 400404 149818 400586 150054
rect 400822 149818 401004 150054
rect 400404 149734 401004 149818
rect 400404 149498 400586 149734
rect 400822 149498 401004 149734
rect 400404 114054 401004 149498
rect 400404 113818 400586 114054
rect 400822 113818 401004 114054
rect 400404 113734 401004 113818
rect 400404 113498 400586 113734
rect 400822 113498 401004 113734
rect 400404 78054 401004 113498
rect 400404 77818 400586 78054
rect 400822 77818 401004 78054
rect 400404 77734 401004 77818
rect 400404 77498 400586 77734
rect 400822 77498 401004 77734
rect 400404 42054 401004 77498
rect 400404 41818 400586 42054
rect 400822 41818 401004 42054
rect 400404 41734 401004 41818
rect 400404 41498 400586 41734
rect 400822 41498 401004 41734
rect 400404 6054 401004 41498
rect 400404 5818 400586 6054
rect 400822 5818 401004 6054
rect 400404 5734 401004 5818
rect 400404 5498 400586 5734
rect 400822 5498 401004 5734
rect 400404 -2186 401004 5498
rect 400404 -2422 400586 -2186
rect 400822 -2422 401004 -2186
rect 400404 -2506 401004 -2422
rect 400404 -2742 400586 -2506
rect 400822 -2742 401004 -2506
rect 400404 -3684 401004 -2742
rect 404004 693654 404604 707962
rect 404004 693418 404186 693654
rect 404422 693418 404604 693654
rect 404004 693334 404604 693418
rect 404004 693098 404186 693334
rect 404422 693098 404604 693334
rect 404004 657654 404604 693098
rect 404004 657418 404186 657654
rect 404422 657418 404604 657654
rect 404004 657334 404604 657418
rect 404004 657098 404186 657334
rect 404422 657098 404604 657334
rect 404004 621654 404604 657098
rect 404004 621418 404186 621654
rect 404422 621418 404604 621654
rect 404004 621334 404604 621418
rect 404004 621098 404186 621334
rect 404422 621098 404604 621334
rect 404004 585654 404604 621098
rect 404004 585418 404186 585654
rect 404422 585418 404604 585654
rect 404004 585334 404604 585418
rect 404004 585098 404186 585334
rect 404422 585098 404604 585334
rect 404004 549654 404604 585098
rect 404004 549418 404186 549654
rect 404422 549418 404604 549654
rect 404004 549334 404604 549418
rect 404004 549098 404186 549334
rect 404422 549098 404604 549334
rect 404004 513654 404604 549098
rect 404004 513418 404186 513654
rect 404422 513418 404604 513654
rect 404004 513334 404604 513418
rect 404004 513098 404186 513334
rect 404422 513098 404604 513334
rect 404004 477654 404604 513098
rect 404004 477418 404186 477654
rect 404422 477418 404604 477654
rect 404004 477334 404604 477418
rect 404004 477098 404186 477334
rect 404422 477098 404604 477334
rect 404004 441654 404604 477098
rect 404004 441418 404186 441654
rect 404422 441418 404604 441654
rect 404004 441334 404604 441418
rect 404004 441098 404186 441334
rect 404422 441098 404604 441334
rect 404004 405654 404604 441098
rect 404004 405418 404186 405654
rect 404422 405418 404604 405654
rect 404004 405334 404604 405418
rect 404004 405098 404186 405334
rect 404422 405098 404604 405334
rect 404004 369654 404604 405098
rect 404004 369418 404186 369654
rect 404422 369418 404604 369654
rect 404004 369334 404604 369418
rect 404004 369098 404186 369334
rect 404422 369098 404604 369334
rect 404004 333654 404604 369098
rect 404004 333418 404186 333654
rect 404422 333418 404604 333654
rect 404004 333334 404604 333418
rect 404004 333098 404186 333334
rect 404422 333098 404604 333334
rect 404004 297654 404604 333098
rect 404004 297418 404186 297654
rect 404422 297418 404604 297654
rect 404004 297334 404604 297418
rect 404004 297098 404186 297334
rect 404422 297098 404604 297334
rect 404004 261654 404604 297098
rect 404004 261418 404186 261654
rect 404422 261418 404604 261654
rect 404004 261334 404604 261418
rect 404004 261098 404186 261334
rect 404422 261098 404604 261334
rect 404004 225654 404604 261098
rect 404004 225418 404186 225654
rect 404422 225418 404604 225654
rect 404004 225334 404604 225418
rect 404004 225098 404186 225334
rect 404422 225098 404604 225334
rect 404004 189654 404604 225098
rect 404004 189418 404186 189654
rect 404422 189418 404604 189654
rect 404004 189334 404604 189418
rect 404004 189098 404186 189334
rect 404422 189098 404604 189334
rect 404004 153654 404604 189098
rect 404004 153418 404186 153654
rect 404422 153418 404604 153654
rect 404004 153334 404604 153418
rect 404004 153098 404186 153334
rect 404422 153098 404604 153334
rect 404004 117654 404604 153098
rect 404004 117418 404186 117654
rect 404422 117418 404604 117654
rect 404004 117334 404604 117418
rect 404004 117098 404186 117334
rect 404422 117098 404604 117334
rect 404004 81654 404604 117098
rect 404004 81418 404186 81654
rect 404422 81418 404604 81654
rect 404004 81334 404604 81418
rect 404004 81098 404186 81334
rect 404422 81098 404604 81334
rect 404004 45654 404604 81098
rect 404004 45418 404186 45654
rect 404422 45418 404604 45654
rect 404004 45334 404604 45418
rect 404004 45098 404186 45334
rect 404422 45098 404604 45334
rect 404004 9654 404604 45098
rect 404004 9418 404186 9654
rect 404422 9418 404604 9654
rect 404004 9334 404604 9418
rect 404004 9098 404186 9334
rect 404422 9098 404604 9334
rect 404004 -4026 404604 9098
rect 404004 -4262 404186 -4026
rect 404422 -4262 404604 -4026
rect 404004 -4346 404604 -4262
rect 404004 -4582 404186 -4346
rect 404422 -4582 404604 -4346
rect 404004 -5524 404604 -4582
rect 407604 697254 408204 709802
rect 425604 711278 426204 711300
rect 425604 711042 425786 711278
rect 426022 711042 426204 711278
rect 425604 710958 426204 711042
rect 425604 710722 425786 710958
rect 426022 710722 426204 710958
rect 422004 709438 422604 709460
rect 422004 709202 422186 709438
rect 422422 709202 422604 709438
rect 422004 709118 422604 709202
rect 422004 708882 422186 709118
rect 422422 708882 422604 709118
rect 418404 707598 419004 707620
rect 418404 707362 418586 707598
rect 418822 707362 419004 707598
rect 418404 707278 419004 707362
rect 418404 707042 418586 707278
rect 418822 707042 419004 707278
rect 407604 697018 407786 697254
rect 408022 697018 408204 697254
rect 407604 696934 408204 697018
rect 407604 696698 407786 696934
rect 408022 696698 408204 696934
rect 407604 661254 408204 696698
rect 407604 661018 407786 661254
rect 408022 661018 408204 661254
rect 407604 660934 408204 661018
rect 407604 660698 407786 660934
rect 408022 660698 408204 660934
rect 407604 625254 408204 660698
rect 407604 625018 407786 625254
rect 408022 625018 408204 625254
rect 407604 624934 408204 625018
rect 407604 624698 407786 624934
rect 408022 624698 408204 624934
rect 407604 589254 408204 624698
rect 407604 589018 407786 589254
rect 408022 589018 408204 589254
rect 407604 588934 408204 589018
rect 407604 588698 407786 588934
rect 408022 588698 408204 588934
rect 407604 553254 408204 588698
rect 407604 553018 407786 553254
rect 408022 553018 408204 553254
rect 407604 552934 408204 553018
rect 407604 552698 407786 552934
rect 408022 552698 408204 552934
rect 407604 517254 408204 552698
rect 407604 517018 407786 517254
rect 408022 517018 408204 517254
rect 407604 516934 408204 517018
rect 407604 516698 407786 516934
rect 408022 516698 408204 516934
rect 407604 481254 408204 516698
rect 407604 481018 407786 481254
rect 408022 481018 408204 481254
rect 407604 480934 408204 481018
rect 407604 480698 407786 480934
rect 408022 480698 408204 480934
rect 407604 445254 408204 480698
rect 407604 445018 407786 445254
rect 408022 445018 408204 445254
rect 407604 444934 408204 445018
rect 407604 444698 407786 444934
rect 408022 444698 408204 444934
rect 407604 409254 408204 444698
rect 407604 409018 407786 409254
rect 408022 409018 408204 409254
rect 407604 408934 408204 409018
rect 407604 408698 407786 408934
rect 408022 408698 408204 408934
rect 407604 373254 408204 408698
rect 407604 373018 407786 373254
rect 408022 373018 408204 373254
rect 407604 372934 408204 373018
rect 407604 372698 407786 372934
rect 408022 372698 408204 372934
rect 407604 337254 408204 372698
rect 407604 337018 407786 337254
rect 408022 337018 408204 337254
rect 407604 336934 408204 337018
rect 407604 336698 407786 336934
rect 408022 336698 408204 336934
rect 407604 301254 408204 336698
rect 407604 301018 407786 301254
rect 408022 301018 408204 301254
rect 407604 300934 408204 301018
rect 407604 300698 407786 300934
rect 408022 300698 408204 300934
rect 407604 265254 408204 300698
rect 407604 265018 407786 265254
rect 408022 265018 408204 265254
rect 407604 264934 408204 265018
rect 407604 264698 407786 264934
rect 408022 264698 408204 264934
rect 407604 229254 408204 264698
rect 407604 229018 407786 229254
rect 408022 229018 408204 229254
rect 407604 228934 408204 229018
rect 407604 228698 407786 228934
rect 408022 228698 408204 228934
rect 407604 193254 408204 228698
rect 407604 193018 407786 193254
rect 408022 193018 408204 193254
rect 407604 192934 408204 193018
rect 407604 192698 407786 192934
rect 408022 192698 408204 192934
rect 407604 157254 408204 192698
rect 407604 157018 407786 157254
rect 408022 157018 408204 157254
rect 407604 156934 408204 157018
rect 407604 156698 407786 156934
rect 408022 156698 408204 156934
rect 407604 121254 408204 156698
rect 407604 121018 407786 121254
rect 408022 121018 408204 121254
rect 407604 120934 408204 121018
rect 407604 120698 407786 120934
rect 408022 120698 408204 120934
rect 407604 85254 408204 120698
rect 407604 85018 407786 85254
rect 408022 85018 408204 85254
rect 407604 84934 408204 85018
rect 407604 84698 407786 84934
rect 408022 84698 408204 84934
rect 407604 49254 408204 84698
rect 407604 49018 407786 49254
rect 408022 49018 408204 49254
rect 407604 48934 408204 49018
rect 407604 48698 407786 48934
rect 408022 48698 408204 48934
rect 407604 13254 408204 48698
rect 407604 13018 407786 13254
rect 408022 13018 408204 13254
rect 407604 12934 408204 13018
rect 407604 12698 407786 12934
rect 408022 12698 408204 12934
rect 389604 -7022 389786 -6786
rect 390022 -7022 390204 -6786
rect 389604 -7106 390204 -7022
rect 389604 -7342 389786 -7106
rect 390022 -7342 390204 -7106
rect 389604 -7364 390204 -7342
rect 407604 -5866 408204 12698
rect 414804 705758 415404 705780
rect 414804 705522 414986 705758
rect 415222 705522 415404 705758
rect 414804 705438 415404 705522
rect 414804 705202 414986 705438
rect 415222 705202 415404 705438
rect 414804 668454 415404 705202
rect 414804 668218 414986 668454
rect 415222 668218 415404 668454
rect 414804 668134 415404 668218
rect 414804 667898 414986 668134
rect 415222 667898 415404 668134
rect 414804 632454 415404 667898
rect 414804 632218 414986 632454
rect 415222 632218 415404 632454
rect 414804 632134 415404 632218
rect 414804 631898 414986 632134
rect 415222 631898 415404 632134
rect 414804 596454 415404 631898
rect 414804 596218 414986 596454
rect 415222 596218 415404 596454
rect 414804 596134 415404 596218
rect 414804 595898 414986 596134
rect 415222 595898 415404 596134
rect 414804 560454 415404 595898
rect 414804 560218 414986 560454
rect 415222 560218 415404 560454
rect 414804 560134 415404 560218
rect 414804 559898 414986 560134
rect 415222 559898 415404 560134
rect 414804 524454 415404 559898
rect 414804 524218 414986 524454
rect 415222 524218 415404 524454
rect 414804 524134 415404 524218
rect 414804 523898 414986 524134
rect 415222 523898 415404 524134
rect 414804 488454 415404 523898
rect 414804 488218 414986 488454
rect 415222 488218 415404 488454
rect 414804 488134 415404 488218
rect 414804 487898 414986 488134
rect 415222 487898 415404 488134
rect 414804 452454 415404 487898
rect 414804 452218 414986 452454
rect 415222 452218 415404 452454
rect 414804 452134 415404 452218
rect 414804 451898 414986 452134
rect 415222 451898 415404 452134
rect 414804 416454 415404 451898
rect 414804 416218 414986 416454
rect 415222 416218 415404 416454
rect 414804 416134 415404 416218
rect 414804 415898 414986 416134
rect 415222 415898 415404 416134
rect 414804 380454 415404 415898
rect 414804 380218 414986 380454
rect 415222 380218 415404 380454
rect 414804 380134 415404 380218
rect 414804 379898 414986 380134
rect 415222 379898 415404 380134
rect 414804 344454 415404 379898
rect 414804 344218 414986 344454
rect 415222 344218 415404 344454
rect 414804 344134 415404 344218
rect 414804 343898 414986 344134
rect 415222 343898 415404 344134
rect 414804 308454 415404 343898
rect 414804 308218 414986 308454
rect 415222 308218 415404 308454
rect 414804 308134 415404 308218
rect 414804 307898 414986 308134
rect 415222 307898 415404 308134
rect 414804 272454 415404 307898
rect 414804 272218 414986 272454
rect 415222 272218 415404 272454
rect 414804 272134 415404 272218
rect 414804 271898 414986 272134
rect 415222 271898 415404 272134
rect 414804 236454 415404 271898
rect 414804 236218 414986 236454
rect 415222 236218 415404 236454
rect 414804 236134 415404 236218
rect 414804 235898 414986 236134
rect 415222 235898 415404 236134
rect 414804 200454 415404 235898
rect 414804 200218 414986 200454
rect 415222 200218 415404 200454
rect 414804 200134 415404 200218
rect 414804 199898 414986 200134
rect 415222 199898 415404 200134
rect 414804 164454 415404 199898
rect 414804 164218 414986 164454
rect 415222 164218 415404 164454
rect 414804 164134 415404 164218
rect 414804 163898 414986 164134
rect 415222 163898 415404 164134
rect 414804 128454 415404 163898
rect 414804 128218 414986 128454
rect 415222 128218 415404 128454
rect 414804 128134 415404 128218
rect 414804 127898 414986 128134
rect 415222 127898 415404 128134
rect 414804 92454 415404 127898
rect 414804 92218 414986 92454
rect 415222 92218 415404 92454
rect 414804 92134 415404 92218
rect 414804 91898 414986 92134
rect 415222 91898 415404 92134
rect 414804 56454 415404 91898
rect 414804 56218 414986 56454
rect 415222 56218 415404 56454
rect 414804 56134 415404 56218
rect 414804 55898 414986 56134
rect 415222 55898 415404 56134
rect 414804 20454 415404 55898
rect 414804 20218 414986 20454
rect 415222 20218 415404 20454
rect 414804 20134 415404 20218
rect 414804 19898 414986 20134
rect 415222 19898 415404 20134
rect 414804 -1266 415404 19898
rect 414804 -1502 414986 -1266
rect 415222 -1502 415404 -1266
rect 414804 -1586 415404 -1502
rect 414804 -1822 414986 -1586
rect 415222 -1822 415404 -1586
rect 414804 -1844 415404 -1822
rect 418404 672054 419004 707042
rect 418404 671818 418586 672054
rect 418822 671818 419004 672054
rect 418404 671734 419004 671818
rect 418404 671498 418586 671734
rect 418822 671498 419004 671734
rect 418404 636054 419004 671498
rect 418404 635818 418586 636054
rect 418822 635818 419004 636054
rect 418404 635734 419004 635818
rect 418404 635498 418586 635734
rect 418822 635498 419004 635734
rect 418404 600054 419004 635498
rect 418404 599818 418586 600054
rect 418822 599818 419004 600054
rect 418404 599734 419004 599818
rect 418404 599498 418586 599734
rect 418822 599498 419004 599734
rect 418404 564054 419004 599498
rect 418404 563818 418586 564054
rect 418822 563818 419004 564054
rect 418404 563734 419004 563818
rect 418404 563498 418586 563734
rect 418822 563498 419004 563734
rect 418404 528054 419004 563498
rect 418404 527818 418586 528054
rect 418822 527818 419004 528054
rect 418404 527734 419004 527818
rect 418404 527498 418586 527734
rect 418822 527498 419004 527734
rect 418404 492054 419004 527498
rect 418404 491818 418586 492054
rect 418822 491818 419004 492054
rect 418404 491734 419004 491818
rect 418404 491498 418586 491734
rect 418822 491498 419004 491734
rect 418404 456054 419004 491498
rect 418404 455818 418586 456054
rect 418822 455818 419004 456054
rect 418404 455734 419004 455818
rect 418404 455498 418586 455734
rect 418822 455498 419004 455734
rect 418404 420054 419004 455498
rect 418404 419818 418586 420054
rect 418822 419818 419004 420054
rect 418404 419734 419004 419818
rect 418404 419498 418586 419734
rect 418822 419498 419004 419734
rect 418404 384054 419004 419498
rect 418404 383818 418586 384054
rect 418822 383818 419004 384054
rect 418404 383734 419004 383818
rect 418404 383498 418586 383734
rect 418822 383498 419004 383734
rect 418404 348054 419004 383498
rect 418404 347818 418586 348054
rect 418822 347818 419004 348054
rect 418404 347734 419004 347818
rect 418404 347498 418586 347734
rect 418822 347498 419004 347734
rect 418404 312054 419004 347498
rect 418404 311818 418586 312054
rect 418822 311818 419004 312054
rect 418404 311734 419004 311818
rect 418404 311498 418586 311734
rect 418822 311498 419004 311734
rect 418404 276054 419004 311498
rect 418404 275818 418586 276054
rect 418822 275818 419004 276054
rect 418404 275734 419004 275818
rect 418404 275498 418586 275734
rect 418822 275498 419004 275734
rect 418404 240054 419004 275498
rect 418404 239818 418586 240054
rect 418822 239818 419004 240054
rect 418404 239734 419004 239818
rect 418404 239498 418586 239734
rect 418822 239498 419004 239734
rect 418404 204054 419004 239498
rect 418404 203818 418586 204054
rect 418822 203818 419004 204054
rect 418404 203734 419004 203818
rect 418404 203498 418586 203734
rect 418822 203498 419004 203734
rect 418404 168054 419004 203498
rect 418404 167818 418586 168054
rect 418822 167818 419004 168054
rect 418404 167734 419004 167818
rect 418404 167498 418586 167734
rect 418822 167498 419004 167734
rect 418404 132054 419004 167498
rect 418404 131818 418586 132054
rect 418822 131818 419004 132054
rect 418404 131734 419004 131818
rect 418404 131498 418586 131734
rect 418822 131498 419004 131734
rect 418404 96054 419004 131498
rect 418404 95818 418586 96054
rect 418822 95818 419004 96054
rect 418404 95734 419004 95818
rect 418404 95498 418586 95734
rect 418822 95498 419004 95734
rect 418404 60054 419004 95498
rect 418404 59818 418586 60054
rect 418822 59818 419004 60054
rect 418404 59734 419004 59818
rect 418404 59498 418586 59734
rect 418822 59498 419004 59734
rect 418404 24054 419004 59498
rect 418404 23818 418586 24054
rect 418822 23818 419004 24054
rect 418404 23734 419004 23818
rect 418404 23498 418586 23734
rect 418822 23498 419004 23734
rect 418404 -3106 419004 23498
rect 418404 -3342 418586 -3106
rect 418822 -3342 419004 -3106
rect 418404 -3426 419004 -3342
rect 418404 -3662 418586 -3426
rect 418822 -3662 419004 -3426
rect 418404 -3684 419004 -3662
rect 422004 675654 422604 708882
rect 422004 675418 422186 675654
rect 422422 675418 422604 675654
rect 422004 675334 422604 675418
rect 422004 675098 422186 675334
rect 422422 675098 422604 675334
rect 422004 639654 422604 675098
rect 422004 639418 422186 639654
rect 422422 639418 422604 639654
rect 422004 639334 422604 639418
rect 422004 639098 422186 639334
rect 422422 639098 422604 639334
rect 422004 603654 422604 639098
rect 422004 603418 422186 603654
rect 422422 603418 422604 603654
rect 422004 603334 422604 603418
rect 422004 603098 422186 603334
rect 422422 603098 422604 603334
rect 422004 567654 422604 603098
rect 422004 567418 422186 567654
rect 422422 567418 422604 567654
rect 422004 567334 422604 567418
rect 422004 567098 422186 567334
rect 422422 567098 422604 567334
rect 422004 531654 422604 567098
rect 422004 531418 422186 531654
rect 422422 531418 422604 531654
rect 422004 531334 422604 531418
rect 422004 531098 422186 531334
rect 422422 531098 422604 531334
rect 422004 495654 422604 531098
rect 422004 495418 422186 495654
rect 422422 495418 422604 495654
rect 422004 495334 422604 495418
rect 422004 495098 422186 495334
rect 422422 495098 422604 495334
rect 422004 459654 422604 495098
rect 422004 459418 422186 459654
rect 422422 459418 422604 459654
rect 422004 459334 422604 459418
rect 422004 459098 422186 459334
rect 422422 459098 422604 459334
rect 422004 423654 422604 459098
rect 422004 423418 422186 423654
rect 422422 423418 422604 423654
rect 422004 423334 422604 423418
rect 422004 423098 422186 423334
rect 422422 423098 422604 423334
rect 422004 387654 422604 423098
rect 422004 387418 422186 387654
rect 422422 387418 422604 387654
rect 422004 387334 422604 387418
rect 422004 387098 422186 387334
rect 422422 387098 422604 387334
rect 422004 351654 422604 387098
rect 422004 351418 422186 351654
rect 422422 351418 422604 351654
rect 422004 351334 422604 351418
rect 422004 351098 422186 351334
rect 422422 351098 422604 351334
rect 422004 315654 422604 351098
rect 422004 315418 422186 315654
rect 422422 315418 422604 315654
rect 422004 315334 422604 315418
rect 422004 315098 422186 315334
rect 422422 315098 422604 315334
rect 422004 279654 422604 315098
rect 422004 279418 422186 279654
rect 422422 279418 422604 279654
rect 422004 279334 422604 279418
rect 422004 279098 422186 279334
rect 422422 279098 422604 279334
rect 422004 243654 422604 279098
rect 422004 243418 422186 243654
rect 422422 243418 422604 243654
rect 422004 243334 422604 243418
rect 422004 243098 422186 243334
rect 422422 243098 422604 243334
rect 422004 207654 422604 243098
rect 422004 207418 422186 207654
rect 422422 207418 422604 207654
rect 422004 207334 422604 207418
rect 422004 207098 422186 207334
rect 422422 207098 422604 207334
rect 422004 171654 422604 207098
rect 422004 171418 422186 171654
rect 422422 171418 422604 171654
rect 422004 171334 422604 171418
rect 422004 171098 422186 171334
rect 422422 171098 422604 171334
rect 422004 135654 422604 171098
rect 422004 135418 422186 135654
rect 422422 135418 422604 135654
rect 422004 135334 422604 135418
rect 422004 135098 422186 135334
rect 422422 135098 422604 135334
rect 422004 99654 422604 135098
rect 422004 99418 422186 99654
rect 422422 99418 422604 99654
rect 422004 99334 422604 99418
rect 422004 99098 422186 99334
rect 422422 99098 422604 99334
rect 422004 63654 422604 99098
rect 422004 63418 422186 63654
rect 422422 63418 422604 63654
rect 422004 63334 422604 63418
rect 422004 63098 422186 63334
rect 422422 63098 422604 63334
rect 422004 27654 422604 63098
rect 422004 27418 422186 27654
rect 422422 27418 422604 27654
rect 422004 27334 422604 27418
rect 422004 27098 422186 27334
rect 422422 27098 422604 27334
rect 422004 -4946 422604 27098
rect 422004 -5182 422186 -4946
rect 422422 -5182 422604 -4946
rect 422004 -5266 422604 -5182
rect 422004 -5502 422186 -5266
rect 422422 -5502 422604 -5266
rect 422004 -5524 422604 -5502
rect 425604 679254 426204 710722
rect 443604 710358 444204 711300
rect 443604 710122 443786 710358
rect 444022 710122 444204 710358
rect 443604 710038 444204 710122
rect 443604 709802 443786 710038
rect 444022 709802 444204 710038
rect 440004 708518 440604 709460
rect 440004 708282 440186 708518
rect 440422 708282 440604 708518
rect 440004 708198 440604 708282
rect 440004 707962 440186 708198
rect 440422 707962 440604 708198
rect 436404 706678 437004 707620
rect 436404 706442 436586 706678
rect 436822 706442 437004 706678
rect 436404 706358 437004 706442
rect 436404 706122 436586 706358
rect 436822 706122 437004 706358
rect 425604 679018 425786 679254
rect 426022 679018 426204 679254
rect 425604 678934 426204 679018
rect 425604 678698 425786 678934
rect 426022 678698 426204 678934
rect 425604 643254 426204 678698
rect 425604 643018 425786 643254
rect 426022 643018 426204 643254
rect 425604 642934 426204 643018
rect 425604 642698 425786 642934
rect 426022 642698 426204 642934
rect 425604 607254 426204 642698
rect 425604 607018 425786 607254
rect 426022 607018 426204 607254
rect 425604 606934 426204 607018
rect 425604 606698 425786 606934
rect 426022 606698 426204 606934
rect 425604 571254 426204 606698
rect 425604 571018 425786 571254
rect 426022 571018 426204 571254
rect 425604 570934 426204 571018
rect 425604 570698 425786 570934
rect 426022 570698 426204 570934
rect 425604 535254 426204 570698
rect 425604 535018 425786 535254
rect 426022 535018 426204 535254
rect 425604 534934 426204 535018
rect 425604 534698 425786 534934
rect 426022 534698 426204 534934
rect 425604 499254 426204 534698
rect 425604 499018 425786 499254
rect 426022 499018 426204 499254
rect 425604 498934 426204 499018
rect 425604 498698 425786 498934
rect 426022 498698 426204 498934
rect 425604 463254 426204 498698
rect 425604 463018 425786 463254
rect 426022 463018 426204 463254
rect 425604 462934 426204 463018
rect 425604 462698 425786 462934
rect 426022 462698 426204 462934
rect 425604 427254 426204 462698
rect 425604 427018 425786 427254
rect 426022 427018 426204 427254
rect 425604 426934 426204 427018
rect 425604 426698 425786 426934
rect 426022 426698 426204 426934
rect 425604 391254 426204 426698
rect 425604 391018 425786 391254
rect 426022 391018 426204 391254
rect 425604 390934 426204 391018
rect 425604 390698 425786 390934
rect 426022 390698 426204 390934
rect 425604 355254 426204 390698
rect 425604 355018 425786 355254
rect 426022 355018 426204 355254
rect 425604 354934 426204 355018
rect 425604 354698 425786 354934
rect 426022 354698 426204 354934
rect 425604 319254 426204 354698
rect 425604 319018 425786 319254
rect 426022 319018 426204 319254
rect 425604 318934 426204 319018
rect 425604 318698 425786 318934
rect 426022 318698 426204 318934
rect 425604 283254 426204 318698
rect 425604 283018 425786 283254
rect 426022 283018 426204 283254
rect 425604 282934 426204 283018
rect 425604 282698 425786 282934
rect 426022 282698 426204 282934
rect 425604 247254 426204 282698
rect 425604 247018 425786 247254
rect 426022 247018 426204 247254
rect 425604 246934 426204 247018
rect 425604 246698 425786 246934
rect 426022 246698 426204 246934
rect 425604 211254 426204 246698
rect 425604 211018 425786 211254
rect 426022 211018 426204 211254
rect 425604 210934 426204 211018
rect 425604 210698 425786 210934
rect 426022 210698 426204 210934
rect 425604 175254 426204 210698
rect 425604 175018 425786 175254
rect 426022 175018 426204 175254
rect 425604 174934 426204 175018
rect 425604 174698 425786 174934
rect 426022 174698 426204 174934
rect 425604 139254 426204 174698
rect 425604 139018 425786 139254
rect 426022 139018 426204 139254
rect 425604 138934 426204 139018
rect 425604 138698 425786 138934
rect 426022 138698 426204 138934
rect 425604 103254 426204 138698
rect 425604 103018 425786 103254
rect 426022 103018 426204 103254
rect 425604 102934 426204 103018
rect 425604 102698 425786 102934
rect 426022 102698 426204 102934
rect 425604 67254 426204 102698
rect 425604 67018 425786 67254
rect 426022 67018 426204 67254
rect 425604 66934 426204 67018
rect 425604 66698 425786 66934
rect 426022 66698 426204 66934
rect 425604 31254 426204 66698
rect 425604 31018 425786 31254
rect 426022 31018 426204 31254
rect 425604 30934 426204 31018
rect 425604 30698 425786 30934
rect 426022 30698 426204 30934
rect 407604 -6102 407786 -5866
rect 408022 -6102 408204 -5866
rect 407604 -6186 408204 -6102
rect 407604 -6422 407786 -6186
rect 408022 -6422 408204 -6186
rect 407604 -7364 408204 -6422
rect 425604 -6786 426204 30698
rect 432804 704838 433404 705780
rect 432804 704602 432986 704838
rect 433222 704602 433404 704838
rect 432804 704518 433404 704602
rect 432804 704282 432986 704518
rect 433222 704282 433404 704518
rect 432804 686454 433404 704282
rect 432804 686218 432986 686454
rect 433222 686218 433404 686454
rect 432804 686134 433404 686218
rect 432804 685898 432986 686134
rect 433222 685898 433404 686134
rect 432804 650454 433404 685898
rect 432804 650218 432986 650454
rect 433222 650218 433404 650454
rect 432804 650134 433404 650218
rect 432804 649898 432986 650134
rect 433222 649898 433404 650134
rect 432804 614454 433404 649898
rect 432804 614218 432986 614454
rect 433222 614218 433404 614454
rect 432804 614134 433404 614218
rect 432804 613898 432986 614134
rect 433222 613898 433404 614134
rect 432804 578454 433404 613898
rect 432804 578218 432986 578454
rect 433222 578218 433404 578454
rect 432804 578134 433404 578218
rect 432804 577898 432986 578134
rect 433222 577898 433404 578134
rect 432804 542454 433404 577898
rect 432804 542218 432986 542454
rect 433222 542218 433404 542454
rect 432804 542134 433404 542218
rect 432804 541898 432986 542134
rect 433222 541898 433404 542134
rect 432804 506454 433404 541898
rect 432804 506218 432986 506454
rect 433222 506218 433404 506454
rect 432804 506134 433404 506218
rect 432804 505898 432986 506134
rect 433222 505898 433404 506134
rect 432804 470454 433404 505898
rect 432804 470218 432986 470454
rect 433222 470218 433404 470454
rect 432804 470134 433404 470218
rect 432804 469898 432986 470134
rect 433222 469898 433404 470134
rect 432804 434454 433404 469898
rect 432804 434218 432986 434454
rect 433222 434218 433404 434454
rect 432804 434134 433404 434218
rect 432804 433898 432986 434134
rect 433222 433898 433404 434134
rect 432804 398454 433404 433898
rect 432804 398218 432986 398454
rect 433222 398218 433404 398454
rect 432804 398134 433404 398218
rect 432804 397898 432986 398134
rect 433222 397898 433404 398134
rect 432804 362454 433404 397898
rect 432804 362218 432986 362454
rect 433222 362218 433404 362454
rect 432804 362134 433404 362218
rect 432804 361898 432986 362134
rect 433222 361898 433404 362134
rect 432804 326454 433404 361898
rect 432804 326218 432986 326454
rect 433222 326218 433404 326454
rect 432804 326134 433404 326218
rect 432804 325898 432986 326134
rect 433222 325898 433404 326134
rect 432804 290454 433404 325898
rect 432804 290218 432986 290454
rect 433222 290218 433404 290454
rect 432804 290134 433404 290218
rect 432804 289898 432986 290134
rect 433222 289898 433404 290134
rect 432804 254454 433404 289898
rect 432804 254218 432986 254454
rect 433222 254218 433404 254454
rect 432804 254134 433404 254218
rect 432804 253898 432986 254134
rect 433222 253898 433404 254134
rect 432804 218454 433404 253898
rect 432804 218218 432986 218454
rect 433222 218218 433404 218454
rect 432804 218134 433404 218218
rect 432804 217898 432986 218134
rect 433222 217898 433404 218134
rect 432804 182454 433404 217898
rect 432804 182218 432986 182454
rect 433222 182218 433404 182454
rect 432804 182134 433404 182218
rect 432804 181898 432986 182134
rect 433222 181898 433404 182134
rect 432804 146454 433404 181898
rect 432804 146218 432986 146454
rect 433222 146218 433404 146454
rect 432804 146134 433404 146218
rect 432804 145898 432986 146134
rect 433222 145898 433404 146134
rect 432804 110454 433404 145898
rect 432804 110218 432986 110454
rect 433222 110218 433404 110454
rect 432804 110134 433404 110218
rect 432804 109898 432986 110134
rect 433222 109898 433404 110134
rect 432804 74454 433404 109898
rect 432804 74218 432986 74454
rect 433222 74218 433404 74454
rect 432804 74134 433404 74218
rect 432804 73898 432986 74134
rect 433222 73898 433404 74134
rect 432804 38454 433404 73898
rect 432804 38218 432986 38454
rect 433222 38218 433404 38454
rect 432804 38134 433404 38218
rect 432804 37898 432986 38134
rect 433222 37898 433404 38134
rect 432804 2454 433404 37898
rect 432804 2218 432986 2454
rect 433222 2218 433404 2454
rect 432804 2134 433404 2218
rect 432804 1898 432986 2134
rect 433222 1898 433404 2134
rect 432804 -346 433404 1898
rect 432804 -582 432986 -346
rect 433222 -582 433404 -346
rect 432804 -666 433404 -582
rect 432804 -902 432986 -666
rect 433222 -902 433404 -666
rect 432804 -1844 433404 -902
rect 436404 690054 437004 706122
rect 436404 689818 436586 690054
rect 436822 689818 437004 690054
rect 436404 689734 437004 689818
rect 436404 689498 436586 689734
rect 436822 689498 437004 689734
rect 436404 654054 437004 689498
rect 436404 653818 436586 654054
rect 436822 653818 437004 654054
rect 436404 653734 437004 653818
rect 436404 653498 436586 653734
rect 436822 653498 437004 653734
rect 436404 618054 437004 653498
rect 436404 617818 436586 618054
rect 436822 617818 437004 618054
rect 436404 617734 437004 617818
rect 436404 617498 436586 617734
rect 436822 617498 437004 617734
rect 436404 582054 437004 617498
rect 436404 581818 436586 582054
rect 436822 581818 437004 582054
rect 436404 581734 437004 581818
rect 436404 581498 436586 581734
rect 436822 581498 437004 581734
rect 436404 546054 437004 581498
rect 436404 545818 436586 546054
rect 436822 545818 437004 546054
rect 436404 545734 437004 545818
rect 436404 545498 436586 545734
rect 436822 545498 437004 545734
rect 436404 510054 437004 545498
rect 436404 509818 436586 510054
rect 436822 509818 437004 510054
rect 436404 509734 437004 509818
rect 436404 509498 436586 509734
rect 436822 509498 437004 509734
rect 436404 474054 437004 509498
rect 436404 473818 436586 474054
rect 436822 473818 437004 474054
rect 436404 473734 437004 473818
rect 436404 473498 436586 473734
rect 436822 473498 437004 473734
rect 436404 438054 437004 473498
rect 436404 437818 436586 438054
rect 436822 437818 437004 438054
rect 436404 437734 437004 437818
rect 436404 437498 436586 437734
rect 436822 437498 437004 437734
rect 436404 402054 437004 437498
rect 436404 401818 436586 402054
rect 436822 401818 437004 402054
rect 436404 401734 437004 401818
rect 436404 401498 436586 401734
rect 436822 401498 437004 401734
rect 436404 366054 437004 401498
rect 436404 365818 436586 366054
rect 436822 365818 437004 366054
rect 436404 365734 437004 365818
rect 436404 365498 436586 365734
rect 436822 365498 437004 365734
rect 436404 330054 437004 365498
rect 436404 329818 436586 330054
rect 436822 329818 437004 330054
rect 436404 329734 437004 329818
rect 436404 329498 436586 329734
rect 436822 329498 437004 329734
rect 436404 294054 437004 329498
rect 436404 293818 436586 294054
rect 436822 293818 437004 294054
rect 436404 293734 437004 293818
rect 436404 293498 436586 293734
rect 436822 293498 437004 293734
rect 436404 258054 437004 293498
rect 436404 257818 436586 258054
rect 436822 257818 437004 258054
rect 436404 257734 437004 257818
rect 436404 257498 436586 257734
rect 436822 257498 437004 257734
rect 436404 222054 437004 257498
rect 436404 221818 436586 222054
rect 436822 221818 437004 222054
rect 436404 221734 437004 221818
rect 436404 221498 436586 221734
rect 436822 221498 437004 221734
rect 436404 186054 437004 221498
rect 436404 185818 436586 186054
rect 436822 185818 437004 186054
rect 436404 185734 437004 185818
rect 436404 185498 436586 185734
rect 436822 185498 437004 185734
rect 436404 150054 437004 185498
rect 436404 149818 436586 150054
rect 436822 149818 437004 150054
rect 436404 149734 437004 149818
rect 436404 149498 436586 149734
rect 436822 149498 437004 149734
rect 436404 114054 437004 149498
rect 436404 113818 436586 114054
rect 436822 113818 437004 114054
rect 436404 113734 437004 113818
rect 436404 113498 436586 113734
rect 436822 113498 437004 113734
rect 436404 78054 437004 113498
rect 436404 77818 436586 78054
rect 436822 77818 437004 78054
rect 436404 77734 437004 77818
rect 436404 77498 436586 77734
rect 436822 77498 437004 77734
rect 436404 42054 437004 77498
rect 436404 41818 436586 42054
rect 436822 41818 437004 42054
rect 436404 41734 437004 41818
rect 436404 41498 436586 41734
rect 436822 41498 437004 41734
rect 436404 6054 437004 41498
rect 436404 5818 436586 6054
rect 436822 5818 437004 6054
rect 436404 5734 437004 5818
rect 436404 5498 436586 5734
rect 436822 5498 437004 5734
rect 436404 -2186 437004 5498
rect 436404 -2422 436586 -2186
rect 436822 -2422 437004 -2186
rect 436404 -2506 437004 -2422
rect 436404 -2742 436586 -2506
rect 436822 -2742 437004 -2506
rect 436404 -3684 437004 -2742
rect 440004 693654 440604 707962
rect 440004 693418 440186 693654
rect 440422 693418 440604 693654
rect 440004 693334 440604 693418
rect 440004 693098 440186 693334
rect 440422 693098 440604 693334
rect 440004 657654 440604 693098
rect 440004 657418 440186 657654
rect 440422 657418 440604 657654
rect 440004 657334 440604 657418
rect 440004 657098 440186 657334
rect 440422 657098 440604 657334
rect 440004 621654 440604 657098
rect 440004 621418 440186 621654
rect 440422 621418 440604 621654
rect 440004 621334 440604 621418
rect 440004 621098 440186 621334
rect 440422 621098 440604 621334
rect 440004 585654 440604 621098
rect 440004 585418 440186 585654
rect 440422 585418 440604 585654
rect 440004 585334 440604 585418
rect 440004 585098 440186 585334
rect 440422 585098 440604 585334
rect 440004 549654 440604 585098
rect 440004 549418 440186 549654
rect 440422 549418 440604 549654
rect 440004 549334 440604 549418
rect 440004 549098 440186 549334
rect 440422 549098 440604 549334
rect 440004 513654 440604 549098
rect 440004 513418 440186 513654
rect 440422 513418 440604 513654
rect 440004 513334 440604 513418
rect 440004 513098 440186 513334
rect 440422 513098 440604 513334
rect 440004 477654 440604 513098
rect 440004 477418 440186 477654
rect 440422 477418 440604 477654
rect 440004 477334 440604 477418
rect 440004 477098 440186 477334
rect 440422 477098 440604 477334
rect 440004 441654 440604 477098
rect 440004 441418 440186 441654
rect 440422 441418 440604 441654
rect 440004 441334 440604 441418
rect 440004 441098 440186 441334
rect 440422 441098 440604 441334
rect 440004 405654 440604 441098
rect 440004 405418 440186 405654
rect 440422 405418 440604 405654
rect 440004 405334 440604 405418
rect 440004 405098 440186 405334
rect 440422 405098 440604 405334
rect 440004 369654 440604 405098
rect 440004 369418 440186 369654
rect 440422 369418 440604 369654
rect 440004 369334 440604 369418
rect 440004 369098 440186 369334
rect 440422 369098 440604 369334
rect 440004 333654 440604 369098
rect 440004 333418 440186 333654
rect 440422 333418 440604 333654
rect 440004 333334 440604 333418
rect 440004 333098 440186 333334
rect 440422 333098 440604 333334
rect 440004 297654 440604 333098
rect 440004 297418 440186 297654
rect 440422 297418 440604 297654
rect 440004 297334 440604 297418
rect 440004 297098 440186 297334
rect 440422 297098 440604 297334
rect 440004 261654 440604 297098
rect 440004 261418 440186 261654
rect 440422 261418 440604 261654
rect 440004 261334 440604 261418
rect 440004 261098 440186 261334
rect 440422 261098 440604 261334
rect 440004 225654 440604 261098
rect 440004 225418 440186 225654
rect 440422 225418 440604 225654
rect 440004 225334 440604 225418
rect 440004 225098 440186 225334
rect 440422 225098 440604 225334
rect 440004 189654 440604 225098
rect 440004 189418 440186 189654
rect 440422 189418 440604 189654
rect 440004 189334 440604 189418
rect 440004 189098 440186 189334
rect 440422 189098 440604 189334
rect 440004 153654 440604 189098
rect 440004 153418 440186 153654
rect 440422 153418 440604 153654
rect 440004 153334 440604 153418
rect 440004 153098 440186 153334
rect 440422 153098 440604 153334
rect 440004 117654 440604 153098
rect 440004 117418 440186 117654
rect 440422 117418 440604 117654
rect 440004 117334 440604 117418
rect 440004 117098 440186 117334
rect 440422 117098 440604 117334
rect 440004 81654 440604 117098
rect 440004 81418 440186 81654
rect 440422 81418 440604 81654
rect 440004 81334 440604 81418
rect 440004 81098 440186 81334
rect 440422 81098 440604 81334
rect 440004 45654 440604 81098
rect 440004 45418 440186 45654
rect 440422 45418 440604 45654
rect 440004 45334 440604 45418
rect 440004 45098 440186 45334
rect 440422 45098 440604 45334
rect 440004 9654 440604 45098
rect 440004 9418 440186 9654
rect 440422 9418 440604 9654
rect 440004 9334 440604 9418
rect 440004 9098 440186 9334
rect 440422 9098 440604 9334
rect 440004 -4026 440604 9098
rect 440004 -4262 440186 -4026
rect 440422 -4262 440604 -4026
rect 440004 -4346 440604 -4262
rect 440004 -4582 440186 -4346
rect 440422 -4582 440604 -4346
rect 440004 -5524 440604 -4582
rect 443604 697254 444204 709802
rect 461604 711278 462204 711300
rect 461604 711042 461786 711278
rect 462022 711042 462204 711278
rect 461604 710958 462204 711042
rect 461604 710722 461786 710958
rect 462022 710722 462204 710958
rect 458004 709438 458604 709460
rect 458004 709202 458186 709438
rect 458422 709202 458604 709438
rect 458004 709118 458604 709202
rect 458004 708882 458186 709118
rect 458422 708882 458604 709118
rect 454404 707598 455004 707620
rect 454404 707362 454586 707598
rect 454822 707362 455004 707598
rect 454404 707278 455004 707362
rect 454404 707042 454586 707278
rect 454822 707042 455004 707278
rect 443604 697018 443786 697254
rect 444022 697018 444204 697254
rect 443604 696934 444204 697018
rect 443604 696698 443786 696934
rect 444022 696698 444204 696934
rect 443604 661254 444204 696698
rect 443604 661018 443786 661254
rect 444022 661018 444204 661254
rect 443604 660934 444204 661018
rect 443604 660698 443786 660934
rect 444022 660698 444204 660934
rect 443604 625254 444204 660698
rect 443604 625018 443786 625254
rect 444022 625018 444204 625254
rect 443604 624934 444204 625018
rect 443604 624698 443786 624934
rect 444022 624698 444204 624934
rect 443604 589254 444204 624698
rect 443604 589018 443786 589254
rect 444022 589018 444204 589254
rect 443604 588934 444204 589018
rect 443604 588698 443786 588934
rect 444022 588698 444204 588934
rect 443604 553254 444204 588698
rect 443604 553018 443786 553254
rect 444022 553018 444204 553254
rect 443604 552934 444204 553018
rect 443604 552698 443786 552934
rect 444022 552698 444204 552934
rect 443604 517254 444204 552698
rect 443604 517018 443786 517254
rect 444022 517018 444204 517254
rect 443604 516934 444204 517018
rect 443604 516698 443786 516934
rect 444022 516698 444204 516934
rect 443604 481254 444204 516698
rect 443604 481018 443786 481254
rect 444022 481018 444204 481254
rect 443604 480934 444204 481018
rect 443604 480698 443786 480934
rect 444022 480698 444204 480934
rect 443604 445254 444204 480698
rect 443604 445018 443786 445254
rect 444022 445018 444204 445254
rect 443604 444934 444204 445018
rect 443604 444698 443786 444934
rect 444022 444698 444204 444934
rect 443604 409254 444204 444698
rect 443604 409018 443786 409254
rect 444022 409018 444204 409254
rect 443604 408934 444204 409018
rect 443604 408698 443786 408934
rect 444022 408698 444204 408934
rect 443604 373254 444204 408698
rect 443604 373018 443786 373254
rect 444022 373018 444204 373254
rect 443604 372934 444204 373018
rect 443604 372698 443786 372934
rect 444022 372698 444204 372934
rect 443604 337254 444204 372698
rect 443604 337018 443786 337254
rect 444022 337018 444204 337254
rect 443604 336934 444204 337018
rect 443604 336698 443786 336934
rect 444022 336698 444204 336934
rect 443604 301254 444204 336698
rect 443604 301018 443786 301254
rect 444022 301018 444204 301254
rect 443604 300934 444204 301018
rect 443604 300698 443786 300934
rect 444022 300698 444204 300934
rect 443604 265254 444204 300698
rect 443604 265018 443786 265254
rect 444022 265018 444204 265254
rect 443604 264934 444204 265018
rect 443604 264698 443786 264934
rect 444022 264698 444204 264934
rect 443604 229254 444204 264698
rect 443604 229018 443786 229254
rect 444022 229018 444204 229254
rect 443604 228934 444204 229018
rect 443604 228698 443786 228934
rect 444022 228698 444204 228934
rect 443604 193254 444204 228698
rect 443604 193018 443786 193254
rect 444022 193018 444204 193254
rect 443604 192934 444204 193018
rect 443604 192698 443786 192934
rect 444022 192698 444204 192934
rect 443604 157254 444204 192698
rect 443604 157018 443786 157254
rect 444022 157018 444204 157254
rect 443604 156934 444204 157018
rect 443604 156698 443786 156934
rect 444022 156698 444204 156934
rect 443604 121254 444204 156698
rect 443604 121018 443786 121254
rect 444022 121018 444204 121254
rect 443604 120934 444204 121018
rect 443604 120698 443786 120934
rect 444022 120698 444204 120934
rect 443604 85254 444204 120698
rect 443604 85018 443786 85254
rect 444022 85018 444204 85254
rect 443604 84934 444204 85018
rect 443604 84698 443786 84934
rect 444022 84698 444204 84934
rect 443604 49254 444204 84698
rect 443604 49018 443786 49254
rect 444022 49018 444204 49254
rect 443604 48934 444204 49018
rect 443604 48698 443786 48934
rect 444022 48698 444204 48934
rect 443604 13254 444204 48698
rect 443604 13018 443786 13254
rect 444022 13018 444204 13254
rect 443604 12934 444204 13018
rect 443604 12698 443786 12934
rect 444022 12698 444204 12934
rect 425604 -7022 425786 -6786
rect 426022 -7022 426204 -6786
rect 425604 -7106 426204 -7022
rect 425604 -7342 425786 -7106
rect 426022 -7342 426204 -7106
rect 425604 -7364 426204 -7342
rect 443604 -5866 444204 12698
rect 450804 705758 451404 705780
rect 450804 705522 450986 705758
rect 451222 705522 451404 705758
rect 450804 705438 451404 705522
rect 450804 705202 450986 705438
rect 451222 705202 451404 705438
rect 450804 668454 451404 705202
rect 450804 668218 450986 668454
rect 451222 668218 451404 668454
rect 450804 668134 451404 668218
rect 450804 667898 450986 668134
rect 451222 667898 451404 668134
rect 450804 632454 451404 667898
rect 450804 632218 450986 632454
rect 451222 632218 451404 632454
rect 450804 632134 451404 632218
rect 450804 631898 450986 632134
rect 451222 631898 451404 632134
rect 450804 596454 451404 631898
rect 450804 596218 450986 596454
rect 451222 596218 451404 596454
rect 450804 596134 451404 596218
rect 450804 595898 450986 596134
rect 451222 595898 451404 596134
rect 450804 560454 451404 595898
rect 450804 560218 450986 560454
rect 451222 560218 451404 560454
rect 450804 560134 451404 560218
rect 450804 559898 450986 560134
rect 451222 559898 451404 560134
rect 450804 524454 451404 559898
rect 450804 524218 450986 524454
rect 451222 524218 451404 524454
rect 450804 524134 451404 524218
rect 450804 523898 450986 524134
rect 451222 523898 451404 524134
rect 450804 488454 451404 523898
rect 450804 488218 450986 488454
rect 451222 488218 451404 488454
rect 450804 488134 451404 488218
rect 450804 487898 450986 488134
rect 451222 487898 451404 488134
rect 450804 452454 451404 487898
rect 450804 452218 450986 452454
rect 451222 452218 451404 452454
rect 450804 452134 451404 452218
rect 450804 451898 450986 452134
rect 451222 451898 451404 452134
rect 450804 416454 451404 451898
rect 450804 416218 450986 416454
rect 451222 416218 451404 416454
rect 450804 416134 451404 416218
rect 450804 415898 450986 416134
rect 451222 415898 451404 416134
rect 450804 380454 451404 415898
rect 450804 380218 450986 380454
rect 451222 380218 451404 380454
rect 450804 380134 451404 380218
rect 450804 379898 450986 380134
rect 451222 379898 451404 380134
rect 450804 344454 451404 379898
rect 450804 344218 450986 344454
rect 451222 344218 451404 344454
rect 450804 344134 451404 344218
rect 450804 343898 450986 344134
rect 451222 343898 451404 344134
rect 450804 308454 451404 343898
rect 450804 308218 450986 308454
rect 451222 308218 451404 308454
rect 450804 308134 451404 308218
rect 450804 307898 450986 308134
rect 451222 307898 451404 308134
rect 450804 272454 451404 307898
rect 450804 272218 450986 272454
rect 451222 272218 451404 272454
rect 450804 272134 451404 272218
rect 450804 271898 450986 272134
rect 451222 271898 451404 272134
rect 450804 236454 451404 271898
rect 450804 236218 450986 236454
rect 451222 236218 451404 236454
rect 450804 236134 451404 236218
rect 450804 235898 450986 236134
rect 451222 235898 451404 236134
rect 450804 200454 451404 235898
rect 450804 200218 450986 200454
rect 451222 200218 451404 200454
rect 450804 200134 451404 200218
rect 450804 199898 450986 200134
rect 451222 199898 451404 200134
rect 450804 164454 451404 199898
rect 450804 164218 450986 164454
rect 451222 164218 451404 164454
rect 450804 164134 451404 164218
rect 450804 163898 450986 164134
rect 451222 163898 451404 164134
rect 450804 128454 451404 163898
rect 450804 128218 450986 128454
rect 451222 128218 451404 128454
rect 450804 128134 451404 128218
rect 450804 127898 450986 128134
rect 451222 127898 451404 128134
rect 450804 92454 451404 127898
rect 450804 92218 450986 92454
rect 451222 92218 451404 92454
rect 450804 92134 451404 92218
rect 450804 91898 450986 92134
rect 451222 91898 451404 92134
rect 450804 56454 451404 91898
rect 450804 56218 450986 56454
rect 451222 56218 451404 56454
rect 450804 56134 451404 56218
rect 450804 55898 450986 56134
rect 451222 55898 451404 56134
rect 450804 20454 451404 55898
rect 450804 20218 450986 20454
rect 451222 20218 451404 20454
rect 450804 20134 451404 20218
rect 450804 19898 450986 20134
rect 451222 19898 451404 20134
rect 450804 -1266 451404 19898
rect 450804 -1502 450986 -1266
rect 451222 -1502 451404 -1266
rect 450804 -1586 451404 -1502
rect 450804 -1822 450986 -1586
rect 451222 -1822 451404 -1586
rect 450804 -1844 451404 -1822
rect 454404 672054 455004 707042
rect 454404 671818 454586 672054
rect 454822 671818 455004 672054
rect 454404 671734 455004 671818
rect 454404 671498 454586 671734
rect 454822 671498 455004 671734
rect 454404 636054 455004 671498
rect 454404 635818 454586 636054
rect 454822 635818 455004 636054
rect 454404 635734 455004 635818
rect 454404 635498 454586 635734
rect 454822 635498 455004 635734
rect 454404 600054 455004 635498
rect 454404 599818 454586 600054
rect 454822 599818 455004 600054
rect 454404 599734 455004 599818
rect 454404 599498 454586 599734
rect 454822 599498 455004 599734
rect 454404 564054 455004 599498
rect 454404 563818 454586 564054
rect 454822 563818 455004 564054
rect 454404 563734 455004 563818
rect 454404 563498 454586 563734
rect 454822 563498 455004 563734
rect 454404 528054 455004 563498
rect 454404 527818 454586 528054
rect 454822 527818 455004 528054
rect 454404 527734 455004 527818
rect 454404 527498 454586 527734
rect 454822 527498 455004 527734
rect 454404 492054 455004 527498
rect 454404 491818 454586 492054
rect 454822 491818 455004 492054
rect 454404 491734 455004 491818
rect 454404 491498 454586 491734
rect 454822 491498 455004 491734
rect 454404 456054 455004 491498
rect 454404 455818 454586 456054
rect 454822 455818 455004 456054
rect 454404 455734 455004 455818
rect 454404 455498 454586 455734
rect 454822 455498 455004 455734
rect 454404 420054 455004 455498
rect 454404 419818 454586 420054
rect 454822 419818 455004 420054
rect 454404 419734 455004 419818
rect 454404 419498 454586 419734
rect 454822 419498 455004 419734
rect 454404 384054 455004 419498
rect 454404 383818 454586 384054
rect 454822 383818 455004 384054
rect 454404 383734 455004 383818
rect 454404 383498 454586 383734
rect 454822 383498 455004 383734
rect 454404 348054 455004 383498
rect 454404 347818 454586 348054
rect 454822 347818 455004 348054
rect 454404 347734 455004 347818
rect 454404 347498 454586 347734
rect 454822 347498 455004 347734
rect 454404 312054 455004 347498
rect 454404 311818 454586 312054
rect 454822 311818 455004 312054
rect 454404 311734 455004 311818
rect 454404 311498 454586 311734
rect 454822 311498 455004 311734
rect 454404 276054 455004 311498
rect 454404 275818 454586 276054
rect 454822 275818 455004 276054
rect 454404 275734 455004 275818
rect 454404 275498 454586 275734
rect 454822 275498 455004 275734
rect 454404 240054 455004 275498
rect 454404 239818 454586 240054
rect 454822 239818 455004 240054
rect 454404 239734 455004 239818
rect 454404 239498 454586 239734
rect 454822 239498 455004 239734
rect 454404 204054 455004 239498
rect 454404 203818 454586 204054
rect 454822 203818 455004 204054
rect 454404 203734 455004 203818
rect 454404 203498 454586 203734
rect 454822 203498 455004 203734
rect 454404 168054 455004 203498
rect 454404 167818 454586 168054
rect 454822 167818 455004 168054
rect 454404 167734 455004 167818
rect 454404 167498 454586 167734
rect 454822 167498 455004 167734
rect 454404 132054 455004 167498
rect 454404 131818 454586 132054
rect 454822 131818 455004 132054
rect 454404 131734 455004 131818
rect 454404 131498 454586 131734
rect 454822 131498 455004 131734
rect 454404 96054 455004 131498
rect 454404 95818 454586 96054
rect 454822 95818 455004 96054
rect 454404 95734 455004 95818
rect 454404 95498 454586 95734
rect 454822 95498 455004 95734
rect 454404 60054 455004 95498
rect 454404 59818 454586 60054
rect 454822 59818 455004 60054
rect 454404 59734 455004 59818
rect 454404 59498 454586 59734
rect 454822 59498 455004 59734
rect 454404 24054 455004 59498
rect 454404 23818 454586 24054
rect 454822 23818 455004 24054
rect 454404 23734 455004 23818
rect 454404 23498 454586 23734
rect 454822 23498 455004 23734
rect 454404 -3106 455004 23498
rect 454404 -3342 454586 -3106
rect 454822 -3342 455004 -3106
rect 454404 -3426 455004 -3342
rect 454404 -3662 454586 -3426
rect 454822 -3662 455004 -3426
rect 454404 -3684 455004 -3662
rect 458004 675654 458604 708882
rect 458004 675418 458186 675654
rect 458422 675418 458604 675654
rect 458004 675334 458604 675418
rect 458004 675098 458186 675334
rect 458422 675098 458604 675334
rect 458004 639654 458604 675098
rect 458004 639418 458186 639654
rect 458422 639418 458604 639654
rect 458004 639334 458604 639418
rect 458004 639098 458186 639334
rect 458422 639098 458604 639334
rect 458004 603654 458604 639098
rect 458004 603418 458186 603654
rect 458422 603418 458604 603654
rect 458004 603334 458604 603418
rect 458004 603098 458186 603334
rect 458422 603098 458604 603334
rect 458004 567654 458604 603098
rect 458004 567418 458186 567654
rect 458422 567418 458604 567654
rect 458004 567334 458604 567418
rect 458004 567098 458186 567334
rect 458422 567098 458604 567334
rect 458004 531654 458604 567098
rect 458004 531418 458186 531654
rect 458422 531418 458604 531654
rect 458004 531334 458604 531418
rect 458004 531098 458186 531334
rect 458422 531098 458604 531334
rect 458004 495654 458604 531098
rect 458004 495418 458186 495654
rect 458422 495418 458604 495654
rect 458004 495334 458604 495418
rect 458004 495098 458186 495334
rect 458422 495098 458604 495334
rect 458004 459654 458604 495098
rect 458004 459418 458186 459654
rect 458422 459418 458604 459654
rect 458004 459334 458604 459418
rect 458004 459098 458186 459334
rect 458422 459098 458604 459334
rect 458004 423654 458604 459098
rect 458004 423418 458186 423654
rect 458422 423418 458604 423654
rect 458004 423334 458604 423418
rect 458004 423098 458186 423334
rect 458422 423098 458604 423334
rect 458004 387654 458604 423098
rect 458004 387418 458186 387654
rect 458422 387418 458604 387654
rect 458004 387334 458604 387418
rect 458004 387098 458186 387334
rect 458422 387098 458604 387334
rect 458004 351654 458604 387098
rect 458004 351418 458186 351654
rect 458422 351418 458604 351654
rect 458004 351334 458604 351418
rect 458004 351098 458186 351334
rect 458422 351098 458604 351334
rect 458004 315654 458604 351098
rect 458004 315418 458186 315654
rect 458422 315418 458604 315654
rect 458004 315334 458604 315418
rect 458004 315098 458186 315334
rect 458422 315098 458604 315334
rect 458004 279654 458604 315098
rect 458004 279418 458186 279654
rect 458422 279418 458604 279654
rect 458004 279334 458604 279418
rect 458004 279098 458186 279334
rect 458422 279098 458604 279334
rect 458004 243654 458604 279098
rect 458004 243418 458186 243654
rect 458422 243418 458604 243654
rect 458004 243334 458604 243418
rect 458004 243098 458186 243334
rect 458422 243098 458604 243334
rect 458004 207654 458604 243098
rect 458004 207418 458186 207654
rect 458422 207418 458604 207654
rect 458004 207334 458604 207418
rect 458004 207098 458186 207334
rect 458422 207098 458604 207334
rect 458004 171654 458604 207098
rect 458004 171418 458186 171654
rect 458422 171418 458604 171654
rect 458004 171334 458604 171418
rect 458004 171098 458186 171334
rect 458422 171098 458604 171334
rect 458004 135654 458604 171098
rect 458004 135418 458186 135654
rect 458422 135418 458604 135654
rect 458004 135334 458604 135418
rect 458004 135098 458186 135334
rect 458422 135098 458604 135334
rect 458004 99654 458604 135098
rect 458004 99418 458186 99654
rect 458422 99418 458604 99654
rect 458004 99334 458604 99418
rect 458004 99098 458186 99334
rect 458422 99098 458604 99334
rect 458004 63654 458604 99098
rect 458004 63418 458186 63654
rect 458422 63418 458604 63654
rect 458004 63334 458604 63418
rect 458004 63098 458186 63334
rect 458422 63098 458604 63334
rect 458004 27654 458604 63098
rect 458004 27418 458186 27654
rect 458422 27418 458604 27654
rect 458004 27334 458604 27418
rect 458004 27098 458186 27334
rect 458422 27098 458604 27334
rect 458004 -4946 458604 27098
rect 458004 -5182 458186 -4946
rect 458422 -5182 458604 -4946
rect 458004 -5266 458604 -5182
rect 458004 -5502 458186 -5266
rect 458422 -5502 458604 -5266
rect 458004 -5524 458604 -5502
rect 461604 679254 462204 710722
rect 479604 710358 480204 711300
rect 479604 710122 479786 710358
rect 480022 710122 480204 710358
rect 479604 710038 480204 710122
rect 479604 709802 479786 710038
rect 480022 709802 480204 710038
rect 476004 708518 476604 709460
rect 476004 708282 476186 708518
rect 476422 708282 476604 708518
rect 476004 708198 476604 708282
rect 476004 707962 476186 708198
rect 476422 707962 476604 708198
rect 472404 706678 473004 707620
rect 472404 706442 472586 706678
rect 472822 706442 473004 706678
rect 472404 706358 473004 706442
rect 472404 706122 472586 706358
rect 472822 706122 473004 706358
rect 461604 679018 461786 679254
rect 462022 679018 462204 679254
rect 461604 678934 462204 679018
rect 461604 678698 461786 678934
rect 462022 678698 462204 678934
rect 461604 643254 462204 678698
rect 461604 643018 461786 643254
rect 462022 643018 462204 643254
rect 461604 642934 462204 643018
rect 461604 642698 461786 642934
rect 462022 642698 462204 642934
rect 461604 607254 462204 642698
rect 461604 607018 461786 607254
rect 462022 607018 462204 607254
rect 461604 606934 462204 607018
rect 461604 606698 461786 606934
rect 462022 606698 462204 606934
rect 461604 571254 462204 606698
rect 461604 571018 461786 571254
rect 462022 571018 462204 571254
rect 461604 570934 462204 571018
rect 461604 570698 461786 570934
rect 462022 570698 462204 570934
rect 461604 535254 462204 570698
rect 461604 535018 461786 535254
rect 462022 535018 462204 535254
rect 461604 534934 462204 535018
rect 461604 534698 461786 534934
rect 462022 534698 462204 534934
rect 461604 499254 462204 534698
rect 461604 499018 461786 499254
rect 462022 499018 462204 499254
rect 461604 498934 462204 499018
rect 461604 498698 461786 498934
rect 462022 498698 462204 498934
rect 461604 463254 462204 498698
rect 461604 463018 461786 463254
rect 462022 463018 462204 463254
rect 461604 462934 462204 463018
rect 461604 462698 461786 462934
rect 462022 462698 462204 462934
rect 461604 427254 462204 462698
rect 461604 427018 461786 427254
rect 462022 427018 462204 427254
rect 461604 426934 462204 427018
rect 461604 426698 461786 426934
rect 462022 426698 462204 426934
rect 461604 391254 462204 426698
rect 461604 391018 461786 391254
rect 462022 391018 462204 391254
rect 461604 390934 462204 391018
rect 461604 390698 461786 390934
rect 462022 390698 462204 390934
rect 461604 355254 462204 390698
rect 461604 355018 461786 355254
rect 462022 355018 462204 355254
rect 461604 354934 462204 355018
rect 461604 354698 461786 354934
rect 462022 354698 462204 354934
rect 461604 319254 462204 354698
rect 461604 319018 461786 319254
rect 462022 319018 462204 319254
rect 461604 318934 462204 319018
rect 461604 318698 461786 318934
rect 462022 318698 462204 318934
rect 461604 283254 462204 318698
rect 461604 283018 461786 283254
rect 462022 283018 462204 283254
rect 461604 282934 462204 283018
rect 461604 282698 461786 282934
rect 462022 282698 462204 282934
rect 461604 247254 462204 282698
rect 461604 247018 461786 247254
rect 462022 247018 462204 247254
rect 461604 246934 462204 247018
rect 461604 246698 461786 246934
rect 462022 246698 462204 246934
rect 461604 211254 462204 246698
rect 461604 211018 461786 211254
rect 462022 211018 462204 211254
rect 461604 210934 462204 211018
rect 461604 210698 461786 210934
rect 462022 210698 462204 210934
rect 461604 175254 462204 210698
rect 461604 175018 461786 175254
rect 462022 175018 462204 175254
rect 461604 174934 462204 175018
rect 461604 174698 461786 174934
rect 462022 174698 462204 174934
rect 461604 139254 462204 174698
rect 461604 139018 461786 139254
rect 462022 139018 462204 139254
rect 461604 138934 462204 139018
rect 461604 138698 461786 138934
rect 462022 138698 462204 138934
rect 461604 103254 462204 138698
rect 461604 103018 461786 103254
rect 462022 103018 462204 103254
rect 461604 102934 462204 103018
rect 461604 102698 461786 102934
rect 462022 102698 462204 102934
rect 461604 67254 462204 102698
rect 461604 67018 461786 67254
rect 462022 67018 462204 67254
rect 461604 66934 462204 67018
rect 461604 66698 461786 66934
rect 462022 66698 462204 66934
rect 461604 31254 462204 66698
rect 461604 31018 461786 31254
rect 462022 31018 462204 31254
rect 461604 30934 462204 31018
rect 461604 30698 461786 30934
rect 462022 30698 462204 30934
rect 443604 -6102 443786 -5866
rect 444022 -6102 444204 -5866
rect 443604 -6186 444204 -6102
rect 443604 -6422 443786 -6186
rect 444022 -6422 444204 -6186
rect 443604 -7364 444204 -6422
rect 461604 -6786 462204 30698
rect 468804 704838 469404 705780
rect 468804 704602 468986 704838
rect 469222 704602 469404 704838
rect 468804 704518 469404 704602
rect 468804 704282 468986 704518
rect 469222 704282 469404 704518
rect 468804 686454 469404 704282
rect 468804 686218 468986 686454
rect 469222 686218 469404 686454
rect 468804 686134 469404 686218
rect 468804 685898 468986 686134
rect 469222 685898 469404 686134
rect 468804 650454 469404 685898
rect 468804 650218 468986 650454
rect 469222 650218 469404 650454
rect 468804 650134 469404 650218
rect 468804 649898 468986 650134
rect 469222 649898 469404 650134
rect 468804 614454 469404 649898
rect 468804 614218 468986 614454
rect 469222 614218 469404 614454
rect 468804 614134 469404 614218
rect 468804 613898 468986 614134
rect 469222 613898 469404 614134
rect 468804 578454 469404 613898
rect 468804 578218 468986 578454
rect 469222 578218 469404 578454
rect 468804 578134 469404 578218
rect 468804 577898 468986 578134
rect 469222 577898 469404 578134
rect 468804 542454 469404 577898
rect 468804 542218 468986 542454
rect 469222 542218 469404 542454
rect 468804 542134 469404 542218
rect 468804 541898 468986 542134
rect 469222 541898 469404 542134
rect 468804 506454 469404 541898
rect 468804 506218 468986 506454
rect 469222 506218 469404 506454
rect 468804 506134 469404 506218
rect 468804 505898 468986 506134
rect 469222 505898 469404 506134
rect 468804 470454 469404 505898
rect 468804 470218 468986 470454
rect 469222 470218 469404 470454
rect 468804 470134 469404 470218
rect 468804 469898 468986 470134
rect 469222 469898 469404 470134
rect 468804 434454 469404 469898
rect 468804 434218 468986 434454
rect 469222 434218 469404 434454
rect 468804 434134 469404 434218
rect 468804 433898 468986 434134
rect 469222 433898 469404 434134
rect 468804 398454 469404 433898
rect 468804 398218 468986 398454
rect 469222 398218 469404 398454
rect 468804 398134 469404 398218
rect 468804 397898 468986 398134
rect 469222 397898 469404 398134
rect 468804 362454 469404 397898
rect 468804 362218 468986 362454
rect 469222 362218 469404 362454
rect 468804 362134 469404 362218
rect 468804 361898 468986 362134
rect 469222 361898 469404 362134
rect 468804 326454 469404 361898
rect 468804 326218 468986 326454
rect 469222 326218 469404 326454
rect 468804 326134 469404 326218
rect 468804 325898 468986 326134
rect 469222 325898 469404 326134
rect 468804 290454 469404 325898
rect 468804 290218 468986 290454
rect 469222 290218 469404 290454
rect 468804 290134 469404 290218
rect 468804 289898 468986 290134
rect 469222 289898 469404 290134
rect 468804 254454 469404 289898
rect 468804 254218 468986 254454
rect 469222 254218 469404 254454
rect 468804 254134 469404 254218
rect 468804 253898 468986 254134
rect 469222 253898 469404 254134
rect 468804 218454 469404 253898
rect 468804 218218 468986 218454
rect 469222 218218 469404 218454
rect 468804 218134 469404 218218
rect 468804 217898 468986 218134
rect 469222 217898 469404 218134
rect 468804 182454 469404 217898
rect 468804 182218 468986 182454
rect 469222 182218 469404 182454
rect 468804 182134 469404 182218
rect 468804 181898 468986 182134
rect 469222 181898 469404 182134
rect 468804 146454 469404 181898
rect 468804 146218 468986 146454
rect 469222 146218 469404 146454
rect 468804 146134 469404 146218
rect 468804 145898 468986 146134
rect 469222 145898 469404 146134
rect 468804 110454 469404 145898
rect 468804 110218 468986 110454
rect 469222 110218 469404 110454
rect 468804 110134 469404 110218
rect 468804 109898 468986 110134
rect 469222 109898 469404 110134
rect 468804 74454 469404 109898
rect 468804 74218 468986 74454
rect 469222 74218 469404 74454
rect 468804 74134 469404 74218
rect 468804 73898 468986 74134
rect 469222 73898 469404 74134
rect 468804 38454 469404 73898
rect 468804 38218 468986 38454
rect 469222 38218 469404 38454
rect 468804 38134 469404 38218
rect 468804 37898 468986 38134
rect 469222 37898 469404 38134
rect 468804 2454 469404 37898
rect 468804 2218 468986 2454
rect 469222 2218 469404 2454
rect 468804 2134 469404 2218
rect 468804 1898 468986 2134
rect 469222 1898 469404 2134
rect 468804 -346 469404 1898
rect 468804 -582 468986 -346
rect 469222 -582 469404 -346
rect 468804 -666 469404 -582
rect 468804 -902 468986 -666
rect 469222 -902 469404 -666
rect 468804 -1844 469404 -902
rect 472404 690054 473004 706122
rect 472404 689818 472586 690054
rect 472822 689818 473004 690054
rect 472404 689734 473004 689818
rect 472404 689498 472586 689734
rect 472822 689498 473004 689734
rect 472404 654054 473004 689498
rect 472404 653818 472586 654054
rect 472822 653818 473004 654054
rect 472404 653734 473004 653818
rect 472404 653498 472586 653734
rect 472822 653498 473004 653734
rect 472404 618054 473004 653498
rect 472404 617818 472586 618054
rect 472822 617818 473004 618054
rect 472404 617734 473004 617818
rect 472404 617498 472586 617734
rect 472822 617498 473004 617734
rect 472404 582054 473004 617498
rect 472404 581818 472586 582054
rect 472822 581818 473004 582054
rect 472404 581734 473004 581818
rect 472404 581498 472586 581734
rect 472822 581498 473004 581734
rect 472404 546054 473004 581498
rect 472404 545818 472586 546054
rect 472822 545818 473004 546054
rect 472404 545734 473004 545818
rect 472404 545498 472586 545734
rect 472822 545498 473004 545734
rect 472404 510054 473004 545498
rect 472404 509818 472586 510054
rect 472822 509818 473004 510054
rect 472404 509734 473004 509818
rect 472404 509498 472586 509734
rect 472822 509498 473004 509734
rect 472404 474054 473004 509498
rect 472404 473818 472586 474054
rect 472822 473818 473004 474054
rect 472404 473734 473004 473818
rect 472404 473498 472586 473734
rect 472822 473498 473004 473734
rect 472404 438054 473004 473498
rect 472404 437818 472586 438054
rect 472822 437818 473004 438054
rect 472404 437734 473004 437818
rect 472404 437498 472586 437734
rect 472822 437498 473004 437734
rect 472404 402054 473004 437498
rect 472404 401818 472586 402054
rect 472822 401818 473004 402054
rect 472404 401734 473004 401818
rect 472404 401498 472586 401734
rect 472822 401498 473004 401734
rect 472404 366054 473004 401498
rect 472404 365818 472586 366054
rect 472822 365818 473004 366054
rect 472404 365734 473004 365818
rect 472404 365498 472586 365734
rect 472822 365498 473004 365734
rect 472404 330054 473004 365498
rect 472404 329818 472586 330054
rect 472822 329818 473004 330054
rect 472404 329734 473004 329818
rect 472404 329498 472586 329734
rect 472822 329498 473004 329734
rect 472404 294054 473004 329498
rect 472404 293818 472586 294054
rect 472822 293818 473004 294054
rect 472404 293734 473004 293818
rect 472404 293498 472586 293734
rect 472822 293498 473004 293734
rect 472404 258054 473004 293498
rect 472404 257818 472586 258054
rect 472822 257818 473004 258054
rect 472404 257734 473004 257818
rect 472404 257498 472586 257734
rect 472822 257498 473004 257734
rect 472404 222054 473004 257498
rect 472404 221818 472586 222054
rect 472822 221818 473004 222054
rect 472404 221734 473004 221818
rect 472404 221498 472586 221734
rect 472822 221498 473004 221734
rect 472404 186054 473004 221498
rect 472404 185818 472586 186054
rect 472822 185818 473004 186054
rect 472404 185734 473004 185818
rect 472404 185498 472586 185734
rect 472822 185498 473004 185734
rect 472404 150054 473004 185498
rect 472404 149818 472586 150054
rect 472822 149818 473004 150054
rect 472404 149734 473004 149818
rect 472404 149498 472586 149734
rect 472822 149498 473004 149734
rect 472404 114054 473004 149498
rect 472404 113818 472586 114054
rect 472822 113818 473004 114054
rect 472404 113734 473004 113818
rect 472404 113498 472586 113734
rect 472822 113498 473004 113734
rect 472404 78054 473004 113498
rect 472404 77818 472586 78054
rect 472822 77818 473004 78054
rect 472404 77734 473004 77818
rect 472404 77498 472586 77734
rect 472822 77498 473004 77734
rect 472404 42054 473004 77498
rect 472404 41818 472586 42054
rect 472822 41818 473004 42054
rect 472404 41734 473004 41818
rect 472404 41498 472586 41734
rect 472822 41498 473004 41734
rect 472404 6054 473004 41498
rect 472404 5818 472586 6054
rect 472822 5818 473004 6054
rect 472404 5734 473004 5818
rect 472404 5498 472586 5734
rect 472822 5498 473004 5734
rect 472404 -2186 473004 5498
rect 472404 -2422 472586 -2186
rect 472822 -2422 473004 -2186
rect 472404 -2506 473004 -2422
rect 472404 -2742 472586 -2506
rect 472822 -2742 473004 -2506
rect 472404 -3684 473004 -2742
rect 476004 693654 476604 707962
rect 476004 693418 476186 693654
rect 476422 693418 476604 693654
rect 476004 693334 476604 693418
rect 476004 693098 476186 693334
rect 476422 693098 476604 693334
rect 476004 657654 476604 693098
rect 476004 657418 476186 657654
rect 476422 657418 476604 657654
rect 476004 657334 476604 657418
rect 476004 657098 476186 657334
rect 476422 657098 476604 657334
rect 476004 621654 476604 657098
rect 476004 621418 476186 621654
rect 476422 621418 476604 621654
rect 476004 621334 476604 621418
rect 476004 621098 476186 621334
rect 476422 621098 476604 621334
rect 476004 585654 476604 621098
rect 476004 585418 476186 585654
rect 476422 585418 476604 585654
rect 476004 585334 476604 585418
rect 476004 585098 476186 585334
rect 476422 585098 476604 585334
rect 476004 549654 476604 585098
rect 476004 549418 476186 549654
rect 476422 549418 476604 549654
rect 476004 549334 476604 549418
rect 476004 549098 476186 549334
rect 476422 549098 476604 549334
rect 476004 513654 476604 549098
rect 476004 513418 476186 513654
rect 476422 513418 476604 513654
rect 476004 513334 476604 513418
rect 476004 513098 476186 513334
rect 476422 513098 476604 513334
rect 476004 477654 476604 513098
rect 476004 477418 476186 477654
rect 476422 477418 476604 477654
rect 476004 477334 476604 477418
rect 476004 477098 476186 477334
rect 476422 477098 476604 477334
rect 476004 441654 476604 477098
rect 476004 441418 476186 441654
rect 476422 441418 476604 441654
rect 476004 441334 476604 441418
rect 476004 441098 476186 441334
rect 476422 441098 476604 441334
rect 476004 405654 476604 441098
rect 476004 405418 476186 405654
rect 476422 405418 476604 405654
rect 476004 405334 476604 405418
rect 476004 405098 476186 405334
rect 476422 405098 476604 405334
rect 476004 369654 476604 405098
rect 476004 369418 476186 369654
rect 476422 369418 476604 369654
rect 476004 369334 476604 369418
rect 476004 369098 476186 369334
rect 476422 369098 476604 369334
rect 476004 333654 476604 369098
rect 476004 333418 476186 333654
rect 476422 333418 476604 333654
rect 476004 333334 476604 333418
rect 476004 333098 476186 333334
rect 476422 333098 476604 333334
rect 476004 297654 476604 333098
rect 476004 297418 476186 297654
rect 476422 297418 476604 297654
rect 476004 297334 476604 297418
rect 476004 297098 476186 297334
rect 476422 297098 476604 297334
rect 476004 261654 476604 297098
rect 476004 261418 476186 261654
rect 476422 261418 476604 261654
rect 476004 261334 476604 261418
rect 476004 261098 476186 261334
rect 476422 261098 476604 261334
rect 476004 225654 476604 261098
rect 476004 225418 476186 225654
rect 476422 225418 476604 225654
rect 476004 225334 476604 225418
rect 476004 225098 476186 225334
rect 476422 225098 476604 225334
rect 476004 189654 476604 225098
rect 476004 189418 476186 189654
rect 476422 189418 476604 189654
rect 476004 189334 476604 189418
rect 476004 189098 476186 189334
rect 476422 189098 476604 189334
rect 476004 153654 476604 189098
rect 476004 153418 476186 153654
rect 476422 153418 476604 153654
rect 476004 153334 476604 153418
rect 476004 153098 476186 153334
rect 476422 153098 476604 153334
rect 476004 117654 476604 153098
rect 476004 117418 476186 117654
rect 476422 117418 476604 117654
rect 476004 117334 476604 117418
rect 476004 117098 476186 117334
rect 476422 117098 476604 117334
rect 476004 81654 476604 117098
rect 476004 81418 476186 81654
rect 476422 81418 476604 81654
rect 476004 81334 476604 81418
rect 476004 81098 476186 81334
rect 476422 81098 476604 81334
rect 476004 45654 476604 81098
rect 476004 45418 476186 45654
rect 476422 45418 476604 45654
rect 476004 45334 476604 45418
rect 476004 45098 476186 45334
rect 476422 45098 476604 45334
rect 476004 9654 476604 45098
rect 476004 9418 476186 9654
rect 476422 9418 476604 9654
rect 476004 9334 476604 9418
rect 476004 9098 476186 9334
rect 476422 9098 476604 9334
rect 476004 -4026 476604 9098
rect 476004 -4262 476186 -4026
rect 476422 -4262 476604 -4026
rect 476004 -4346 476604 -4262
rect 476004 -4582 476186 -4346
rect 476422 -4582 476604 -4346
rect 476004 -5524 476604 -4582
rect 479604 697254 480204 709802
rect 497604 711278 498204 711300
rect 497604 711042 497786 711278
rect 498022 711042 498204 711278
rect 497604 710958 498204 711042
rect 497604 710722 497786 710958
rect 498022 710722 498204 710958
rect 494004 709438 494604 709460
rect 494004 709202 494186 709438
rect 494422 709202 494604 709438
rect 494004 709118 494604 709202
rect 494004 708882 494186 709118
rect 494422 708882 494604 709118
rect 490404 707598 491004 707620
rect 490404 707362 490586 707598
rect 490822 707362 491004 707598
rect 490404 707278 491004 707362
rect 490404 707042 490586 707278
rect 490822 707042 491004 707278
rect 479604 697018 479786 697254
rect 480022 697018 480204 697254
rect 479604 696934 480204 697018
rect 479604 696698 479786 696934
rect 480022 696698 480204 696934
rect 479604 661254 480204 696698
rect 479604 661018 479786 661254
rect 480022 661018 480204 661254
rect 479604 660934 480204 661018
rect 479604 660698 479786 660934
rect 480022 660698 480204 660934
rect 479604 625254 480204 660698
rect 479604 625018 479786 625254
rect 480022 625018 480204 625254
rect 479604 624934 480204 625018
rect 479604 624698 479786 624934
rect 480022 624698 480204 624934
rect 479604 589254 480204 624698
rect 479604 589018 479786 589254
rect 480022 589018 480204 589254
rect 479604 588934 480204 589018
rect 479604 588698 479786 588934
rect 480022 588698 480204 588934
rect 479604 553254 480204 588698
rect 479604 553018 479786 553254
rect 480022 553018 480204 553254
rect 479604 552934 480204 553018
rect 479604 552698 479786 552934
rect 480022 552698 480204 552934
rect 479604 517254 480204 552698
rect 479604 517018 479786 517254
rect 480022 517018 480204 517254
rect 479604 516934 480204 517018
rect 479604 516698 479786 516934
rect 480022 516698 480204 516934
rect 479604 481254 480204 516698
rect 479604 481018 479786 481254
rect 480022 481018 480204 481254
rect 479604 480934 480204 481018
rect 479604 480698 479786 480934
rect 480022 480698 480204 480934
rect 479604 445254 480204 480698
rect 479604 445018 479786 445254
rect 480022 445018 480204 445254
rect 479604 444934 480204 445018
rect 479604 444698 479786 444934
rect 480022 444698 480204 444934
rect 479604 409254 480204 444698
rect 479604 409018 479786 409254
rect 480022 409018 480204 409254
rect 479604 408934 480204 409018
rect 479604 408698 479786 408934
rect 480022 408698 480204 408934
rect 479604 373254 480204 408698
rect 479604 373018 479786 373254
rect 480022 373018 480204 373254
rect 479604 372934 480204 373018
rect 479604 372698 479786 372934
rect 480022 372698 480204 372934
rect 479604 337254 480204 372698
rect 479604 337018 479786 337254
rect 480022 337018 480204 337254
rect 479604 336934 480204 337018
rect 479604 336698 479786 336934
rect 480022 336698 480204 336934
rect 479604 301254 480204 336698
rect 479604 301018 479786 301254
rect 480022 301018 480204 301254
rect 479604 300934 480204 301018
rect 479604 300698 479786 300934
rect 480022 300698 480204 300934
rect 479604 265254 480204 300698
rect 479604 265018 479786 265254
rect 480022 265018 480204 265254
rect 479604 264934 480204 265018
rect 479604 264698 479786 264934
rect 480022 264698 480204 264934
rect 479604 229254 480204 264698
rect 479604 229018 479786 229254
rect 480022 229018 480204 229254
rect 479604 228934 480204 229018
rect 479604 228698 479786 228934
rect 480022 228698 480204 228934
rect 479604 193254 480204 228698
rect 479604 193018 479786 193254
rect 480022 193018 480204 193254
rect 479604 192934 480204 193018
rect 479604 192698 479786 192934
rect 480022 192698 480204 192934
rect 479604 157254 480204 192698
rect 479604 157018 479786 157254
rect 480022 157018 480204 157254
rect 479604 156934 480204 157018
rect 479604 156698 479786 156934
rect 480022 156698 480204 156934
rect 479604 121254 480204 156698
rect 479604 121018 479786 121254
rect 480022 121018 480204 121254
rect 479604 120934 480204 121018
rect 479604 120698 479786 120934
rect 480022 120698 480204 120934
rect 479604 85254 480204 120698
rect 479604 85018 479786 85254
rect 480022 85018 480204 85254
rect 479604 84934 480204 85018
rect 479604 84698 479786 84934
rect 480022 84698 480204 84934
rect 479604 49254 480204 84698
rect 479604 49018 479786 49254
rect 480022 49018 480204 49254
rect 479604 48934 480204 49018
rect 479604 48698 479786 48934
rect 480022 48698 480204 48934
rect 479604 13254 480204 48698
rect 479604 13018 479786 13254
rect 480022 13018 480204 13254
rect 479604 12934 480204 13018
rect 479604 12698 479786 12934
rect 480022 12698 480204 12934
rect 461604 -7022 461786 -6786
rect 462022 -7022 462204 -6786
rect 461604 -7106 462204 -7022
rect 461604 -7342 461786 -7106
rect 462022 -7342 462204 -7106
rect 461604 -7364 462204 -7342
rect 479604 -5866 480204 12698
rect 486804 705758 487404 705780
rect 486804 705522 486986 705758
rect 487222 705522 487404 705758
rect 486804 705438 487404 705522
rect 486804 705202 486986 705438
rect 487222 705202 487404 705438
rect 486804 668454 487404 705202
rect 486804 668218 486986 668454
rect 487222 668218 487404 668454
rect 486804 668134 487404 668218
rect 486804 667898 486986 668134
rect 487222 667898 487404 668134
rect 486804 632454 487404 667898
rect 486804 632218 486986 632454
rect 487222 632218 487404 632454
rect 486804 632134 487404 632218
rect 486804 631898 486986 632134
rect 487222 631898 487404 632134
rect 486804 596454 487404 631898
rect 486804 596218 486986 596454
rect 487222 596218 487404 596454
rect 486804 596134 487404 596218
rect 486804 595898 486986 596134
rect 487222 595898 487404 596134
rect 486804 560454 487404 595898
rect 486804 560218 486986 560454
rect 487222 560218 487404 560454
rect 486804 560134 487404 560218
rect 486804 559898 486986 560134
rect 487222 559898 487404 560134
rect 486804 524454 487404 559898
rect 486804 524218 486986 524454
rect 487222 524218 487404 524454
rect 486804 524134 487404 524218
rect 486804 523898 486986 524134
rect 487222 523898 487404 524134
rect 486804 488454 487404 523898
rect 486804 488218 486986 488454
rect 487222 488218 487404 488454
rect 486804 488134 487404 488218
rect 486804 487898 486986 488134
rect 487222 487898 487404 488134
rect 486804 452454 487404 487898
rect 486804 452218 486986 452454
rect 487222 452218 487404 452454
rect 486804 452134 487404 452218
rect 486804 451898 486986 452134
rect 487222 451898 487404 452134
rect 486804 416454 487404 451898
rect 486804 416218 486986 416454
rect 487222 416218 487404 416454
rect 486804 416134 487404 416218
rect 486804 415898 486986 416134
rect 487222 415898 487404 416134
rect 486804 380454 487404 415898
rect 486804 380218 486986 380454
rect 487222 380218 487404 380454
rect 486804 380134 487404 380218
rect 486804 379898 486986 380134
rect 487222 379898 487404 380134
rect 486804 344454 487404 379898
rect 486804 344218 486986 344454
rect 487222 344218 487404 344454
rect 486804 344134 487404 344218
rect 486804 343898 486986 344134
rect 487222 343898 487404 344134
rect 486804 308454 487404 343898
rect 486804 308218 486986 308454
rect 487222 308218 487404 308454
rect 486804 308134 487404 308218
rect 486804 307898 486986 308134
rect 487222 307898 487404 308134
rect 486804 272454 487404 307898
rect 486804 272218 486986 272454
rect 487222 272218 487404 272454
rect 486804 272134 487404 272218
rect 486804 271898 486986 272134
rect 487222 271898 487404 272134
rect 486804 236454 487404 271898
rect 486804 236218 486986 236454
rect 487222 236218 487404 236454
rect 486804 236134 487404 236218
rect 486804 235898 486986 236134
rect 487222 235898 487404 236134
rect 486804 200454 487404 235898
rect 486804 200218 486986 200454
rect 487222 200218 487404 200454
rect 486804 200134 487404 200218
rect 486804 199898 486986 200134
rect 487222 199898 487404 200134
rect 486804 164454 487404 199898
rect 486804 164218 486986 164454
rect 487222 164218 487404 164454
rect 486804 164134 487404 164218
rect 486804 163898 486986 164134
rect 487222 163898 487404 164134
rect 486804 128454 487404 163898
rect 486804 128218 486986 128454
rect 487222 128218 487404 128454
rect 486804 128134 487404 128218
rect 486804 127898 486986 128134
rect 487222 127898 487404 128134
rect 486804 92454 487404 127898
rect 486804 92218 486986 92454
rect 487222 92218 487404 92454
rect 486804 92134 487404 92218
rect 486804 91898 486986 92134
rect 487222 91898 487404 92134
rect 486804 56454 487404 91898
rect 486804 56218 486986 56454
rect 487222 56218 487404 56454
rect 486804 56134 487404 56218
rect 486804 55898 486986 56134
rect 487222 55898 487404 56134
rect 486804 20454 487404 55898
rect 486804 20218 486986 20454
rect 487222 20218 487404 20454
rect 486804 20134 487404 20218
rect 486804 19898 486986 20134
rect 487222 19898 487404 20134
rect 486804 -1266 487404 19898
rect 486804 -1502 486986 -1266
rect 487222 -1502 487404 -1266
rect 486804 -1586 487404 -1502
rect 486804 -1822 486986 -1586
rect 487222 -1822 487404 -1586
rect 486804 -1844 487404 -1822
rect 490404 672054 491004 707042
rect 490404 671818 490586 672054
rect 490822 671818 491004 672054
rect 490404 671734 491004 671818
rect 490404 671498 490586 671734
rect 490822 671498 491004 671734
rect 490404 636054 491004 671498
rect 490404 635818 490586 636054
rect 490822 635818 491004 636054
rect 490404 635734 491004 635818
rect 490404 635498 490586 635734
rect 490822 635498 491004 635734
rect 490404 600054 491004 635498
rect 490404 599818 490586 600054
rect 490822 599818 491004 600054
rect 490404 599734 491004 599818
rect 490404 599498 490586 599734
rect 490822 599498 491004 599734
rect 490404 564054 491004 599498
rect 490404 563818 490586 564054
rect 490822 563818 491004 564054
rect 490404 563734 491004 563818
rect 490404 563498 490586 563734
rect 490822 563498 491004 563734
rect 490404 528054 491004 563498
rect 490404 527818 490586 528054
rect 490822 527818 491004 528054
rect 490404 527734 491004 527818
rect 490404 527498 490586 527734
rect 490822 527498 491004 527734
rect 490404 492054 491004 527498
rect 490404 491818 490586 492054
rect 490822 491818 491004 492054
rect 490404 491734 491004 491818
rect 490404 491498 490586 491734
rect 490822 491498 491004 491734
rect 490404 456054 491004 491498
rect 490404 455818 490586 456054
rect 490822 455818 491004 456054
rect 490404 455734 491004 455818
rect 490404 455498 490586 455734
rect 490822 455498 491004 455734
rect 490404 420054 491004 455498
rect 490404 419818 490586 420054
rect 490822 419818 491004 420054
rect 490404 419734 491004 419818
rect 490404 419498 490586 419734
rect 490822 419498 491004 419734
rect 490404 384054 491004 419498
rect 490404 383818 490586 384054
rect 490822 383818 491004 384054
rect 490404 383734 491004 383818
rect 490404 383498 490586 383734
rect 490822 383498 491004 383734
rect 490404 348054 491004 383498
rect 490404 347818 490586 348054
rect 490822 347818 491004 348054
rect 490404 347734 491004 347818
rect 490404 347498 490586 347734
rect 490822 347498 491004 347734
rect 490404 312054 491004 347498
rect 490404 311818 490586 312054
rect 490822 311818 491004 312054
rect 490404 311734 491004 311818
rect 490404 311498 490586 311734
rect 490822 311498 491004 311734
rect 490404 276054 491004 311498
rect 490404 275818 490586 276054
rect 490822 275818 491004 276054
rect 490404 275734 491004 275818
rect 490404 275498 490586 275734
rect 490822 275498 491004 275734
rect 490404 240054 491004 275498
rect 490404 239818 490586 240054
rect 490822 239818 491004 240054
rect 490404 239734 491004 239818
rect 490404 239498 490586 239734
rect 490822 239498 491004 239734
rect 490404 204054 491004 239498
rect 490404 203818 490586 204054
rect 490822 203818 491004 204054
rect 490404 203734 491004 203818
rect 490404 203498 490586 203734
rect 490822 203498 491004 203734
rect 490404 168054 491004 203498
rect 490404 167818 490586 168054
rect 490822 167818 491004 168054
rect 490404 167734 491004 167818
rect 490404 167498 490586 167734
rect 490822 167498 491004 167734
rect 490404 132054 491004 167498
rect 490404 131818 490586 132054
rect 490822 131818 491004 132054
rect 490404 131734 491004 131818
rect 490404 131498 490586 131734
rect 490822 131498 491004 131734
rect 490404 96054 491004 131498
rect 490404 95818 490586 96054
rect 490822 95818 491004 96054
rect 490404 95734 491004 95818
rect 490404 95498 490586 95734
rect 490822 95498 491004 95734
rect 490404 60054 491004 95498
rect 490404 59818 490586 60054
rect 490822 59818 491004 60054
rect 490404 59734 491004 59818
rect 490404 59498 490586 59734
rect 490822 59498 491004 59734
rect 490404 24054 491004 59498
rect 490404 23818 490586 24054
rect 490822 23818 491004 24054
rect 490404 23734 491004 23818
rect 490404 23498 490586 23734
rect 490822 23498 491004 23734
rect 490404 -3106 491004 23498
rect 490404 -3342 490586 -3106
rect 490822 -3342 491004 -3106
rect 490404 -3426 491004 -3342
rect 490404 -3662 490586 -3426
rect 490822 -3662 491004 -3426
rect 490404 -3684 491004 -3662
rect 494004 675654 494604 708882
rect 494004 675418 494186 675654
rect 494422 675418 494604 675654
rect 494004 675334 494604 675418
rect 494004 675098 494186 675334
rect 494422 675098 494604 675334
rect 494004 639654 494604 675098
rect 494004 639418 494186 639654
rect 494422 639418 494604 639654
rect 494004 639334 494604 639418
rect 494004 639098 494186 639334
rect 494422 639098 494604 639334
rect 494004 603654 494604 639098
rect 494004 603418 494186 603654
rect 494422 603418 494604 603654
rect 494004 603334 494604 603418
rect 494004 603098 494186 603334
rect 494422 603098 494604 603334
rect 494004 567654 494604 603098
rect 494004 567418 494186 567654
rect 494422 567418 494604 567654
rect 494004 567334 494604 567418
rect 494004 567098 494186 567334
rect 494422 567098 494604 567334
rect 494004 531654 494604 567098
rect 494004 531418 494186 531654
rect 494422 531418 494604 531654
rect 494004 531334 494604 531418
rect 494004 531098 494186 531334
rect 494422 531098 494604 531334
rect 494004 495654 494604 531098
rect 494004 495418 494186 495654
rect 494422 495418 494604 495654
rect 494004 495334 494604 495418
rect 494004 495098 494186 495334
rect 494422 495098 494604 495334
rect 494004 459654 494604 495098
rect 494004 459418 494186 459654
rect 494422 459418 494604 459654
rect 494004 459334 494604 459418
rect 494004 459098 494186 459334
rect 494422 459098 494604 459334
rect 494004 423654 494604 459098
rect 494004 423418 494186 423654
rect 494422 423418 494604 423654
rect 494004 423334 494604 423418
rect 494004 423098 494186 423334
rect 494422 423098 494604 423334
rect 494004 387654 494604 423098
rect 494004 387418 494186 387654
rect 494422 387418 494604 387654
rect 494004 387334 494604 387418
rect 494004 387098 494186 387334
rect 494422 387098 494604 387334
rect 494004 351654 494604 387098
rect 494004 351418 494186 351654
rect 494422 351418 494604 351654
rect 494004 351334 494604 351418
rect 494004 351098 494186 351334
rect 494422 351098 494604 351334
rect 494004 315654 494604 351098
rect 494004 315418 494186 315654
rect 494422 315418 494604 315654
rect 494004 315334 494604 315418
rect 494004 315098 494186 315334
rect 494422 315098 494604 315334
rect 494004 279654 494604 315098
rect 494004 279418 494186 279654
rect 494422 279418 494604 279654
rect 494004 279334 494604 279418
rect 494004 279098 494186 279334
rect 494422 279098 494604 279334
rect 494004 243654 494604 279098
rect 494004 243418 494186 243654
rect 494422 243418 494604 243654
rect 494004 243334 494604 243418
rect 494004 243098 494186 243334
rect 494422 243098 494604 243334
rect 494004 207654 494604 243098
rect 494004 207418 494186 207654
rect 494422 207418 494604 207654
rect 494004 207334 494604 207418
rect 494004 207098 494186 207334
rect 494422 207098 494604 207334
rect 494004 171654 494604 207098
rect 494004 171418 494186 171654
rect 494422 171418 494604 171654
rect 494004 171334 494604 171418
rect 494004 171098 494186 171334
rect 494422 171098 494604 171334
rect 494004 135654 494604 171098
rect 494004 135418 494186 135654
rect 494422 135418 494604 135654
rect 494004 135334 494604 135418
rect 494004 135098 494186 135334
rect 494422 135098 494604 135334
rect 494004 99654 494604 135098
rect 494004 99418 494186 99654
rect 494422 99418 494604 99654
rect 494004 99334 494604 99418
rect 494004 99098 494186 99334
rect 494422 99098 494604 99334
rect 494004 63654 494604 99098
rect 494004 63418 494186 63654
rect 494422 63418 494604 63654
rect 494004 63334 494604 63418
rect 494004 63098 494186 63334
rect 494422 63098 494604 63334
rect 494004 27654 494604 63098
rect 494004 27418 494186 27654
rect 494422 27418 494604 27654
rect 494004 27334 494604 27418
rect 494004 27098 494186 27334
rect 494422 27098 494604 27334
rect 494004 -4946 494604 27098
rect 494004 -5182 494186 -4946
rect 494422 -5182 494604 -4946
rect 494004 -5266 494604 -5182
rect 494004 -5502 494186 -5266
rect 494422 -5502 494604 -5266
rect 494004 -5524 494604 -5502
rect 497604 679254 498204 710722
rect 515604 710358 516204 711300
rect 515604 710122 515786 710358
rect 516022 710122 516204 710358
rect 515604 710038 516204 710122
rect 515604 709802 515786 710038
rect 516022 709802 516204 710038
rect 512004 708518 512604 709460
rect 512004 708282 512186 708518
rect 512422 708282 512604 708518
rect 512004 708198 512604 708282
rect 512004 707962 512186 708198
rect 512422 707962 512604 708198
rect 508404 706678 509004 707620
rect 508404 706442 508586 706678
rect 508822 706442 509004 706678
rect 508404 706358 509004 706442
rect 508404 706122 508586 706358
rect 508822 706122 509004 706358
rect 497604 679018 497786 679254
rect 498022 679018 498204 679254
rect 497604 678934 498204 679018
rect 497604 678698 497786 678934
rect 498022 678698 498204 678934
rect 497604 643254 498204 678698
rect 497604 643018 497786 643254
rect 498022 643018 498204 643254
rect 497604 642934 498204 643018
rect 497604 642698 497786 642934
rect 498022 642698 498204 642934
rect 497604 607254 498204 642698
rect 497604 607018 497786 607254
rect 498022 607018 498204 607254
rect 497604 606934 498204 607018
rect 497604 606698 497786 606934
rect 498022 606698 498204 606934
rect 497604 571254 498204 606698
rect 497604 571018 497786 571254
rect 498022 571018 498204 571254
rect 497604 570934 498204 571018
rect 497604 570698 497786 570934
rect 498022 570698 498204 570934
rect 497604 535254 498204 570698
rect 497604 535018 497786 535254
rect 498022 535018 498204 535254
rect 497604 534934 498204 535018
rect 497604 534698 497786 534934
rect 498022 534698 498204 534934
rect 497604 499254 498204 534698
rect 497604 499018 497786 499254
rect 498022 499018 498204 499254
rect 497604 498934 498204 499018
rect 497604 498698 497786 498934
rect 498022 498698 498204 498934
rect 497604 463254 498204 498698
rect 497604 463018 497786 463254
rect 498022 463018 498204 463254
rect 497604 462934 498204 463018
rect 497604 462698 497786 462934
rect 498022 462698 498204 462934
rect 497604 427254 498204 462698
rect 497604 427018 497786 427254
rect 498022 427018 498204 427254
rect 497604 426934 498204 427018
rect 497604 426698 497786 426934
rect 498022 426698 498204 426934
rect 497604 391254 498204 426698
rect 497604 391018 497786 391254
rect 498022 391018 498204 391254
rect 497604 390934 498204 391018
rect 497604 390698 497786 390934
rect 498022 390698 498204 390934
rect 497604 355254 498204 390698
rect 497604 355018 497786 355254
rect 498022 355018 498204 355254
rect 497604 354934 498204 355018
rect 497604 354698 497786 354934
rect 498022 354698 498204 354934
rect 497604 319254 498204 354698
rect 497604 319018 497786 319254
rect 498022 319018 498204 319254
rect 497604 318934 498204 319018
rect 497604 318698 497786 318934
rect 498022 318698 498204 318934
rect 497604 283254 498204 318698
rect 497604 283018 497786 283254
rect 498022 283018 498204 283254
rect 497604 282934 498204 283018
rect 497604 282698 497786 282934
rect 498022 282698 498204 282934
rect 497604 247254 498204 282698
rect 497604 247018 497786 247254
rect 498022 247018 498204 247254
rect 497604 246934 498204 247018
rect 497604 246698 497786 246934
rect 498022 246698 498204 246934
rect 497604 211254 498204 246698
rect 497604 211018 497786 211254
rect 498022 211018 498204 211254
rect 497604 210934 498204 211018
rect 497604 210698 497786 210934
rect 498022 210698 498204 210934
rect 497604 175254 498204 210698
rect 497604 175018 497786 175254
rect 498022 175018 498204 175254
rect 497604 174934 498204 175018
rect 497604 174698 497786 174934
rect 498022 174698 498204 174934
rect 497604 139254 498204 174698
rect 497604 139018 497786 139254
rect 498022 139018 498204 139254
rect 497604 138934 498204 139018
rect 497604 138698 497786 138934
rect 498022 138698 498204 138934
rect 497604 103254 498204 138698
rect 497604 103018 497786 103254
rect 498022 103018 498204 103254
rect 497604 102934 498204 103018
rect 497604 102698 497786 102934
rect 498022 102698 498204 102934
rect 497604 67254 498204 102698
rect 497604 67018 497786 67254
rect 498022 67018 498204 67254
rect 497604 66934 498204 67018
rect 497604 66698 497786 66934
rect 498022 66698 498204 66934
rect 497604 31254 498204 66698
rect 497604 31018 497786 31254
rect 498022 31018 498204 31254
rect 497604 30934 498204 31018
rect 497604 30698 497786 30934
rect 498022 30698 498204 30934
rect 479604 -6102 479786 -5866
rect 480022 -6102 480204 -5866
rect 479604 -6186 480204 -6102
rect 479604 -6422 479786 -6186
rect 480022 -6422 480204 -6186
rect 479604 -7364 480204 -6422
rect 497604 -6786 498204 30698
rect 504804 704838 505404 705780
rect 504804 704602 504986 704838
rect 505222 704602 505404 704838
rect 504804 704518 505404 704602
rect 504804 704282 504986 704518
rect 505222 704282 505404 704518
rect 504804 686454 505404 704282
rect 504804 686218 504986 686454
rect 505222 686218 505404 686454
rect 504804 686134 505404 686218
rect 504804 685898 504986 686134
rect 505222 685898 505404 686134
rect 504804 650454 505404 685898
rect 504804 650218 504986 650454
rect 505222 650218 505404 650454
rect 504804 650134 505404 650218
rect 504804 649898 504986 650134
rect 505222 649898 505404 650134
rect 504804 614454 505404 649898
rect 504804 614218 504986 614454
rect 505222 614218 505404 614454
rect 504804 614134 505404 614218
rect 504804 613898 504986 614134
rect 505222 613898 505404 614134
rect 504804 578454 505404 613898
rect 504804 578218 504986 578454
rect 505222 578218 505404 578454
rect 504804 578134 505404 578218
rect 504804 577898 504986 578134
rect 505222 577898 505404 578134
rect 504804 542454 505404 577898
rect 504804 542218 504986 542454
rect 505222 542218 505404 542454
rect 504804 542134 505404 542218
rect 504804 541898 504986 542134
rect 505222 541898 505404 542134
rect 504804 506454 505404 541898
rect 504804 506218 504986 506454
rect 505222 506218 505404 506454
rect 504804 506134 505404 506218
rect 504804 505898 504986 506134
rect 505222 505898 505404 506134
rect 504804 470454 505404 505898
rect 504804 470218 504986 470454
rect 505222 470218 505404 470454
rect 504804 470134 505404 470218
rect 504804 469898 504986 470134
rect 505222 469898 505404 470134
rect 504804 434454 505404 469898
rect 504804 434218 504986 434454
rect 505222 434218 505404 434454
rect 504804 434134 505404 434218
rect 504804 433898 504986 434134
rect 505222 433898 505404 434134
rect 504804 398454 505404 433898
rect 504804 398218 504986 398454
rect 505222 398218 505404 398454
rect 504804 398134 505404 398218
rect 504804 397898 504986 398134
rect 505222 397898 505404 398134
rect 504804 362454 505404 397898
rect 504804 362218 504986 362454
rect 505222 362218 505404 362454
rect 504804 362134 505404 362218
rect 504804 361898 504986 362134
rect 505222 361898 505404 362134
rect 504804 326454 505404 361898
rect 504804 326218 504986 326454
rect 505222 326218 505404 326454
rect 504804 326134 505404 326218
rect 504804 325898 504986 326134
rect 505222 325898 505404 326134
rect 504804 290454 505404 325898
rect 504804 290218 504986 290454
rect 505222 290218 505404 290454
rect 504804 290134 505404 290218
rect 504804 289898 504986 290134
rect 505222 289898 505404 290134
rect 504804 254454 505404 289898
rect 504804 254218 504986 254454
rect 505222 254218 505404 254454
rect 504804 254134 505404 254218
rect 504804 253898 504986 254134
rect 505222 253898 505404 254134
rect 504804 218454 505404 253898
rect 504804 218218 504986 218454
rect 505222 218218 505404 218454
rect 504804 218134 505404 218218
rect 504804 217898 504986 218134
rect 505222 217898 505404 218134
rect 504804 182454 505404 217898
rect 504804 182218 504986 182454
rect 505222 182218 505404 182454
rect 504804 182134 505404 182218
rect 504804 181898 504986 182134
rect 505222 181898 505404 182134
rect 504804 146454 505404 181898
rect 504804 146218 504986 146454
rect 505222 146218 505404 146454
rect 504804 146134 505404 146218
rect 504804 145898 504986 146134
rect 505222 145898 505404 146134
rect 504804 110454 505404 145898
rect 504804 110218 504986 110454
rect 505222 110218 505404 110454
rect 504804 110134 505404 110218
rect 504804 109898 504986 110134
rect 505222 109898 505404 110134
rect 504804 74454 505404 109898
rect 504804 74218 504986 74454
rect 505222 74218 505404 74454
rect 504804 74134 505404 74218
rect 504804 73898 504986 74134
rect 505222 73898 505404 74134
rect 504804 38454 505404 73898
rect 504804 38218 504986 38454
rect 505222 38218 505404 38454
rect 504804 38134 505404 38218
rect 504804 37898 504986 38134
rect 505222 37898 505404 38134
rect 504804 2454 505404 37898
rect 504804 2218 504986 2454
rect 505222 2218 505404 2454
rect 504804 2134 505404 2218
rect 504804 1898 504986 2134
rect 505222 1898 505404 2134
rect 504804 -346 505404 1898
rect 504804 -582 504986 -346
rect 505222 -582 505404 -346
rect 504804 -666 505404 -582
rect 504804 -902 504986 -666
rect 505222 -902 505404 -666
rect 504804 -1844 505404 -902
rect 508404 690054 509004 706122
rect 508404 689818 508586 690054
rect 508822 689818 509004 690054
rect 508404 689734 509004 689818
rect 508404 689498 508586 689734
rect 508822 689498 509004 689734
rect 508404 654054 509004 689498
rect 508404 653818 508586 654054
rect 508822 653818 509004 654054
rect 508404 653734 509004 653818
rect 508404 653498 508586 653734
rect 508822 653498 509004 653734
rect 508404 618054 509004 653498
rect 508404 617818 508586 618054
rect 508822 617818 509004 618054
rect 508404 617734 509004 617818
rect 508404 617498 508586 617734
rect 508822 617498 509004 617734
rect 508404 582054 509004 617498
rect 508404 581818 508586 582054
rect 508822 581818 509004 582054
rect 508404 581734 509004 581818
rect 508404 581498 508586 581734
rect 508822 581498 509004 581734
rect 508404 546054 509004 581498
rect 508404 545818 508586 546054
rect 508822 545818 509004 546054
rect 508404 545734 509004 545818
rect 508404 545498 508586 545734
rect 508822 545498 509004 545734
rect 508404 510054 509004 545498
rect 508404 509818 508586 510054
rect 508822 509818 509004 510054
rect 508404 509734 509004 509818
rect 508404 509498 508586 509734
rect 508822 509498 509004 509734
rect 508404 474054 509004 509498
rect 508404 473818 508586 474054
rect 508822 473818 509004 474054
rect 508404 473734 509004 473818
rect 508404 473498 508586 473734
rect 508822 473498 509004 473734
rect 508404 438054 509004 473498
rect 508404 437818 508586 438054
rect 508822 437818 509004 438054
rect 508404 437734 509004 437818
rect 508404 437498 508586 437734
rect 508822 437498 509004 437734
rect 508404 402054 509004 437498
rect 508404 401818 508586 402054
rect 508822 401818 509004 402054
rect 508404 401734 509004 401818
rect 508404 401498 508586 401734
rect 508822 401498 509004 401734
rect 508404 366054 509004 401498
rect 508404 365818 508586 366054
rect 508822 365818 509004 366054
rect 508404 365734 509004 365818
rect 508404 365498 508586 365734
rect 508822 365498 509004 365734
rect 508404 330054 509004 365498
rect 508404 329818 508586 330054
rect 508822 329818 509004 330054
rect 508404 329734 509004 329818
rect 508404 329498 508586 329734
rect 508822 329498 509004 329734
rect 508404 294054 509004 329498
rect 508404 293818 508586 294054
rect 508822 293818 509004 294054
rect 508404 293734 509004 293818
rect 508404 293498 508586 293734
rect 508822 293498 509004 293734
rect 508404 258054 509004 293498
rect 508404 257818 508586 258054
rect 508822 257818 509004 258054
rect 508404 257734 509004 257818
rect 508404 257498 508586 257734
rect 508822 257498 509004 257734
rect 508404 222054 509004 257498
rect 508404 221818 508586 222054
rect 508822 221818 509004 222054
rect 508404 221734 509004 221818
rect 508404 221498 508586 221734
rect 508822 221498 509004 221734
rect 508404 186054 509004 221498
rect 508404 185818 508586 186054
rect 508822 185818 509004 186054
rect 508404 185734 509004 185818
rect 508404 185498 508586 185734
rect 508822 185498 509004 185734
rect 508404 150054 509004 185498
rect 508404 149818 508586 150054
rect 508822 149818 509004 150054
rect 508404 149734 509004 149818
rect 508404 149498 508586 149734
rect 508822 149498 509004 149734
rect 508404 114054 509004 149498
rect 508404 113818 508586 114054
rect 508822 113818 509004 114054
rect 508404 113734 509004 113818
rect 508404 113498 508586 113734
rect 508822 113498 509004 113734
rect 508404 78054 509004 113498
rect 508404 77818 508586 78054
rect 508822 77818 509004 78054
rect 508404 77734 509004 77818
rect 508404 77498 508586 77734
rect 508822 77498 509004 77734
rect 508404 42054 509004 77498
rect 508404 41818 508586 42054
rect 508822 41818 509004 42054
rect 508404 41734 509004 41818
rect 508404 41498 508586 41734
rect 508822 41498 509004 41734
rect 508404 6054 509004 41498
rect 508404 5818 508586 6054
rect 508822 5818 509004 6054
rect 508404 5734 509004 5818
rect 508404 5498 508586 5734
rect 508822 5498 509004 5734
rect 508404 -2186 509004 5498
rect 508404 -2422 508586 -2186
rect 508822 -2422 509004 -2186
rect 508404 -2506 509004 -2422
rect 508404 -2742 508586 -2506
rect 508822 -2742 509004 -2506
rect 508404 -3684 509004 -2742
rect 512004 693654 512604 707962
rect 512004 693418 512186 693654
rect 512422 693418 512604 693654
rect 512004 693334 512604 693418
rect 512004 693098 512186 693334
rect 512422 693098 512604 693334
rect 512004 657654 512604 693098
rect 512004 657418 512186 657654
rect 512422 657418 512604 657654
rect 512004 657334 512604 657418
rect 512004 657098 512186 657334
rect 512422 657098 512604 657334
rect 512004 621654 512604 657098
rect 512004 621418 512186 621654
rect 512422 621418 512604 621654
rect 512004 621334 512604 621418
rect 512004 621098 512186 621334
rect 512422 621098 512604 621334
rect 512004 585654 512604 621098
rect 512004 585418 512186 585654
rect 512422 585418 512604 585654
rect 512004 585334 512604 585418
rect 512004 585098 512186 585334
rect 512422 585098 512604 585334
rect 512004 549654 512604 585098
rect 512004 549418 512186 549654
rect 512422 549418 512604 549654
rect 512004 549334 512604 549418
rect 512004 549098 512186 549334
rect 512422 549098 512604 549334
rect 512004 513654 512604 549098
rect 512004 513418 512186 513654
rect 512422 513418 512604 513654
rect 512004 513334 512604 513418
rect 512004 513098 512186 513334
rect 512422 513098 512604 513334
rect 512004 477654 512604 513098
rect 512004 477418 512186 477654
rect 512422 477418 512604 477654
rect 512004 477334 512604 477418
rect 512004 477098 512186 477334
rect 512422 477098 512604 477334
rect 512004 441654 512604 477098
rect 512004 441418 512186 441654
rect 512422 441418 512604 441654
rect 512004 441334 512604 441418
rect 512004 441098 512186 441334
rect 512422 441098 512604 441334
rect 512004 405654 512604 441098
rect 512004 405418 512186 405654
rect 512422 405418 512604 405654
rect 512004 405334 512604 405418
rect 512004 405098 512186 405334
rect 512422 405098 512604 405334
rect 512004 369654 512604 405098
rect 512004 369418 512186 369654
rect 512422 369418 512604 369654
rect 512004 369334 512604 369418
rect 512004 369098 512186 369334
rect 512422 369098 512604 369334
rect 512004 333654 512604 369098
rect 512004 333418 512186 333654
rect 512422 333418 512604 333654
rect 512004 333334 512604 333418
rect 512004 333098 512186 333334
rect 512422 333098 512604 333334
rect 512004 297654 512604 333098
rect 512004 297418 512186 297654
rect 512422 297418 512604 297654
rect 512004 297334 512604 297418
rect 512004 297098 512186 297334
rect 512422 297098 512604 297334
rect 512004 261654 512604 297098
rect 512004 261418 512186 261654
rect 512422 261418 512604 261654
rect 512004 261334 512604 261418
rect 512004 261098 512186 261334
rect 512422 261098 512604 261334
rect 512004 225654 512604 261098
rect 512004 225418 512186 225654
rect 512422 225418 512604 225654
rect 512004 225334 512604 225418
rect 512004 225098 512186 225334
rect 512422 225098 512604 225334
rect 512004 189654 512604 225098
rect 512004 189418 512186 189654
rect 512422 189418 512604 189654
rect 512004 189334 512604 189418
rect 512004 189098 512186 189334
rect 512422 189098 512604 189334
rect 512004 153654 512604 189098
rect 512004 153418 512186 153654
rect 512422 153418 512604 153654
rect 512004 153334 512604 153418
rect 512004 153098 512186 153334
rect 512422 153098 512604 153334
rect 512004 117654 512604 153098
rect 512004 117418 512186 117654
rect 512422 117418 512604 117654
rect 512004 117334 512604 117418
rect 512004 117098 512186 117334
rect 512422 117098 512604 117334
rect 512004 81654 512604 117098
rect 512004 81418 512186 81654
rect 512422 81418 512604 81654
rect 512004 81334 512604 81418
rect 512004 81098 512186 81334
rect 512422 81098 512604 81334
rect 512004 45654 512604 81098
rect 512004 45418 512186 45654
rect 512422 45418 512604 45654
rect 512004 45334 512604 45418
rect 512004 45098 512186 45334
rect 512422 45098 512604 45334
rect 512004 9654 512604 45098
rect 512004 9418 512186 9654
rect 512422 9418 512604 9654
rect 512004 9334 512604 9418
rect 512004 9098 512186 9334
rect 512422 9098 512604 9334
rect 512004 -4026 512604 9098
rect 512004 -4262 512186 -4026
rect 512422 -4262 512604 -4026
rect 512004 -4346 512604 -4262
rect 512004 -4582 512186 -4346
rect 512422 -4582 512604 -4346
rect 512004 -5524 512604 -4582
rect 515604 697254 516204 709802
rect 533604 711278 534204 711300
rect 533604 711042 533786 711278
rect 534022 711042 534204 711278
rect 533604 710958 534204 711042
rect 533604 710722 533786 710958
rect 534022 710722 534204 710958
rect 530004 709438 530604 709460
rect 530004 709202 530186 709438
rect 530422 709202 530604 709438
rect 530004 709118 530604 709202
rect 530004 708882 530186 709118
rect 530422 708882 530604 709118
rect 526404 707598 527004 707620
rect 526404 707362 526586 707598
rect 526822 707362 527004 707598
rect 526404 707278 527004 707362
rect 526404 707042 526586 707278
rect 526822 707042 527004 707278
rect 515604 697018 515786 697254
rect 516022 697018 516204 697254
rect 515604 696934 516204 697018
rect 515604 696698 515786 696934
rect 516022 696698 516204 696934
rect 515604 661254 516204 696698
rect 515604 661018 515786 661254
rect 516022 661018 516204 661254
rect 515604 660934 516204 661018
rect 515604 660698 515786 660934
rect 516022 660698 516204 660934
rect 515604 625254 516204 660698
rect 515604 625018 515786 625254
rect 516022 625018 516204 625254
rect 515604 624934 516204 625018
rect 515604 624698 515786 624934
rect 516022 624698 516204 624934
rect 515604 589254 516204 624698
rect 515604 589018 515786 589254
rect 516022 589018 516204 589254
rect 515604 588934 516204 589018
rect 515604 588698 515786 588934
rect 516022 588698 516204 588934
rect 515604 553254 516204 588698
rect 515604 553018 515786 553254
rect 516022 553018 516204 553254
rect 515604 552934 516204 553018
rect 515604 552698 515786 552934
rect 516022 552698 516204 552934
rect 515604 517254 516204 552698
rect 515604 517018 515786 517254
rect 516022 517018 516204 517254
rect 515604 516934 516204 517018
rect 515604 516698 515786 516934
rect 516022 516698 516204 516934
rect 515604 481254 516204 516698
rect 515604 481018 515786 481254
rect 516022 481018 516204 481254
rect 515604 480934 516204 481018
rect 515604 480698 515786 480934
rect 516022 480698 516204 480934
rect 515604 445254 516204 480698
rect 515604 445018 515786 445254
rect 516022 445018 516204 445254
rect 515604 444934 516204 445018
rect 515604 444698 515786 444934
rect 516022 444698 516204 444934
rect 515604 409254 516204 444698
rect 515604 409018 515786 409254
rect 516022 409018 516204 409254
rect 515604 408934 516204 409018
rect 515604 408698 515786 408934
rect 516022 408698 516204 408934
rect 515604 373254 516204 408698
rect 515604 373018 515786 373254
rect 516022 373018 516204 373254
rect 515604 372934 516204 373018
rect 515604 372698 515786 372934
rect 516022 372698 516204 372934
rect 515604 337254 516204 372698
rect 515604 337018 515786 337254
rect 516022 337018 516204 337254
rect 515604 336934 516204 337018
rect 515604 336698 515786 336934
rect 516022 336698 516204 336934
rect 515604 301254 516204 336698
rect 515604 301018 515786 301254
rect 516022 301018 516204 301254
rect 515604 300934 516204 301018
rect 515604 300698 515786 300934
rect 516022 300698 516204 300934
rect 515604 265254 516204 300698
rect 515604 265018 515786 265254
rect 516022 265018 516204 265254
rect 515604 264934 516204 265018
rect 515604 264698 515786 264934
rect 516022 264698 516204 264934
rect 515604 229254 516204 264698
rect 515604 229018 515786 229254
rect 516022 229018 516204 229254
rect 515604 228934 516204 229018
rect 515604 228698 515786 228934
rect 516022 228698 516204 228934
rect 515604 193254 516204 228698
rect 515604 193018 515786 193254
rect 516022 193018 516204 193254
rect 515604 192934 516204 193018
rect 515604 192698 515786 192934
rect 516022 192698 516204 192934
rect 515604 157254 516204 192698
rect 515604 157018 515786 157254
rect 516022 157018 516204 157254
rect 515604 156934 516204 157018
rect 515604 156698 515786 156934
rect 516022 156698 516204 156934
rect 515604 121254 516204 156698
rect 515604 121018 515786 121254
rect 516022 121018 516204 121254
rect 515604 120934 516204 121018
rect 515604 120698 515786 120934
rect 516022 120698 516204 120934
rect 515604 85254 516204 120698
rect 515604 85018 515786 85254
rect 516022 85018 516204 85254
rect 515604 84934 516204 85018
rect 515604 84698 515786 84934
rect 516022 84698 516204 84934
rect 515604 49254 516204 84698
rect 515604 49018 515786 49254
rect 516022 49018 516204 49254
rect 515604 48934 516204 49018
rect 515604 48698 515786 48934
rect 516022 48698 516204 48934
rect 515604 13254 516204 48698
rect 515604 13018 515786 13254
rect 516022 13018 516204 13254
rect 515604 12934 516204 13018
rect 515604 12698 515786 12934
rect 516022 12698 516204 12934
rect 497604 -7022 497786 -6786
rect 498022 -7022 498204 -6786
rect 497604 -7106 498204 -7022
rect 497604 -7342 497786 -7106
rect 498022 -7342 498204 -7106
rect 497604 -7364 498204 -7342
rect 515604 -5866 516204 12698
rect 522804 705758 523404 705780
rect 522804 705522 522986 705758
rect 523222 705522 523404 705758
rect 522804 705438 523404 705522
rect 522804 705202 522986 705438
rect 523222 705202 523404 705438
rect 522804 668454 523404 705202
rect 522804 668218 522986 668454
rect 523222 668218 523404 668454
rect 522804 668134 523404 668218
rect 522804 667898 522986 668134
rect 523222 667898 523404 668134
rect 522804 632454 523404 667898
rect 522804 632218 522986 632454
rect 523222 632218 523404 632454
rect 522804 632134 523404 632218
rect 522804 631898 522986 632134
rect 523222 631898 523404 632134
rect 522804 596454 523404 631898
rect 522804 596218 522986 596454
rect 523222 596218 523404 596454
rect 522804 596134 523404 596218
rect 522804 595898 522986 596134
rect 523222 595898 523404 596134
rect 522804 560454 523404 595898
rect 522804 560218 522986 560454
rect 523222 560218 523404 560454
rect 522804 560134 523404 560218
rect 522804 559898 522986 560134
rect 523222 559898 523404 560134
rect 522804 524454 523404 559898
rect 522804 524218 522986 524454
rect 523222 524218 523404 524454
rect 522804 524134 523404 524218
rect 522804 523898 522986 524134
rect 523222 523898 523404 524134
rect 522804 488454 523404 523898
rect 522804 488218 522986 488454
rect 523222 488218 523404 488454
rect 522804 488134 523404 488218
rect 522804 487898 522986 488134
rect 523222 487898 523404 488134
rect 522804 452454 523404 487898
rect 522804 452218 522986 452454
rect 523222 452218 523404 452454
rect 522804 452134 523404 452218
rect 522804 451898 522986 452134
rect 523222 451898 523404 452134
rect 522804 416454 523404 451898
rect 522804 416218 522986 416454
rect 523222 416218 523404 416454
rect 522804 416134 523404 416218
rect 522804 415898 522986 416134
rect 523222 415898 523404 416134
rect 522804 380454 523404 415898
rect 522804 380218 522986 380454
rect 523222 380218 523404 380454
rect 522804 380134 523404 380218
rect 522804 379898 522986 380134
rect 523222 379898 523404 380134
rect 522804 344454 523404 379898
rect 522804 344218 522986 344454
rect 523222 344218 523404 344454
rect 522804 344134 523404 344218
rect 522804 343898 522986 344134
rect 523222 343898 523404 344134
rect 522804 308454 523404 343898
rect 522804 308218 522986 308454
rect 523222 308218 523404 308454
rect 522804 308134 523404 308218
rect 522804 307898 522986 308134
rect 523222 307898 523404 308134
rect 522804 272454 523404 307898
rect 522804 272218 522986 272454
rect 523222 272218 523404 272454
rect 522804 272134 523404 272218
rect 522804 271898 522986 272134
rect 523222 271898 523404 272134
rect 522804 236454 523404 271898
rect 522804 236218 522986 236454
rect 523222 236218 523404 236454
rect 522804 236134 523404 236218
rect 522804 235898 522986 236134
rect 523222 235898 523404 236134
rect 522804 200454 523404 235898
rect 522804 200218 522986 200454
rect 523222 200218 523404 200454
rect 522804 200134 523404 200218
rect 522804 199898 522986 200134
rect 523222 199898 523404 200134
rect 522804 164454 523404 199898
rect 522804 164218 522986 164454
rect 523222 164218 523404 164454
rect 522804 164134 523404 164218
rect 522804 163898 522986 164134
rect 523222 163898 523404 164134
rect 522804 128454 523404 163898
rect 522804 128218 522986 128454
rect 523222 128218 523404 128454
rect 522804 128134 523404 128218
rect 522804 127898 522986 128134
rect 523222 127898 523404 128134
rect 522804 92454 523404 127898
rect 522804 92218 522986 92454
rect 523222 92218 523404 92454
rect 522804 92134 523404 92218
rect 522804 91898 522986 92134
rect 523222 91898 523404 92134
rect 522804 56454 523404 91898
rect 522804 56218 522986 56454
rect 523222 56218 523404 56454
rect 522804 56134 523404 56218
rect 522804 55898 522986 56134
rect 523222 55898 523404 56134
rect 522804 20454 523404 55898
rect 522804 20218 522986 20454
rect 523222 20218 523404 20454
rect 522804 20134 523404 20218
rect 522804 19898 522986 20134
rect 523222 19898 523404 20134
rect 522804 -1266 523404 19898
rect 522804 -1502 522986 -1266
rect 523222 -1502 523404 -1266
rect 522804 -1586 523404 -1502
rect 522804 -1822 522986 -1586
rect 523222 -1822 523404 -1586
rect 522804 -1844 523404 -1822
rect 526404 672054 527004 707042
rect 526404 671818 526586 672054
rect 526822 671818 527004 672054
rect 526404 671734 527004 671818
rect 526404 671498 526586 671734
rect 526822 671498 527004 671734
rect 526404 636054 527004 671498
rect 526404 635818 526586 636054
rect 526822 635818 527004 636054
rect 526404 635734 527004 635818
rect 526404 635498 526586 635734
rect 526822 635498 527004 635734
rect 526404 600054 527004 635498
rect 526404 599818 526586 600054
rect 526822 599818 527004 600054
rect 526404 599734 527004 599818
rect 526404 599498 526586 599734
rect 526822 599498 527004 599734
rect 526404 564054 527004 599498
rect 526404 563818 526586 564054
rect 526822 563818 527004 564054
rect 526404 563734 527004 563818
rect 526404 563498 526586 563734
rect 526822 563498 527004 563734
rect 526404 528054 527004 563498
rect 526404 527818 526586 528054
rect 526822 527818 527004 528054
rect 526404 527734 527004 527818
rect 526404 527498 526586 527734
rect 526822 527498 527004 527734
rect 526404 492054 527004 527498
rect 526404 491818 526586 492054
rect 526822 491818 527004 492054
rect 526404 491734 527004 491818
rect 526404 491498 526586 491734
rect 526822 491498 527004 491734
rect 526404 456054 527004 491498
rect 526404 455818 526586 456054
rect 526822 455818 527004 456054
rect 526404 455734 527004 455818
rect 526404 455498 526586 455734
rect 526822 455498 527004 455734
rect 526404 420054 527004 455498
rect 526404 419818 526586 420054
rect 526822 419818 527004 420054
rect 526404 419734 527004 419818
rect 526404 419498 526586 419734
rect 526822 419498 527004 419734
rect 526404 384054 527004 419498
rect 526404 383818 526586 384054
rect 526822 383818 527004 384054
rect 526404 383734 527004 383818
rect 526404 383498 526586 383734
rect 526822 383498 527004 383734
rect 526404 348054 527004 383498
rect 526404 347818 526586 348054
rect 526822 347818 527004 348054
rect 526404 347734 527004 347818
rect 526404 347498 526586 347734
rect 526822 347498 527004 347734
rect 526404 312054 527004 347498
rect 526404 311818 526586 312054
rect 526822 311818 527004 312054
rect 526404 311734 527004 311818
rect 526404 311498 526586 311734
rect 526822 311498 527004 311734
rect 526404 276054 527004 311498
rect 526404 275818 526586 276054
rect 526822 275818 527004 276054
rect 526404 275734 527004 275818
rect 526404 275498 526586 275734
rect 526822 275498 527004 275734
rect 526404 240054 527004 275498
rect 526404 239818 526586 240054
rect 526822 239818 527004 240054
rect 526404 239734 527004 239818
rect 526404 239498 526586 239734
rect 526822 239498 527004 239734
rect 526404 204054 527004 239498
rect 526404 203818 526586 204054
rect 526822 203818 527004 204054
rect 526404 203734 527004 203818
rect 526404 203498 526586 203734
rect 526822 203498 527004 203734
rect 526404 168054 527004 203498
rect 526404 167818 526586 168054
rect 526822 167818 527004 168054
rect 526404 167734 527004 167818
rect 526404 167498 526586 167734
rect 526822 167498 527004 167734
rect 526404 132054 527004 167498
rect 526404 131818 526586 132054
rect 526822 131818 527004 132054
rect 526404 131734 527004 131818
rect 526404 131498 526586 131734
rect 526822 131498 527004 131734
rect 526404 96054 527004 131498
rect 526404 95818 526586 96054
rect 526822 95818 527004 96054
rect 526404 95734 527004 95818
rect 526404 95498 526586 95734
rect 526822 95498 527004 95734
rect 526404 60054 527004 95498
rect 526404 59818 526586 60054
rect 526822 59818 527004 60054
rect 526404 59734 527004 59818
rect 526404 59498 526586 59734
rect 526822 59498 527004 59734
rect 526404 24054 527004 59498
rect 526404 23818 526586 24054
rect 526822 23818 527004 24054
rect 526404 23734 527004 23818
rect 526404 23498 526586 23734
rect 526822 23498 527004 23734
rect 526404 -3106 527004 23498
rect 526404 -3342 526586 -3106
rect 526822 -3342 527004 -3106
rect 526404 -3426 527004 -3342
rect 526404 -3662 526586 -3426
rect 526822 -3662 527004 -3426
rect 526404 -3684 527004 -3662
rect 530004 675654 530604 708882
rect 530004 675418 530186 675654
rect 530422 675418 530604 675654
rect 530004 675334 530604 675418
rect 530004 675098 530186 675334
rect 530422 675098 530604 675334
rect 530004 639654 530604 675098
rect 530004 639418 530186 639654
rect 530422 639418 530604 639654
rect 530004 639334 530604 639418
rect 530004 639098 530186 639334
rect 530422 639098 530604 639334
rect 530004 603654 530604 639098
rect 530004 603418 530186 603654
rect 530422 603418 530604 603654
rect 530004 603334 530604 603418
rect 530004 603098 530186 603334
rect 530422 603098 530604 603334
rect 530004 567654 530604 603098
rect 530004 567418 530186 567654
rect 530422 567418 530604 567654
rect 530004 567334 530604 567418
rect 530004 567098 530186 567334
rect 530422 567098 530604 567334
rect 530004 531654 530604 567098
rect 530004 531418 530186 531654
rect 530422 531418 530604 531654
rect 530004 531334 530604 531418
rect 530004 531098 530186 531334
rect 530422 531098 530604 531334
rect 530004 495654 530604 531098
rect 530004 495418 530186 495654
rect 530422 495418 530604 495654
rect 530004 495334 530604 495418
rect 530004 495098 530186 495334
rect 530422 495098 530604 495334
rect 530004 459654 530604 495098
rect 530004 459418 530186 459654
rect 530422 459418 530604 459654
rect 530004 459334 530604 459418
rect 530004 459098 530186 459334
rect 530422 459098 530604 459334
rect 530004 423654 530604 459098
rect 530004 423418 530186 423654
rect 530422 423418 530604 423654
rect 530004 423334 530604 423418
rect 530004 423098 530186 423334
rect 530422 423098 530604 423334
rect 530004 387654 530604 423098
rect 530004 387418 530186 387654
rect 530422 387418 530604 387654
rect 530004 387334 530604 387418
rect 530004 387098 530186 387334
rect 530422 387098 530604 387334
rect 530004 351654 530604 387098
rect 530004 351418 530186 351654
rect 530422 351418 530604 351654
rect 530004 351334 530604 351418
rect 530004 351098 530186 351334
rect 530422 351098 530604 351334
rect 530004 315654 530604 351098
rect 530004 315418 530186 315654
rect 530422 315418 530604 315654
rect 530004 315334 530604 315418
rect 530004 315098 530186 315334
rect 530422 315098 530604 315334
rect 530004 279654 530604 315098
rect 530004 279418 530186 279654
rect 530422 279418 530604 279654
rect 530004 279334 530604 279418
rect 530004 279098 530186 279334
rect 530422 279098 530604 279334
rect 530004 243654 530604 279098
rect 530004 243418 530186 243654
rect 530422 243418 530604 243654
rect 530004 243334 530604 243418
rect 530004 243098 530186 243334
rect 530422 243098 530604 243334
rect 530004 207654 530604 243098
rect 530004 207418 530186 207654
rect 530422 207418 530604 207654
rect 530004 207334 530604 207418
rect 530004 207098 530186 207334
rect 530422 207098 530604 207334
rect 530004 171654 530604 207098
rect 530004 171418 530186 171654
rect 530422 171418 530604 171654
rect 530004 171334 530604 171418
rect 530004 171098 530186 171334
rect 530422 171098 530604 171334
rect 530004 135654 530604 171098
rect 530004 135418 530186 135654
rect 530422 135418 530604 135654
rect 530004 135334 530604 135418
rect 530004 135098 530186 135334
rect 530422 135098 530604 135334
rect 530004 99654 530604 135098
rect 530004 99418 530186 99654
rect 530422 99418 530604 99654
rect 530004 99334 530604 99418
rect 530004 99098 530186 99334
rect 530422 99098 530604 99334
rect 530004 63654 530604 99098
rect 530004 63418 530186 63654
rect 530422 63418 530604 63654
rect 530004 63334 530604 63418
rect 530004 63098 530186 63334
rect 530422 63098 530604 63334
rect 530004 27654 530604 63098
rect 530004 27418 530186 27654
rect 530422 27418 530604 27654
rect 530004 27334 530604 27418
rect 530004 27098 530186 27334
rect 530422 27098 530604 27334
rect 530004 -4946 530604 27098
rect 530004 -5182 530186 -4946
rect 530422 -5182 530604 -4946
rect 530004 -5266 530604 -5182
rect 530004 -5502 530186 -5266
rect 530422 -5502 530604 -5266
rect 530004 -5524 530604 -5502
rect 533604 679254 534204 710722
rect 551604 710358 552204 711300
rect 551604 710122 551786 710358
rect 552022 710122 552204 710358
rect 551604 710038 552204 710122
rect 551604 709802 551786 710038
rect 552022 709802 552204 710038
rect 548004 708518 548604 709460
rect 548004 708282 548186 708518
rect 548422 708282 548604 708518
rect 548004 708198 548604 708282
rect 548004 707962 548186 708198
rect 548422 707962 548604 708198
rect 544404 706678 545004 707620
rect 544404 706442 544586 706678
rect 544822 706442 545004 706678
rect 544404 706358 545004 706442
rect 544404 706122 544586 706358
rect 544822 706122 545004 706358
rect 533604 679018 533786 679254
rect 534022 679018 534204 679254
rect 533604 678934 534204 679018
rect 533604 678698 533786 678934
rect 534022 678698 534204 678934
rect 533604 643254 534204 678698
rect 533604 643018 533786 643254
rect 534022 643018 534204 643254
rect 533604 642934 534204 643018
rect 533604 642698 533786 642934
rect 534022 642698 534204 642934
rect 533604 607254 534204 642698
rect 533604 607018 533786 607254
rect 534022 607018 534204 607254
rect 533604 606934 534204 607018
rect 533604 606698 533786 606934
rect 534022 606698 534204 606934
rect 533604 571254 534204 606698
rect 533604 571018 533786 571254
rect 534022 571018 534204 571254
rect 533604 570934 534204 571018
rect 533604 570698 533786 570934
rect 534022 570698 534204 570934
rect 533604 535254 534204 570698
rect 533604 535018 533786 535254
rect 534022 535018 534204 535254
rect 533604 534934 534204 535018
rect 533604 534698 533786 534934
rect 534022 534698 534204 534934
rect 533604 499254 534204 534698
rect 533604 499018 533786 499254
rect 534022 499018 534204 499254
rect 533604 498934 534204 499018
rect 533604 498698 533786 498934
rect 534022 498698 534204 498934
rect 533604 463254 534204 498698
rect 533604 463018 533786 463254
rect 534022 463018 534204 463254
rect 533604 462934 534204 463018
rect 533604 462698 533786 462934
rect 534022 462698 534204 462934
rect 533604 427254 534204 462698
rect 533604 427018 533786 427254
rect 534022 427018 534204 427254
rect 533604 426934 534204 427018
rect 533604 426698 533786 426934
rect 534022 426698 534204 426934
rect 533604 391254 534204 426698
rect 533604 391018 533786 391254
rect 534022 391018 534204 391254
rect 533604 390934 534204 391018
rect 533604 390698 533786 390934
rect 534022 390698 534204 390934
rect 533604 355254 534204 390698
rect 533604 355018 533786 355254
rect 534022 355018 534204 355254
rect 533604 354934 534204 355018
rect 533604 354698 533786 354934
rect 534022 354698 534204 354934
rect 533604 319254 534204 354698
rect 533604 319018 533786 319254
rect 534022 319018 534204 319254
rect 533604 318934 534204 319018
rect 533604 318698 533786 318934
rect 534022 318698 534204 318934
rect 533604 283254 534204 318698
rect 533604 283018 533786 283254
rect 534022 283018 534204 283254
rect 533604 282934 534204 283018
rect 533604 282698 533786 282934
rect 534022 282698 534204 282934
rect 533604 247254 534204 282698
rect 533604 247018 533786 247254
rect 534022 247018 534204 247254
rect 533604 246934 534204 247018
rect 533604 246698 533786 246934
rect 534022 246698 534204 246934
rect 533604 211254 534204 246698
rect 533604 211018 533786 211254
rect 534022 211018 534204 211254
rect 533604 210934 534204 211018
rect 533604 210698 533786 210934
rect 534022 210698 534204 210934
rect 533604 175254 534204 210698
rect 533604 175018 533786 175254
rect 534022 175018 534204 175254
rect 533604 174934 534204 175018
rect 533604 174698 533786 174934
rect 534022 174698 534204 174934
rect 533604 139254 534204 174698
rect 533604 139018 533786 139254
rect 534022 139018 534204 139254
rect 533604 138934 534204 139018
rect 533604 138698 533786 138934
rect 534022 138698 534204 138934
rect 533604 103254 534204 138698
rect 533604 103018 533786 103254
rect 534022 103018 534204 103254
rect 533604 102934 534204 103018
rect 533604 102698 533786 102934
rect 534022 102698 534204 102934
rect 533604 67254 534204 102698
rect 533604 67018 533786 67254
rect 534022 67018 534204 67254
rect 533604 66934 534204 67018
rect 533604 66698 533786 66934
rect 534022 66698 534204 66934
rect 533604 31254 534204 66698
rect 533604 31018 533786 31254
rect 534022 31018 534204 31254
rect 533604 30934 534204 31018
rect 533604 30698 533786 30934
rect 534022 30698 534204 30934
rect 515604 -6102 515786 -5866
rect 516022 -6102 516204 -5866
rect 515604 -6186 516204 -6102
rect 515604 -6422 515786 -6186
rect 516022 -6422 516204 -6186
rect 515604 -7364 516204 -6422
rect 533604 -6786 534204 30698
rect 540804 704838 541404 705780
rect 540804 704602 540986 704838
rect 541222 704602 541404 704838
rect 540804 704518 541404 704602
rect 540804 704282 540986 704518
rect 541222 704282 541404 704518
rect 540804 686454 541404 704282
rect 540804 686218 540986 686454
rect 541222 686218 541404 686454
rect 540804 686134 541404 686218
rect 540804 685898 540986 686134
rect 541222 685898 541404 686134
rect 540804 650454 541404 685898
rect 540804 650218 540986 650454
rect 541222 650218 541404 650454
rect 540804 650134 541404 650218
rect 540804 649898 540986 650134
rect 541222 649898 541404 650134
rect 540804 614454 541404 649898
rect 540804 614218 540986 614454
rect 541222 614218 541404 614454
rect 540804 614134 541404 614218
rect 540804 613898 540986 614134
rect 541222 613898 541404 614134
rect 540804 578454 541404 613898
rect 540804 578218 540986 578454
rect 541222 578218 541404 578454
rect 540804 578134 541404 578218
rect 540804 577898 540986 578134
rect 541222 577898 541404 578134
rect 540804 542454 541404 577898
rect 540804 542218 540986 542454
rect 541222 542218 541404 542454
rect 540804 542134 541404 542218
rect 540804 541898 540986 542134
rect 541222 541898 541404 542134
rect 540804 506454 541404 541898
rect 540804 506218 540986 506454
rect 541222 506218 541404 506454
rect 540804 506134 541404 506218
rect 540804 505898 540986 506134
rect 541222 505898 541404 506134
rect 540804 470454 541404 505898
rect 540804 470218 540986 470454
rect 541222 470218 541404 470454
rect 540804 470134 541404 470218
rect 540804 469898 540986 470134
rect 541222 469898 541404 470134
rect 540804 434454 541404 469898
rect 540804 434218 540986 434454
rect 541222 434218 541404 434454
rect 540804 434134 541404 434218
rect 540804 433898 540986 434134
rect 541222 433898 541404 434134
rect 540804 398454 541404 433898
rect 540804 398218 540986 398454
rect 541222 398218 541404 398454
rect 540804 398134 541404 398218
rect 540804 397898 540986 398134
rect 541222 397898 541404 398134
rect 540804 362454 541404 397898
rect 540804 362218 540986 362454
rect 541222 362218 541404 362454
rect 540804 362134 541404 362218
rect 540804 361898 540986 362134
rect 541222 361898 541404 362134
rect 540804 326454 541404 361898
rect 540804 326218 540986 326454
rect 541222 326218 541404 326454
rect 540804 326134 541404 326218
rect 540804 325898 540986 326134
rect 541222 325898 541404 326134
rect 540804 290454 541404 325898
rect 540804 290218 540986 290454
rect 541222 290218 541404 290454
rect 540804 290134 541404 290218
rect 540804 289898 540986 290134
rect 541222 289898 541404 290134
rect 540804 254454 541404 289898
rect 540804 254218 540986 254454
rect 541222 254218 541404 254454
rect 540804 254134 541404 254218
rect 540804 253898 540986 254134
rect 541222 253898 541404 254134
rect 540804 218454 541404 253898
rect 540804 218218 540986 218454
rect 541222 218218 541404 218454
rect 540804 218134 541404 218218
rect 540804 217898 540986 218134
rect 541222 217898 541404 218134
rect 540804 182454 541404 217898
rect 540804 182218 540986 182454
rect 541222 182218 541404 182454
rect 540804 182134 541404 182218
rect 540804 181898 540986 182134
rect 541222 181898 541404 182134
rect 540804 146454 541404 181898
rect 540804 146218 540986 146454
rect 541222 146218 541404 146454
rect 540804 146134 541404 146218
rect 540804 145898 540986 146134
rect 541222 145898 541404 146134
rect 540804 110454 541404 145898
rect 540804 110218 540986 110454
rect 541222 110218 541404 110454
rect 540804 110134 541404 110218
rect 540804 109898 540986 110134
rect 541222 109898 541404 110134
rect 540804 74454 541404 109898
rect 540804 74218 540986 74454
rect 541222 74218 541404 74454
rect 540804 74134 541404 74218
rect 540804 73898 540986 74134
rect 541222 73898 541404 74134
rect 540804 38454 541404 73898
rect 540804 38218 540986 38454
rect 541222 38218 541404 38454
rect 540804 38134 541404 38218
rect 540804 37898 540986 38134
rect 541222 37898 541404 38134
rect 540804 2454 541404 37898
rect 540804 2218 540986 2454
rect 541222 2218 541404 2454
rect 540804 2134 541404 2218
rect 540804 1898 540986 2134
rect 541222 1898 541404 2134
rect 540804 -346 541404 1898
rect 540804 -582 540986 -346
rect 541222 -582 541404 -346
rect 540804 -666 541404 -582
rect 540804 -902 540986 -666
rect 541222 -902 541404 -666
rect 540804 -1844 541404 -902
rect 544404 690054 545004 706122
rect 544404 689818 544586 690054
rect 544822 689818 545004 690054
rect 544404 689734 545004 689818
rect 544404 689498 544586 689734
rect 544822 689498 545004 689734
rect 544404 654054 545004 689498
rect 544404 653818 544586 654054
rect 544822 653818 545004 654054
rect 544404 653734 545004 653818
rect 544404 653498 544586 653734
rect 544822 653498 545004 653734
rect 544404 618054 545004 653498
rect 544404 617818 544586 618054
rect 544822 617818 545004 618054
rect 544404 617734 545004 617818
rect 544404 617498 544586 617734
rect 544822 617498 545004 617734
rect 544404 582054 545004 617498
rect 544404 581818 544586 582054
rect 544822 581818 545004 582054
rect 544404 581734 545004 581818
rect 544404 581498 544586 581734
rect 544822 581498 545004 581734
rect 544404 546054 545004 581498
rect 544404 545818 544586 546054
rect 544822 545818 545004 546054
rect 544404 545734 545004 545818
rect 544404 545498 544586 545734
rect 544822 545498 545004 545734
rect 544404 510054 545004 545498
rect 544404 509818 544586 510054
rect 544822 509818 545004 510054
rect 544404 509734 545004 509818
rect 544404 509498 544586 509734
rect 544822 509498 545004 509734
rect 544404 474054 545004 509498
rect 544404 473818 544586 474054
rect 544822 473818 545004 474054
rect 544404 473734 545004 473818
rect 544404 473498 544586 473734
rect 544822 473498 545004 473734
rect 544404 438054 545004 473498
rect 544404 437818 544586 438054
rect 544822 437818 545004 438054
rect 544404 437734 545004 437818
rect 544404 437498 544586 437734
rect 544822 437498 545004 437734
rect 544404 402054 545004 437498
rect 544404 401818 544586 402054
rect 544822 401818 545004 402054
rect 544404 401734 545004 401818
rect 544404 401498 544586 401734
rect 544822 401498 545004 401734
rect 544404 366054 545004 401498
rect 544404 365818 544586 366054
rect 544822 365818 545004 366054
rect 544404 365734 545004 365818
rect 544404 365498 544586 365734
rect 544822 365498 545004 365734
rect 544404 330054 545004 365498
rect 544404 329818 544586 330054
rect 544822 329818 545004 330054
rect 544404 329734 545004 329818
rect 544404 329498 544586 329734
rect 544822 329498 545004 329734
rect 544404 294054 545004 329498
rect 544404 293818 544586 294054
rect 544822 293818 545004 294054
rect 544404 293734 545004 293818
rect 544404 293498 544586 293734
rect 544822 293498 545004 293734
rect 544404 258054 545004 293498
rect 544404 257818 544586 258054
rect 544822 257818 545004 258054
rect 544404 257734 545004 257818
rect 544404 257498 544586 257734
rect 544822 257498 545004 257734
rect 544404 222054 545004 257498
rect 544404 221818 544586 222054
rect 544822 221818 545004 222054
rect 544404 221734 545004 221818
rect 544404 221498 544586 221734
rect 544822 221498 545004 221734
rect 544404 186054 545004 221498
rect 544404 185818 544586 186054
rect 544822 185818 545004 186054
rect 544404 185734 545004 185818
rect 544404 185498 544586 185734
rect 544822 185498 545004 185734
rect 544404 150054 545004 185498
rect 544404 149818 544586 150054
rect 544822 149818 545004 150054
rect 544404 149734 545004 149818
rect 544404 149498 544586 149734
rect 544822 149498 545004 149734
rect 544404 114054 545004 149498
rect 544404 113818 544586 114054
rect 544822 113818 545004 114054
rect 544404 113734 545004 113818
rect 544404 113498 544586 113734
rect 544822 113498 545004 113734
rect 544404 78054 545004 113498
rect 544404 77818 544586 78054
rect 544822 77818 545004 78054
rect 544404 77734 545004 77818
rect 544404 77498 544586 77734
rect 544822 77498 545004 77734
rect 544404 42054 545004 77498
rect 544404 41818 544586 42054
rect 544822 41818 545004 42054
rect 544404 41734 545004 41818
rect 544404 41498 544586 41734
rect 544822 41498 545004 41734
rect 544404 6054 545004 41498
rect 544404 5818 544586 6054
rect 544822 5818 545004 6054
rect 544404 5734 545004 5818
rect 544404 5498 544586 5734
rect 544822 5498 545004 5734
rect 544404 -2186 545004 5498
rect 544404 -2422 544586 -2186
rect 544822 -2422 545004 -2186
rect 544404 -2506 545004 -2422
rect 544404 -2742 544586 -2506
rect 544822 -2742 545004 -2506
rect 544404 -3684 545004 -2742
rect 548004 693654 548604 707962
rect 548004 693418 548186 693654
rect 548422 693418 548604 693654
rect 548004 693334 548604 693418
rect 548004 693098 548186 693334
rect 548422 693098 548604 693334
rect 548004 657654 548604 693098
rect 548004 657418 548186 657654
rect 548422 657418 548604 657654
rect 548004 657334 548604 657418
rect 548004 657098 548186 657334
rect 548422 657098 548604 657334
rect 548004 621654 548604 657098
rect 548004 621418 548186 621654
rect 548422 621418 548604 621654
rect 548004 621334 548604 621418
rect 548004 621098 548186 621334
rect 548422 621098 548604 621334
rect 548004 585654 548604 621098
rect 548004 585418 548186 585654
rect 548422 585418 548604 585654
rect 548004 585334 548604 585418
rect 548004 585098 548186 585334
rect 548422 585098 548604 585334
rect 548004 549654 548604 585098
rect 548004 549418 548186 549654
rect 548422 549418 548604 549654
rect 548004 549334 548604 549418
rect 548004 549098 548186 549334
rect 548422 549098 548604 549334
rect 548004 513654 548604 549098
rect 548004 513418 548186 513654
rect 548422 513418 548604 513654
rect 548004 513334 548604 513418
rect 548004 513098 548186 513334
rect 548422 513098 548604 513334
rect 548004 477654 548604 513098
rect 548004 477418 548186 477654
rect 548422 477418 548604 477654
rect 548004 477334 548604 477418
rect 548004 477098 548186 477334
rect 548422 477098 548604 477334
rect 548004 441654 548604 477098
rect 548004 441418 548186 441654
rect 548422 441418 548604 441654
rect 548004 441334 548604 441418
rect 548004 441098 548186 441334
rect 548422 441098 548604 441334
rect 548004 405654 548604 441098
rect 548004 405418 548186 405654
rect 548422 405418 548604 405654
rect 548004 405334 548604 405418
rect 548004 405098 548186 405334
rect 548422 405098 548604 405334
rect 548004 369654 548604 405098
rect 548004 369418 548186 369654
rect 548422 369418 548604 369654
rect 548004 369334 548604 369418
rect 548004 369098 548186 369334
rect 548422 369098 548604 369334
rect 548004 333654 548604 369098
rect 548004 333418 548186 333654
rect 548422 333418 548604 333654
rect 548004 333334 548604 333418
rect 548004 333098 548186 333334
rect 548422 333098 548604 333334
rect 548004 297654 548604 333098
rect 548004 297418 548186 297654
rect 548422 297418 548604 297654
rect 548004 297334 548604 297418
rect 548004 297098 548186 297334
rect 548422 297098 548604 297334
rect 548004 261654 548604 297098
rect 548004 261418 548186 261654
rect 548422 261418 548604 261654
rect 548004 261334 548604 261418
rect 548004 261098 548186 261334
rect 548422 261098 548604 261334
rect 548004 225654 548604 261098
rect 548004 225418 548186 225654
rect 548422 225418 548604 225654
rect 548004 225334 548604 225418
rect 548004 225098 548186 225334
rect 548422 225098 548604 225334
rect 548004 189654 548604 225098
rect 548004 189418 548186 189654
rect 548422 189418 548604 189654
rect 548004 189334 548604 189418
rect 548004 189098 548186 189334
rect 548422 189098 548604 189334
rect 548004 153654 548604 189098
rect 548004 153418 548186 153654
rect 548422 153418 548604 153654
rect 548004 153334 548604 153418
rect 548004 153098 548186 153334
rect 548422 153098 548604 153334
rect 548004 117654 548604 153098
rect 548004 117418 548186 117654
rect 548422 117418 548604 117654
rect 548004 117334 548604 117418
rect 548004 117098 548186 117334
rect 548422 117098 548604 117334
rect 548004 81654 548604 117098
rect 548004 81418 548186 81654
rect 548422 81418 548604 81654
rect 548004 81334 548604 81418
rect 548004 81098 548186 81334
rect 548422 81098 548604 81334
rect 548004 45654 548604 81098
rect 548004 45418 548186 45654
rect 548422 45418 548604 45654
rect 548004 45334 548604 45418
rect 548004 45098 548186 45334
rect 548422 45098 548604 45334
rect 548004 9654 548604 45098
rect 548004 9418 548186 9654
rect 548422 9418 548604 9654
rect 548004 9334 548604 9418
rect 548004 9098 548186 9334
rect 548422 9098 548604 9334
rect 548004 -4026 548604 9098
rect 548004 -4262 548186 -4026
rect 548422 -4262 548604 -4026
rect 548004 -4346 548604 -4262
rect 548004 -4582 548186 -4346
rect 548422 -4582 548604 -4346
rect 548004 -5524 548604 -4582
rect 551604 697254 552204 709802
rect 569604 711278 570204 711300
rect 569604 711042 569786 711278
rect 570022 711042 570204 711278
rect 569604 710958 570204 711042
rect 569604 710722 569786 710958
rect 570022 710722 570204 710958
rect 566004 709438 566604 709460
rect 566004 709202 566186 709438
rect 566422 709202 566604 709438
rect 566004 709118 566604 709202
rect 566004 708882 566186 709118
rect 566422 708882 566604 709118
rect 562404 707598 563004 707620
rect 562404 707362 562586 707598
rect 562822 707362 563004 707598
rect 562404 707278 563004 707362
rect 562404 707042 562586 707278
rect 562822 707042 563004 707278
rect 551604 697018 551786 697254
rect 552022 697018 552204 697254
rect 551604 696934 552204 697018
rect 551604 696698 551786 696934
rect 552022 696698 552204 696934
rect 551604 661254 552204 696698
rect 551604 661018 551786 661254
rect 552022 661018 552204 661254
rect 551604 660934 552204 661018
rect 551604 660698 551786 660934
rect 552022 660698 552204 660934
rect 551604 625254 552204 660698
rect 551604 625018 551786 625254
rect 552022 625018 552204 625254
rect 551604 624934 552204 625018
rect 551604 624698 551786 624934
rect 552022 624698 552204 624934
rect 551604 589254 552204 624698
rect 551604 589018 551786 589254
rect 552022 589018 552204 589254
rect 551604 588934 552204 589018
rect 551604 588698 551786 588934
rect 552022 588698 552204 588934
rect 551604 553254 552204 588698
rect 551604 553018 551786 553254
rect 552022 553018 552204 553254
rect 551604 552934 552204 553018
rect 551604 552698 551786 552934
rect 552022 552698 552204 552934
rect 551604 517254 552204 552698
rect 551604 517018 551786 517254
rect 552022 517018 552204 517254
rect 551604 516934 552204 517018
rect 551604 516698 551786 516934
rect 552022 516698 552204 516934
rect 551604 481254 552204 516698
rect 551604 481018 551786 481254
rect 552022 481018 552204 481254
rect 551604 480934 552204 481018
rect 551604 480698 551786 480934
rect 552022 480698 552204 480934
rect 551604 445254 552204 480698
rect 551604 445018 551786 445254
rect 552022 445018 552204 445254
rect 551604 444934 552204 445018
rect 551604 444698 551786 444934
rect 552022 444698 552204 444934
rect 551604 409254 552204 444698
rect 551604 409018 551786 409254
rect 552022 409018 552204 409254
rect 551604 408934 552204 409018
rect 551604 408698 551786 408934
rect 552022 408698 552204 408934
rect 551604 373254 552204 408698
rect 551604 373018 551786 373254
rect 552022 373018 552204 373254
rect 551604 372934 552204 373018
rect 551604 372698 551786 372934
rect 552022 372698 552204 372934
rect 551604 337254 552204 372698
rect 551604 337018 551786 337254
rect 552022 337018 552204 337254
rect 551604 336934 552204 337018
rect 551604 336698 551786 336934
rect 552022 336698 552204 336934
rect 551604 301254 552204 336698
rect 551604 301018 551786 301254
rect 552022 301018 552204 301254
rect 551604 300934 552204 301018
rect 551604 300698 551786 300934
rect 552022 300698 552204 300934
rect 551604 265254 552204 300698
rect 551604 265018 551786 265254
rect 552022 265018 552204 265254
rect 551604 264934 552204 265018
rect 551604 264698 551786 264934
rect 552022 264698 552204 264934
rect 551604 229254 552204 264698
rect 551604 229018 551786 229254
rect 552022 229018 552204 229254
rect 551604 228934 552204 229018
rect 551604 228698 551786 228934
rect 552022 228698 552204 228934
rect 551604 193254 552204 228698
rect 551604 193018 551786 193254
rect 552022 193018 552204 193254
rect 551604 192934 552204 193018
rect 551604 192698 551786 192934
rect 552022 192698 552204 192934
rect 551604 157254 552204 192698
rect 551604 157018 551786 157254
rect 552022 157018 552204 157254
rect 551604 156934 552204 157018
rect 551604 156698 551786 156934
rect 552022 156698 552204 156934
rect 551604 121254 552204 156698
rect 551604 121018 551786 121254
rect 552022 121018 552204 121254
rect 551604 120934 552204 121018
rect 551604 120698 551786 120934
rect 552022 120698 552204 120934
rect 551604 85254 552204 120698
rect 551604 85018 551786 85254
rect 552022 85018 552204 85254
rect 551604 84934 552204 85018
rect 551604 84698 551786 84934
rect 552022 84698 552204 84934
rect 551604 49254 552204 84698
rect 551604 49018 551786 49254
rect 552022 49018 552204 49254
rect 551604 48934 552204 49018
rect 551604 48698 551786 48934
rect 552022 48698 552204 48934
rect 551604 13254 552204 48698
rect 551604 13018 551786 13254
rect 552022 13018 552204 13254
rect 551604 12934 552204 13018
rect 551604 12698 551786 12934
rect 552022 12698 552204 12934
rect 533604 -7022 533786 -6786
rect 534022 -7022 534204 -6786
rect 533604 -7106 534204 -7022
rect 533604 -7342 533786 -7106
rect 534022 -7342 534204 -7106
rect 533604 -7364 534204 -7342
rect 551604 -5866 552204 12698
rect 558804 705758 559404 705780
rect 558804 705522 558986 705758
rect 559222 705522 559404 705758
rect 558804 705438 559404 705522
rect 558804 705202 558986 705438
rect 559222 705202 559404 705438
rect 558804 668454 559404 705202
rect 558804 668218 558986 668454
rect 559222 668218 559404 668454
rect 558804 668134 559404 668218
rect 558804 667898 558986 668134
rect 559222 667898 559404 668134
rect 558804 632454 559404 667898
rect 558804 632218 558986 632454
rect 559222 632218 559404 632454
rect 558804 632134 559404 632218
rect 558804 631898 558986 632134
rect 559222 631898 559404 632134
rect 558804 596454 559404 631898
rect 558804 596218 558986 596454
rect 559222 596218 559404 596454
rect 558804 596134 559404 596218
rect 558804 595898 558986 596134
rect 559222 595898 559404 596134
rect 558804 560454 559404 595898
rect 558804 560218 558986 560454
rect 559222 560218 559404 560454
rect 558804 560134 559404 560218
rect 558804 559898 558986 560134
rect 559222 559898 559404 560134
rect 558804 524454 559404 559898
rect 558804 524218 558986 524454
rect 559222 524218 559404 524454
rect 558804 524134 559404 524218
rect 558804 523898 558986 524134
rect 559222 523898 559404 524134
rect 558804 488454 559404 523898
rect 558804 488218 558986 488454
rect 559222 488218 559404 488454
rect 558804 488134 559404 488218
rect 558804 487898 558986 488134
rect 559222 487898 559404 488134
rect 558804 452454 559404 487898
rect 558804 452218 558986 452454
rect 559222 452218 559404 452454
rect 558804 452134 559404 452218
rect 558804 451898 558986 452134
rect 559222 451898 559404 452134
rect 558804 416454 559404 451898
rect 558804 416218 558986 416454
rect 559222 416218 559404 416454
rect 558804 416134 559404 416218
rect 558804 415898 558986 416134
rect 559222 415898 559404 416134
rect 558804 380454 559404 415898
rect 558804 380218 558986 380454
rect 559222 380218 559404 380454
rect 558804 380134 559404 380218
rect 558804 379898 558986 380134
rect 559222 379898 559404 380134
rect 558804 344454 559404 379898
rect 558804 344218 558986 344454
rect 559222 344218 559404 344454
rect 558804 344134 559404 344218
rect 558804 343898 558986 344134
rect 559222 343898 559404 344134
rect 558804 308454 559404 343898
rect 558804 308218 558986 308454
rect 559222 308218 559404 308454
rect 558804 308134 559404 308218
rect 558804 307898 558986 308134
rect 559222 307898 559404 308134
rect 558804 272454 559404 307898
rect 558804 272218 558986 272454
rect 559222 272218 559404 272454
rect 558804 272134 559404 272218
rect 558804 271898 558986 272134
rect 559222 271898 559404 272134
rect 558804 236454 559404 271898
rect 558804 236218 558986 236454
rect 559222 236218 559404 236454
rect 558804 236134 559404 236218
rect 558804 235898 558986 236134
rect 559222 235898 559404 236134
rect 558804 200454 559404 235898
rect 558804 200218 558986 200454
rect 559222 200218 559404 200454
rect 558804 200134 559404 200218
rect 558804 199898 558986 200134
rect 559222 199898 559404 200134
rect 558804 164454 559404 199898
rect 558804 164218 558986 164454
rect 559222 164218 559404 164454
rect 558804 164134 559404 164218
rect 558804 163898 558986 164134
rect 559222 163898 559404 164134
rect 558804 128454 559404 163898
rect 558804 128218 558986 128454
rect 559222 128218 559404 128454
rect 558804 128134 559404 128218
rect 558804 127898 558986 128134
rect 559222 127898 559404 128134
rect 558804 92454 559404 127898
rect 558804 92218 558986 92454
rect 559222 92218 559404 92454
rect 558804 92134 559404 92218
rect 558804 91898 558986 92134
rect 559222 91898 559404 92134
rect 558804 56454 559404 91898
rect 558804 56218 558986 56454
rect 559222 56218 559404 56454
rect 558804 56134 559404 56218
rect 558804 55898 558986 56134
rect 559222 55898 559404 56134
rect 558804 20454 559404 55898
rect 558804 20218 558986 20454
rect 559222 20218 559404 20454
rect 558804 20134 559404 20218
rect 558804 19898 558986 20134
rect 559222 19898 559404 20134
rect 558804 -1266 559404 19898
rect 558804 -1502 558986 -1266
rect 559222 -1502 559404 -1266
rect 558804 -1586 559404 -1502
rect 558804 -1822 558986 -1586
rect 559222 -1822 559404 -1586
rect 558804 -1844 559404 -1822
rect 562404 672054 563004 707042
rect 562404 671818 562586 672054
rect 562822 671818 563004 672054
rect 562404 671734 563004 671818
rect 562404 671498 562586 671734
rect 562822 671498 563004 671734
rect 562404 636054 563004 671498
rect 562404 635818 562586 636054
rect 562822 635818 563004 636054
rect 562404 635734 563004 635818
rect 562404 635498 562586 635734
rect 562822 635498 563004 635734
rect 562404 600054 563004 635498
rect 562404 599818 562586 600054
rect 562822 599818 563004 600054
rect 562404 599734 563004 599818
rect 562404 599498 562586 599734
rect 562822 599498 563004 599734
rect 562404 564054 563004 599498
rect 562404 563818 562586 564054
rect 562822 563818 563004 564054
rect 562404 563734 563004 563818
rect 562404 563498 562586 563734
rect 562822 563498 563004 563734
rect 562404 528054 563004 563498
rect 562404 527818 562586 528054
rect 562822 527818 563004 528054
rect 562404 527734 563004 527818
rect 562404 527498 562586 527734
rect 562822 527498 563004 527734
rect 562404 492054 563004 527498
rect 562404 491818 562586 492054
rect 562822 491818 563004 492054
rect 562404 491734 563004 491818
rect 562404 491498 562586 491734
rect 562822 491498 563004 491734
rect 562404 456054 563004 491498
rect 562404 455818 562586 456054
rect 562822 455818 563004 456054
rect 562404 455734 563004 455818
rect 562404 455498 562586 455734
rect 562822 455498 563004 455734
rect 562404 420054 563004 455498
rect 562404 419818 562586 420054
rect 562822 419818 563004 420054
rect 562404 419734 563004 419818
rect 562404 419498 562586 419734
rect 562822 419498 563004 419734
rect 562404 384054 563004 419498
rect 562404 383818 562586 384054
rect 562822 383818 563004 384054
rect 562404 383734 563004 383818
rect 562404 383498 562586 383734
rect 562822 383498 563004 383734
rect 562404 348054 563004 383498
rect 562404 347818 562586 348054
rect 562822 347818 563004 348054
rect 562404 347734 563004 347818
rect 562404 347498 562586 347734
rect 562822 347498 563004 347734
rect 562404 312054 563004 347498
rect 562404 311818 562586 312054
rect 562822 311818 563004 312054
rect 562404 311734 563004 311818
rect 562404 311498 562586 311734
rect 562822 311498 563004 311734
rect 562404 276054 563004 311498
rect 562404 275818 562586 276054
rect 562822 275818 563004 276054
rect 562404 275734 563004 275818
rect 562404 275498 562586 275734
rect 562822 275498 563004 275734
rect 562404 240054 563004 275498
rect 562404 239818 562586 240054
rect 562822 239818 563004 240054
rect 562404 239734 563004 239818
rect 562404 239498 562586 239734
rect 562822 239498 563004 239734
rect 562404 204054 563004 239498
rect 562404 203818 562586 204054
rect 562822 203818 563004 204054
rect 562404 203734 563004 203818
rect 562404 203498 562586 203734
rect 562822 203498 563004 203734
rect 562404 168054 563004 203498
rect 562404 167818 562586 168054
rect 562822 167818 563004 168054
rect 562404 167734 563004 167818
rect 562404 167498 562586 167734
rect 562822 167498 563004 167734
rect 562404 132054 563004 167498
rect 562404 131818 562586 132054
rect 562822 131818 563004 132054
rect 562404 131734 563004 131818
rect 562404 131498 562586 131734
rect 562822 131498 563004 131734
rect 562404 96054 563004 131498
rect 562404 95818 562586 96054
rect 562822 95818 563004 96054
rect 562404 95734 563004 95818
rect 562404 95498 562586 95734
rect 562822 95498 563004 95734
rect 562404 60054 563004 95498
rect 562404 59818 562586 60054
rect 562822 59818 563004 60054
rect 562404 59734 563004 59818
rect 562404 59498 562586 59734
rect 562822 59498 563004 59734
rect 562404 24054 563004 59498
rect 562404 23818 562586 24054
rect 562822 23818 563004 24054
rect 562404 23734 563004 23818
rect 562404 23498 562586 23734
rect 562822 23498 563004 23734
rect 562404 -3106 563004 23498
rect 562404 -3342 562586 -3106
rect 562822 -3342 563004 -3106
rect 562404 -3426 563004 -3342
rect 562404 -3662 562586 -3426
rect 562822 -3662 563004 -3426
rect 562404 -3684 563004 -3662
rect 566004 675654 566604 708882
rect 566004 675418 566186 675654
rect 566422 675418 566604 675654
rect 566004 675334 566604 675418
rect 566004 675098 566186 675334
rect 566422 675098 566604 675334
rect 566004 639654 566604 675098
rect 566004 639418 566186 639654
rect 566422 639418 566604 639654
rect 566004 639334 566604 639418
rect 566004 639098 566186 639334
rect 566422 639098 566604 639334
rect 566004 603654 566604 639098
rect 566004 603418 566186 603654
rect 566422 603418 566604 603654
rect 566004 603334 566604 603418
rect 566004 603098 566186 603334
rect 566422 603098 566604 603334
rect 566004 567654 566604 603098
rect 566004 567418 566186 567654
rect 566422 567418 566604 567654
rect 566004 567334 566604 567418
rect 566004 567098 566186 567334
rect 566422 567098 566604 567334
rect 566004 531654 566604 567098
rect 566004 531418 566186 531654
rect 566422 531418 566604 531654
rect 566004 531334 566604 531418
rect 566004 531098 566186 531334
rect 566422 531098 566604 531334
rect 566004 495654 566604 531098
rect 566004 495418 566186 495654
rect 566422 495418 566604 495654
rect 566004 495334 566604 495418
rect 566004 495098 566186 495334
rect 566422 495098 566604 495334
rect 566004 459654 566604 495098
rect 566004 459418 566186 459654
rect 566422 459418 566604 459654
rect 566004 459334 566604 459418
rect 566004 459098 566186 459334
rect 566422 459098 566604 459334
rect 566004 423654 566604 459098
rect 566004 423418 566186 423654
rect 566422 423418 566604 423654
rect 566004 423334 566604 423418
rect 566004 423098 566186 423334
rect 566422 423098 566604 423334
rect 566004 387654 566604 423098
rect 566004 387418 566186 387654
rect 566422 387418 566604 387654
rect 566004 387334 566604 387418
rect 566004 387098 566186 387334
rect 566422 387098 566604 387334
rect 566004 351654 566604 387098
rect 566004 351418 566186 351654
rect 566422 351418 566604 351654
rect 566004 351334 566604 351418
rect 566004 351098 566186 351334
rect 566422 351098 566604 351334
rect 566004 315654 566604 351098
rect 566004 315418 566186 315654
rect 566422 315418 566604 315654
rect 566004 315334 566604 315418
rect 566004 315098 566186 315334
rect 566422 315098 566604 315334
rect 566004 279654 566604 315098
rect 566004 279418 566186 279654
rect 566422 279418 566604 279654
rect 566004 279334 566604 279418
rect 566004 279098 566186 279334
rect 566422 279098 566604 279334
rect 566004 243654 566604 279098
rect 566004 243418 566186 243654
rect 566422 243418 566604 243654
rect 566004 243334 566604 243418
rect 566004 243098 566186 243334
rect 566422 243098 566604 243334
rect 566004 207654 566604 243098
rect 566004 207418 566186 207654
rect 566422 207418 566604 207654
rect 566004 207334 566604 207418
rect 566004 207098 566186 207334
rect 566422 207098 566604 207334
rect 566004 171654 566604 207098
rect 566004 171418 566186 171654
rect 566422 171418 566604 171654
rect 566004 171334 566604 171418
rect 566004 171098 566186 171334
rect 566422 171098 566604 171334
rect 566004 135654 566604 171098
rect 566004 135418 566186 135654
rect 566422 135418 566604 135654
rect 566004 135334 566604 135418
rect 566004 135098 566186 135334
rect 566422 135098 566604 135334
rect 566004 99654 566604 135098
rect 566004 99418 566186 99654
rect 566422 99418 566604 99654
rect 566004 99334 566604 99418
rect 566004 99098 566186 99334
rect 566422 99098 566604 99334
rect 566004 63654 566604 99098
rect 566004 63418 566186 63654
rect 566422 63418 566604 63654
rect 566004 63334 566604 63418
rect 566004 63098 566186 63334
rect 566422 63098 566604 63334
rect 566004 27654 566604 63098
rect 566004 27418 566186 27654
rect 566422 27418 566604 27654
rect 566004 27334 566604 27418
rect 566004 27098 566186 27334
rect 566422 27098 566604 27334
rect 566004 -4946 566604 27098
rect 566004 -5182 566186 -4946
rect 566422 -5182 566604 -4946
rect 566004 -5266 566604 -5182
rect 566004 -5502 566186 -5266
rect 566422 -5502 566604 -5266
rect 566004 -5524 566604 -5502
rect 569604 679254 570204 710722
rect 591760 711278 592360 711300
rect 591760 711042 591942 711278
rect 592178 711042 592360 711278
rect 591760 710958 592360 711042
rect 591760 710722 591942 710958
rect 592178 710722 592360 710958
rect 590840 710358 591440 710380
rect 590840 710122 591022 710358
rect 591258 710122 591440 710358
rect 590840 710038 591440 710122
rect 590840 709802 591022 710038
rect 591258 709802 591440 710038
rect 589920 709438 590520 709460
rect 589920 709202 590102 709438
rect 590338 709202 590520 709438
rect 589920 709118 590520 709202
rect 589920 708882 590102 709118
rect 590338 708882 590520 709118
rect 589000 708518 589600 708540
rect 589000 708282 589182 708518
rect 589418 708282 589600 708518
rect 589000 708198 589600 708282
rect 589000 707962 589182 708198
rect 589418 707962 589600 708198
rect 580404 706678 581004 707620
rect 588080 707598 588680 707620
rect 588080 707362 588262 707598
rect 588498 707362 588680 707598
rect 588080 707278 588680 707362
rect 588080 707042 588262 707278
rect 588498 707042 588680 707278
rect 580404 706442 580586 706678
rect 580822 706442 581004 706678
rect 580404 706358 581004 706442
rect 580404 706122 580586 706358
rect 580822 706122 581004 706358
rect 569604 679018 569786 679254
rect 570022 679018 570204 679254
rect 569604 678934 570204 679018
rect 569604 678698 569786 678934
rect 570022 678698 570204 678934
rect 569604 643254 570204 678698
rect 569604 643018 569786 643254
rect 570022 643018 570204 643254
rect 569604 642934 570204 643018
rect 569604 642698 569786 642934
rect 570022 642698 570204 642934
rect 569604 607254 570204 642698
rect 569604 607018 569786 607254
rect 570022 607018 570204 607254
rect 569604 606934 570204 607018
rect 569604 606698 569786 606934
rect 570022 606698 570204 606934
rect 569604 571254 570204 606698
rect 569604 571018 569786 571254
rect 570022 571018 570204 571254
rect 569604 570934 570204 571018
rect 569604 570698 569786 570934
rect 570022 570698 570204 570934
rect 569604 535254 570204 570698
rect 569604 535018 569786 535254
rect 570022 535018 570204 535254
rect 569604 534934 570204 535018
rect 569604 534698 569786 534934
rect 570022 534698 570204 534934
rect 569604 499254 570204 534698
rect 569604 499018 569786 499254
rect 570022 499018 570204 499254
rect 569604 498934 570204 499018
rect 569604 498698 569786 498934
rect 570022 498698 570204 498934
rect 569604 463254 570204 498698
rect 569604 463018 569786 463254
rect 570022 463018 570204 463254
rect 569604 462934 570204 463018
rect 569604 462698 569786 462934
rect 570022 462698 570204 462934
rect 569604 427254 570204 462698
rect 569604 427018 569786 427254
rect 570022 427018 570204 427254
rect 569604 426934 570204 427018
rect 569604 426698 569786 426934
rect 570022 426698 570204 426934
rect 569604 391254 570204 426698
rect 569604 391018 569786 391254
rect 570022 391018 570204 391254
rect 569604 390934 570204 391018
rect 569604 390698 569786 390934
rect 570022 390698 570204 390934
rect 569604 355254 570204 390698
rect 569604 355018 569786 355254
rect 570022 355018 570204 355254
rect 569604 354934 570204 355018
rect 569604 354698 569786 354934
rect 570022 354698 570204 354934
rect 569604 319254 570204 354698
rect 569604 319018 569786 319254
rect 570022 319018 570204 319254
rect 569604 318934 570204 319018
rect 569604 318698 569786 318934
rect 570022 318698 570204 318934
rect 569604 283254 570204 318698
rect 569604 283018 569786 283254
rect 570022 283018 570204 283254
rect 569604 282934 570204 283018
rect 569604 282698 569786 282934
rect 570022 282698 570204 282934
rect 569604 247254 570204 282698
rect 569604 247018 569786 247254
rect 570022 247018 570204 247254
rect 569604 246934 570204 247018
rect 569604 246698 569786 246934
rect 570022 246698 570204 246934
rect 569604 211254 570204 246698
rect 569604 211018 569786 211254
rect 570022 211018 570204 211254
rect 569604 210934 570204 211018
rect 569604 210698 569786 210934
rect 570022 210698 570204 210934
rect 569604 175254 570204 210698
rect 569604 175018 569786 175254
rect 570022 175018 570204 175254
rect 569604 174934 570204 175018
rect 569604 174698 569786 174934
rect 570022 174698 570204 174934
rect 569604 139254 570204 174698
rect 569604 139018 569786 139254
rect 570022 139018 570204 139254
rect 569604 138934 570204 139018
rect 569604 138698 569786 138934
rect 570022 138698 570204 138934
rect 569604 103254 570204 138698
rect 569604 103018 569786 103254
rect 570022 103018 570204 103254
rect 569604 102934 570204 103018
rect 569604 102698 569786 102934
rect 570022 102698 570204 102934
rect 569604 67254 570204 102698
rect 569604 67018 569786 67254
rect 570022 67018 570204 67254
rect 569604 66934 570204 67018
rect 569604 66698 569786 66934
rect 570022 66698 570204 66934
rect 569604 31254 570204 66698
rect 569604 31018 569786 31254
rect 570022 31018 570204 31254
rect 569604 30934 570204 31018
rect 569604 30698 569786 30934
rect 570022 30698 570204 30934
rect 551604 -6102 551786 -5866
rect 552022 -6102 552204 -5866
rect 551604 -6186 552204 -6102
rect 551604 -6422 551786 -6186
rect 552022 -6422 552204 -6186
rect 551604 -7364 552204 -6422
rect 569604 -6786 570204 30698
rect 576804 704838 577404 705780
rect 576804 704602 576986 704838
rect 577222 704602 577404 704838
rect 576804 704518 577404 704602
rect 576804 704282 576986 704518
rect 577222 704282 577404 704518
rect 576804 686454 577404 704282
rect 576804 686218 576986 686454
rect 577222 686218 577404 686454
rect 576804 686134 577404 686218
rect 576804 685898 576986 686134
rect 577222 685898 577404 686134
rect 576804 650454 577404 685898
rect 576804 650218 576986 650454
rect 577222 650218 577404 650454
rect 576804 650134 577404 650218
rect 576804 649898 576986 650134
rect 577222 649898 577404 650134
rect 576804 614454 577404 649898
rect 576804 614218 576986 614454
rect 577222 614218 577404 614454
rect 576804 614134 577404 614218
rect 576804 613898 576986 614134
rect 577222 613898 577404 614134
rect 576804 578454 577404 613898
rect 576804 578218 576986 578454
rect 577222 578218 577404 578454
rect 576804 578134 577404 578218
rect 576804 577898 576986 578134
rect 577222 577898 577404 578134
rect 576804 542454 577404 577898
rect 576804 542218 576986 542454
rect 577222 542218 577404 542454
rect 576804 542134 577404 542218
rect 576804 541898 576986 542134
rect 577222 541898 577404 542134
rect 576804 506454 577404 541898
rect 576804 506218 576986 506454
rect 577222 506218 577404 506454
rect 576804 506134 577404 506218
rect 576804 505898 576986 506134
rect 577222 505898 577404 506134
rect 576804 470454 577404 505898
rect 576804 470218 576986 470454
rect 577222 470218 577404 470454
rect 576804 470134 577404 470218
rect 576804 469898 576986 470134
rect 577222 469898 577404 470134
rect 576804 434454 577404 469898
rect 576804 434218 576986 434454
rect 577222 434218 577404 434454
rect 576804 434134 577404 434218
rect 576804 433898 576986 434134
rect 577222 433898 577404 434134
rect 576804 398454 577404 433898
rect 576804 398218 576986 398454
rect 577222 398218 577404 398454
rect 576804 398134 577404 398218
rect 576804 397898 576986 398134
rect 577222 397898 577404 398134
rect 576804 362454 577404 397898
rect 576804 362218 576986 362454
rect 577222 362218 577404 362454
rect 576804 362134 577404 362218
rect 576804 361898 576986 362134
rect 577222 361898 577404 362134
rect 576804 326454 577404 361898
rect 576804 326218 576986 326454
rect 577222 326218 577404 326454
rect 576804 326134 577404 326218
rect 576804 325898 576986 326134
rect 577222 325898 577404 326134
rect 576804 290454 577404 325898
rect 576804 290218 576986 290454
rect 577222 290218 577404 290454
rect 576804 290134 577404 290218
rect 576804 289898 576986 290134
rect 577222 289898 577404 290134
rect 576804 254454 577404 289898
rect 576804 254218 576986 254454
rect 577222 254218 577404 254454
rect 576804 254134 577404 254218
rect 576804 253898 576986 254134
rect 577222 253898 577404 254134
rect 576804 218454 577404 253898
rect 576804 218218 576986 218454
rect 577222 218218 577404 218454
rect 576804 218134 577404 218218
rect 576804 217898 576986 218134
rect 577222 217898 577404 218134
rect 576804 182454 577404 217898
rect 576804 182218 576986 182454
rect 577222 182218 577404 182454
rect 576804 182134 577404 182218
rect 576804 181898 576986 182134
rect 577222 181898 577404 182134
rect 576804 146454 577404 181898
rect 576804 146218 576986 146454
rect 577222 146218 577404 146454
rect 576804 146134 577404 146218
rect 576804 145898 576986 146134
rect 577222 145898 577404 146134
rect 576804 110454 577404 145898
rect 576804 110218 576986 110454
rect 577222 110218 577404 110454
rect 576804 110134 577404 110218
rect 576804 109898 576986 110134
rect 577222 109898 577404 110134
rect 576804 74454 577404 109898
rect 576804 74218 576986 74454
rect 577222 74218 577404 74454
rect 576804 74134 577404 74218
rect 576804 73898 576986 74134
rect 577222 73898 577404 74134
rect 576804 38454 577404 73898
rect 576804 38218 576986 38454
rect 577222 38218 577404 38454
rect 576804 38134 577404 38218
rect 576804 37898 576986 38134
rect 577222 37898 577404 38134
rect 576804 2454 577404 37898
rect 576804 2218 576986 2454
rect 577222 2218 577404 2454
rect 576804 2134 577404 2218
rect 576804 1898 576986 2134
rect 577222 1898 577404 2134
rect 576804 -346 577404 1898
rect 576804 -582 576986 -346
rect 577222 -582 577404 -346
rect 576804 -666 577404 -582
rect 576804 -902 576986 -666
rect 577222 -902 577404 -666
rect 576804 -1844 577404 -902
rect 580404 690054 581004 706122
rect 587160 706678 587760 706700
rect 587160 706442 587342 706678
rect 587578 706442 587760 706678
rect 587160 706358 587760 706442
rect 587160 706122 587342 706358
rect 587578 706122 587760 706358
rect 586240 705758 586840 705780
rect 586240 705522 586422 705758
rect 586658 705522 586840 705758
rect 586240 705438 586840 705522
rect 586240 705202 586422 705438
rect 586658 705202 586840 705438
rect 580404 689818 580586 690054
rect 580822 689818 581004 690054
rect 580404 689734 581004 689818
rect 580404 689498 580586 689734
rect 580822 689498 581004 689734
rect 580404 654054 581004 689498
rect 580404 653818 580586 654054
rect 580822 653818 581004 654054
rect 580404 653734 581004 653818
rect 580404 653498 580586 653734
rect 580822 653498 581004 653734
rect 580404 618054 581004 653498
rect 580404 617818 580586 618054
rect 580822 617818 581004 618054
rect 580404 617734 581004 617818
rect 580404 617498 580586 617734
rect 580822 617498 581004 617734
rect 580404 582054 581004 617498
rect 580404 581818 580586 582054
rect 580822 581818 581004 582054
rect 580404 581734 581004 581818
rect 580404 581498 580586 581734
rect 580822 581498 581004 581734
rect 580404 546054 581004 581498
rect 580404 545818 580586 546054
rect 580822 545818 581004 546054
rect 580404 545734 581004 545818
rect 580404 545498 580586 545734
rect 580822 545498 581004 545734
rect 580404 510054 581004 545498
rect 580404 509818 580586 510054
rect 580822 509818 581004 510054
rect 580404 509734 581004 509818
rect 580404 509498 580586 509734
rect 580822 509498 581004 509734
rect 580404 474054 581004 509498
rect 580404 473818 580586 474054
rect 580822 473818 581004 474054
rect 580404 473734 581004 473818
rect 580404 473498 580586 473734
rect 580822 473498 581004 473734
rect 580404 438054 581004 473498
rect 580404 437818 580586 438054
rect 580822 437818 581004 438054
rect 580404 437734 581004 437818
rect 580404 437498 580586 437734
rect 580822 437498 581004 437734
rect 580404 402054 581004 437498
rect 580404 401818 580586 402054
rect 580822 401818 581004 402054
rect 580404 401734 581004 401818
rect 580404 401498 580586 401734
rect 580822 401498 581004 401734
rect 580404 366054 581004 401498
rect 580404 365818 580586 366054
rect 580822 365818 581004 366054
rect 580404 365734 581004 365818
rect 580404 365498 580586 365734
rect 580822 365498 581004 365734
rect 580404 330054 581004 365498
rect 580404 329818 580586 330054
rect 580822 329818 581004 330054
rect 580404 329734 581004 329818
rect 580404 329498 580586 329734
rect 580822 329498 581004 329734
rect 580404 294054 581004 329498
rect 580404 293818 580586 294054
rect 580822 293818 581004 294054
rect 580404 293734 581004 293818
rect 580404 293498 580586 293734
rect 580822 293498 581004 293734
rect 580404 258054 581004 293498
rect 580404 257818 580586 258054
rect 580822 257818 581004 258054
rect 580404 257734 581004 257818
rect 580404 257498 580586 257734
rect 580822 257498 581004 257734
rect 580404 222054 581004 257498
rect 580404 221818 580586 222054
rect 580822 221818 581004 222054
rect 580404 221734 581004 221818
rect 580404 221498 580586 221734
rect 580822 221498 581004 221734
rect 580404 186054 581004 221498
rect 580404 185818 580586 186054
rect 580822 185818 581004 186054
rect 580404 185734 581004 185818
rect 580404 185498 580586 185734
rect 580822 185498 581004 185734
rect 580404 150054 581004 185498
rect 580404 149818 580586 150054
rect 580822 149818 581004 150054
rect 580404 149734 581004 149818
rect 580404 149498 580586 149734
rect 580822 149498 581004 149734
rect 580404 114054 581004 149498
rect 580404 113818 580586 114054
rect 580822 113818 581004 114054
rect 580404 113734 581004 113818
rect 580404 113498 580586 113734
rect 580822 113498 581004 113734
rect 580404 78054 581004 113498
rect 580404 77818 580586 78054
rect 580822 77818 581004 78054
rect 580404 77734 581004 77818
rect 580404 77498 580586 77734
rect 580822 77498 581004 77734
rect 580404 42054 581004 77498
rect 580404 41818 580586 42054
rect 580822 41818 581004 42054
rect 580404 41734 581004 41818
rect 580404 41498 580586 41734
rect 580822 41498 581004 41734
rect 580404 6054 581004 41498
rect 580404 5818 580586 6054
rect 580822 5818 581004 6054
rect 580404 5734 581004 5818
rect 580404 5498 580586 5734
rect 580822 5498 581004 5734
rect 580404 -2186 581004 5498
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 686454 585920 704282
rect 585320 686218 585502 686454
rect 585738 686218 585920 686454
rect 585320 686134 585920 686218
rect 585320 685898 585502 686134
rect 585738 685898 585920 686134
rect 585320 650454 585920 685898
rect 585320 650218 585502 650454
rect 585738 650218 585920 650454
rect 585320 650134 585920 650218
rect 585320 649898 585502 650134
rect 585738 649898 585920 650134
rect 585320 614454 585920 649898
rect 585320 614218 585502 614454
rect 585738 614218 585920 614454
rect 585320 614134 585920 614218
rect 585320 613898 585502 614134
rect 585738 613898 585920 614134
rect 585320 578454 585920 613898
rect 585320 578218 585502 578454
rect 585738 578218 585920 578454
rect 585320 578134 585920 578218
rect 585320 577898 585502 578134
rect 585738 577898 585920 578134
rect 585320 542454 585920 577898
rect 585320 542218 585502 542454
rect 585738 542218 585920 542454
rect 585320 542134 585920 542218
rect 585320 541898 585502 542134
rect 585738 541898 585920 542134
rect 585320 506454 585920 541898
rect 585320 506218 585502 506454
rect 585738 506218 585920 506454
rect 585320 506134 585920 506218
rect 585320 505898 585502 506134
rect 585738 505898 585920 506134
rect 585320 470454 585920 505898
rect 585320 470218 585502 470454
rect 585738 470218 585920 470454
rect 585320 470134 585920 470218
rect 585320 469898 585502 470134
rect 585738 469898 585920 470134
rect 585320 434454 585920 469898
rect 585320 434218 585502 434454
rect 585738 434218 585920 434454
rect 585320 434134 585920 434218
rect 585320 433898 585502 434134
rect 585738 433898 585920 434134
rect 585320 398454 585920 433898
rect 585320 398218 585502 398454
rect 585738 398218 585920 398454
rect 585320 398134 585920 398218
rect 585320 397898 585502 398134
rect 585738 397898 585920 398134
rect 585320 362454 585920 397898
rect 585320 362218 585502 362454
rect 585738 362218 585920 362454
rect 585320 362134 585920 362218
rect 585320 361898 585502 362134
rect 585738 361898 585920 362134
rect 585320 326454 585920 361898
rect 585320 326218 585502 326454
rect 585738 326218 585920 326454
rect 585320 326134 585920 326218
rect 585320 325898 585502 326134
rect 585738 325898 585920 326134
rect 585320 290454 585920 325898
rect 585320 290218 585502 290454
rect 585738 290218 585920 290454
rect 585320 290134 585920 290218
rect 585320 289898 585502 290134
rect 585738 289898 585920 290134
rect 585320 254454 585920 289898
rect 585320 254218 585502 254454
rect 585738 254218 585920 254454
rect 585320 254134 585920 254218
rect 585320 253898 585502 254134
rect 585738 253898 585920 254134
rect 585320 218454 585920 253898
rect 585320 218218 585502 218454
rect 585738 218218 585920 218454
rect 585320 218134 585920 218218
rect 585320 217898 585502 218134
rect 585738 217898 585920 218134
rect 585320 182454 585920 217898
rect 585320 182218 585502 182454
rect 585738 182218 585920 182454
rect 585320 182134 585920 182218
rect 585320 181898 585502 182134
rect 585738 181898 585920 182134
rect 585320 146454 585920 181898
rect 585320 146218 585502 146454
rect 585738 146218 585920 146454
rect 585320 146134 585920 146218
rect 585320 145898 585502 146134
rect 585738 145898 585920 146134
rect 585320 110454 585920 145898
rect 585320 110218 585502 110454
rect 585738 110218 585920 110454
rect 585320 110134 585920 110218
rect 585320 109898 585502 110134
rect 585738 109898 585920 110134
rect 585320 74454 585920 109898
rect 585320 74218 585502 74454
rect 585738 74218 585920 74454
rect 585320 74134 585920 74218
rect 585320 73898 585502 74134
rect 585738 73898 585920 74134
rect 585320 38454 585920 73898
rect 585320 38218 585502 38454
rect 585738 38218 585920 38454
rect 585320 38134 585920 38218
rect 585320 37898 585502 38134
rect 585738 37898 585920 38134
rect 585320 2454 585920 37898
rect 585320 2218 585502 2454
rect 585738 2218 585920 2454
rect 585320 2134 585920 2218
rect 585320 1898 585502 2134
rect 585738 1898 585920 2134
rect 585320 -346 585920 1898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586240 668454 586840 705202
rect 586240 668218 586422 668454
rect 586658 668218 586840 668454
rect 586240 668134 586840 668218
rect 586240 667898 586422 668134
rect 586658 667898 586840 668134
rect 586240 632454 586840 667898
rect 586240 632218 586422 632454
rect 586658 632218 586840 632454
rect 586240 632134 586840 632218
rect 586240 631898 586422 632134
rect 586658 631898 586840 632134
rect 586240 596454 586840 631898
rect 586240 596218 586422 596454
rect 586658 596218 586840 596454
rect 586240 596134 586840 596218
rect 586240 595898 586422 596134
rect 586658 595898 586840 596134
rect 586240 560454 586840 595898
rect 586240 560218 586422 560454
rect 586658 560218 586840 560454
rect 586240 560134 586840 560218
rect 586240 559898 586422 560134
rect 586658 559898 586840 560134
rect 586240 524454 586840 559898
rect 586240 524218 586422 524454
rect 586658 524218 586840 524454
rect 586240 524134 586840 524218
rect 586240 523898 586422 524134
rect 586658 523898 586840 524134
rect 586240 488454 586840 523898
rect 586240 488218 586422 488454
rect 586658 488218 586840 488454
rect 586240 488134 586840 488218
rect 586240 487898 586422 488134
rect 586658 487898 586840 488134
rect 586240 452454 586840 487898
rect 586240 452218 586422 452454
rect 586658 452218 586840 452454
rect 586240 452134 586840 452218
rect 586240 451898 586422 452134
rect 586658 451898 586840 452134
rect 586240 416454 586840 451898
rect 586240 416218 586422 416454
rect 586658 416218 586840 416454
rect 586240 416134 586840 416218
rect 586240 415898 586422 416134
rect 586658 415898 586840 416134
rect 586240 380454 586840 415898
rect 586240 380218 586422 380454
rect 586658 380218 586840 380454
rect 586240 380134 586840 380218
rect 586240 379898 586422 380134
rect 586658 379898 586840 380134
rect 586240 344454 586840 379898
rect 586240 344218 586422 344454
rect 586658 344218 586840 344454
rect 586240 344134 586840 344218
rect 586240 343898 586422 344134
rect 586658 343898 586840 344134
rect 586240 308454 586840 343898
rect 586240 308218 586422 308454
rect 586658 308218 586840 308454
rect 586240 308134 586840 308218
rect 586240 307898 586422 308134
rect 586658 307898 586840 308134
rect 586240 272454 586840 307898
rect 586240 272218 586422 272454
rect 586658 272218 586840 272454
rect 586240 272134 586840 272218
rect 586240 271898 586422 272134
rect 586658 271898 586840 272134
rect 586240 236454 586840 271898
rect 586240 236218 586422 236454
rect 586658 236218 586840 236454
rect 586240 236134 586840 236218
rect 586240 235898 586422 236134
rect 586658 235898 586840 236134
rect 586240 200454 586840 235898
rect 586240 200218 586422 200454
rect 586658 200218 586840 200454
rect 586240 200134 586840 200218
rect 586240 199898 586422 200134
rect 586658 199898 586840 200134
rect 586240 164454 586840 199898
rect 586240 164218 586422 164454
rect 586658 164218 586840 164454
rect 586240 164134 586840 164218
rect 586240 163898 586422 164134
rect 586658 163898 586840 164134
rect 586240 128454 586840 163898
rect 586240 128218 586422 128454
rect 586658 128218 586840 128454
rect 586240 128134 586840 128218
rect 586240 127898 586422 128134
rect 586658 127898 586840 128134
rect 586240 92454 586840 127898
rect 586240 92218 586422 92454
rect 586658 92218 586840 92454
rect 586240 92134 586840 92218
rect 586240 91898 586422 92134
rect 586658 91898 586840 92134
rect 586240 56454 586840 91898
rect 586240 56218 586422 56454
rect 586658 56218 586840 56454
rect 586240 56134 586840 56218
rect 586240 55898 586422 56134
rect 586658 55898 586840 56134
rect 586240 20454 586840 55898
rect 586240 20218 586422 20454
rect 586658 20218 586840 20454
rect 586240 20134 586840 20218
rect 586240 19898 586422 20134
rect 586658 19898 586840 20134
rect 586240 -1266 586840 19898
rect 586240 -1502 586422 -1266
rect 586658 -1502 586840 -1266
rect 586240 -1586 586840 -1502
rect 586240 -1822 586422 -1586
rect 586658 -1822 586840 -1586
rect 586240 -1844 586840 -1822
rect 587160 690054 587760 706122
rect 587160 689818 587342 690054
rect 587578 689818 587760 690054
rect 587160 689734 587760 689818
rect 587160 689498 587342 689734
rect 587578 689498 587760 689734
rect 587160 654054 587760 689498
rect 587160 653818 587342 654054
rect 587578 653818 587760 654054
rect 587160 653734 587760 653818
rect 587160 653498 587342 653734
rect 587578 653498 587760 653734
rect 587160 618054 587760 653498
rect 587160 617818 587342 618054
rect 587578 617818 587760 618054
rect 587160 617734 587760 617818
rect 587160 617498 587342 617734
rect 587578 617498 587760 617734
rect 587160 582054 587760 617498
rect 587160 581818 587342 582054
rect 587578 581818 587760 582054
rect 587160 581734 587760 581818
rect 587160 581498 587342 581734
rect 587578 581498 587760 581734
rect 587160 546054 587760 581498
rect 587160 545818 587342 546054
rect 587578 545818 587760 546054
rect 587160 545734 587760 545818
rect 587160 545498 587342 545734
rect 587578 545498 587760 545734
rect 587160 510054 587760 545498
rect 587160 509818 587342 510054
rect 587578 509818 587760 510054
rect 587160 509734 587760 509818
rect 587160 509498 587342 509734
rect 587578 509498 587760 509734
rect 587160 474054 587760 509498
rect 587160 473818 587342 474054
rect 587578 473818 587760 474054
rect 587160 473734 587760 473818
rect 587160 473498 587342 473734
rect 587578 473498 587760 473734
rect 587160 438054 587760 473498
rect 587160 437818 587342 438054
rect 587578 437818 587760 438054
rect 587160 437734 587760 437818
rect 587160 437498 587342 437734
rect 587578 437498 587760 437734
rect 587160 402054 587760 437498
rect 587160 401818 587342 402054
rect 587578 401818 587760 402054
rect 587160 401734 587760 401818
rect 587160 401498 587342 401734
rect 587578 401498 587760 401734
rect 587160 366054 587760 401498
rect 587160 365818 587342 366054
rect 587578 365818 587760 366054
rect 587160 365734 587760 365818
rect 587160 365498 587342 365734
rect 587578 365498 587760 365734
rect 587160 330054 587760 365498
rect 587160 329818 587342 330054
rect 587578 329818 587760 330054
rect 587160 329734 587760 329818
rect 587160 329498 587342 329734
rect 587578 329498 587760 329734
rect 587160 294054 587760 329498
rect 587160 293818 587342 294054
rect 587578 293818 587760 294054
rect 587160 293734 587760 293818
rect 587160 293498 587342 293734
rect 587578 293498 587760 293734
rect 587160 258054 587760 293498
rect 587160 257818 587342 258054
rect 587578 257818 587760 258054
rect 587160 257734 587760 257818
rect 587160 257498 587342 257734
rect 587578 257498 587760 257734
rect 587160 222054 587760 257498
rect 587160 221818 587342 222054
rect 587578 221818 587760 222054
rect 587160 221734 587760 221818
rect 587160 221498 587342 221734
rect 587578 221498 587760 221734
rect 587160 186054 587760 221498
rect 587160 185818 587342 186054
rect 587578 185818 587760 186054
rect 587160 185734 587760 185818
rect 587160 185498 587342 185734
rect 587578 185498 587760 185734
rect 587160 150054 587760 185498
rect 587160 149818 587342 150054
rect 587578 149818 587760 150054
rect 587160 149734 587760 149818
rect 587160 149498 587342 149734
rect 587578 149498 587760 149734
rect 587160 114054 587760 149498
rect 587160 113818 587342 114054
rect 587578 113818 587760 114054
rect 587160 113734 587760 113818
rect 587160 113498 587342 113734
rect 587578 113498 587760 113734
rect 587160 78054 587760 113498
rect 587160 77818 587342 78054
rect 587578 77818 587760 78054
rect 587160 77734 587760 77818
rect 587160 77498 587342 77734
rect 587578 77498 587760 77734
rect 587160 42054 587760 77498
rect 587160 41818 587342 42054
rect 587578 41818 587760 42054
rect 587160 41734 587760 41818
rect 587160 41498 587342 41734
rect 587578 41498 587760 41734
rect 587160 6054 587760 41498
rect 587160 5818 587342 6054
rect 587578 5818 587760 6054
rect 587160 5734 587760 5818
rect 587160 5498 587342 5734
rect 587578 5498 587760 5734
rect 580404 -2422 580586 -2186
rect 580822 -2422 581004 -2186
rect 580404 -2506 581004 -2422
rect 580404 -2742 580586 -2506
rect 580822 -2742 581004 -2506
rect 580404 -3684 581004 -2742
rect 587160 -2186 587760 5498
rect 587160 -2422 587342 -2186
rect 587578 -2422 587760 -2186
rect 587160 -2506 587760 -2422
rect 587160 -2742 587342 -2506
rect 587578 -2742 587760 -2506
rect 587160 -2764 587760 -2742
rect 588080 672054 588680 707042
rect 588080 671818 588262 672054
rect 588498 671818 588680 672054
rect 588080 671734 588680 671818
rect 588080 671498 588262 671734
rect 588498 671498 588680 671734
rect 588080 636054 588680 671498
rect 588080 635818 588262 636054
rect 588498 635818 588680 636054
rect 588080 635734 588680 635818
rect 588080 635498 588262 635734
rect 588498 635498 588680 635734
rect 588080 600054 588680 635498
rect 588080 599818 588262 600054
rect 588498 599818 588680 600054
rect 588080 599734 588680 599818
rect 588080 599498 588262 599734
rect 588498 599498 588680 599734
rect 588080 564054 588680 599498
rect 588080 563818 588262 564054
rect 588498 563818 588680 564054
rect 588080 563734 588680 563818
rect 588080 563498 588262 563734
rect 588498 563498 588680 563734
rect 588080 528054 588680 563498
rect 588080 527818 588262 528054
rect 588498 527818 588680 528054
rect 588080 527734 588680 527818
rect 588080 527498 588262 527734
rect 588498 527498 588680 527734
rect 588080 492054 588680 527498
rect 588080 491818 588262 492054
rect 588498 491818 588680 492054
rect 588080 491734 588680 491818
rect 588080 491498 588262 491734
rect 588498 491498 588680 491734
rect 588080 456054 588680 491498
rect 588080 455818 588262 456054
rect 588498 455818 588680 456054
rect 588080 455734 588680 455818
rect 588080 455498 588262 455734
rect 588498 455498 588680 455734
rect 588080 420054 588680 455498
rect 588080 419818 588262 420054
rect 588498 419818 588680 420054
rect 588080 419734 588680 419818
rect 588080 419498 588262 419734
rect 588498 419498 588680 419734
rect 588080 384054 588680 419498
rect 588080 383818 588262 384054
rect 588498 383818 588680 384054
rect 588080 383734 588680 383818
rect 588080 383498 588262 383734
rect 588498 383498 588680 383734
rect 588080 348054 588680 383498
rect 588080 347818 588262 348054
rect 588498 347818 588680 348054
rect 588080 347734 588680 347818
rect 588080 347498 588262 347734
rect 588498 347498 588680 347734
rect 588080 312054 588680 347498
rect 588080 311818 588262 312054
rect 588498 311818 588680 312054
rect 588080 311734 588680 311818
rect 588080 311498 588262 311734
rect 588498 311498 588680 311734
rect 588080 276054 588680 311498
rect 588080 275818 588262 276054
rect 588498 275818 588680 276054
rect 588080 275734 588680 275818
rect 588080 275498 588262 275734
rect 588498 275498 588680 275734
rect 588080 240054 588680 275498
rect 588080 239818 588262 240054
rect 588498 239818 588680 240054
rect 588080 239734 588680 239818
rect 588080 239498 588262 239734
rect 588498 239498 588680 239734
rect 588080 204054 588680 239498
rect 588080 203818 588262 204054
rect 588498 203818 588680 204054
rect 588080 203734 588680 203818
rect 588080 203498 588262 203734
rect 588498 203498 588680 203734
rect 588080 168054 588680 203498
rect 588080 167818 588262 168054
rect 588498 167818 588680 168054
rect 588080 167734 588680 167818
rect 588080 167498 588262 167734
rect 588498 167498 588680 167734
rect 588080 132054 588680 167498
rect 588080 131818 588262 132054
rect 588498 131818 588680 132054
rect 588080 131734 588680 131818
rect 588080 131498 588262 131734
rect 588498 131498 588680 131734
rect 588080 96054 588680 131498
rect 588080 95818 588262 96054
rect 588498 95818 588680 96054
rect 588080 95734 588680 95818
rect 588080 95498 588262 95734
rect 588498 95498 588680 95734
rect 588080 60054 588680 95498
rect 588080 59818 588262 60054
rect 588498 59818 588680 60054
rect 588080 59734 588680 59818
rect 588080 59498 588262 59734
rect 588498 59498 588680 59734
rect 588080 24054 588680 59498
rect 588080 23818 588262 24054
rect 588498 23818 588680 24054
rect 588080 23734 588680 23818
rect 588080 23498 588262 23734
rect 588498 23498 588680 23734
rect 588080 -3106 588680 23498
rect 588080 -3342 588262 -3106
rect 588498 -3342 588680 -3106
rect 588080 -3426 588680 -3342
rect 588080 -3662 588262 -3426
rect 588498 -3662 588680 -3426
rect 588080 -3684 588680 -3662
rect 589000 693654 589600 707962
rect 589000 693418 589182 693654
rect 589418 693418 589600 693654
rect 589000 693334 589600 693418
rect 589000 693098 589182 693334
rect 589418 693098 589600 693334
rect 589000 657654 589600 693098
rect 589000 657418 589182 657654
rect 589418 657418 589600 657654
rect 589000 657334 589600 657418
rect 589000 657098 589182 657334
rect 589418 657098 589600 657334
rect 589000 621654 589600 657098
rect 589000 621418 589182 621654
rect 589418 621418 589600 621654
rect 589000 621334 589600 621418
rect 589000 621098 589182 621334
rect 589418 621098 589600 621334
rect 589000 585654 589600 621098
rect 589000 585418 589182 585654
rect 589418 585418 589600 585654
rect 589000 585334 589600 585418
rect 589000 585098 589182 585334
rect 589418 585098 589600 585334
rect 589000 549654 589600 585098
rect 589000 549418 589182 549654
rect 589418 549418 589600 549654
rect 589000 549334 589600 549418
rect 589000 549098 589182 549334
rect 589418 549098 589600 549334
rect 589000 513654 589600 549098
rect 589000 513418 589182 513654
rect 589418 513418 589600 513654
rect 589000 513334 589600 513418
rect 589000 513098 589182 513334
rect 589418 513098 589600 513334
rect 589000 477654 589600 513098
rect 589000 477418 589182 477654
rect 589418 477418 589600 477654
rect 589000 477334 589600 477418
rect 589000 477098 589182 477334
rect 589418 477098 589600 477334
rect 589000 441654 589600 477098
rect 589000 441418 589182 441654
rect 589418 441418 589600 441654
rect 589000 441334 589600 441418
rect 589000 441098 589182 441334
rect 589418 441098 589600 441334
rect 589000 405654 589600 441098
rect 589000 405418 589182 405654
rect 589418 405418 589600 405654
rect 589000 405334 589600 405418
rect 589000 405098 589182 405334
rect 589418 405098 589600 405334
rect 589000 369654 589600 405098
rect 589000 369418 589182 369654
rect 589418 369418 589600 369654
rect 589000 369334 589600 369418
rect 589000 369098 589182 369334
rect 589418 369098 589600 369334
rect 589000 333654 589600 369098
rect 589000 333418 589182 333654
rect 589418 333418 589600 333654
rect 589000 333334 589600 333418
rect 589000 333098 589182 333334
rect 589418 333098 589600 333334
rect 589000 297654 589600 333098
rect 589000 297418 589182 297654
rect 589418 297418 589600 297654
rect 589000 297334 589600 297418
rect 589000 297098 589182 297334
rect 589418 297098 589600 297334
rect 589000 261654 589600 297098
rect 589000 261418 589182 261654
rect 589418 261418 589600 261654
rect 589000 261334 589600 261418
rect 589000 261098 589182 261334
rect 589418 261098 589600 261334
rect 589000 225654 589600 261098
rect 589000 225418 589182 225654
rect 589418 225418 589600 225654
rect 589000 225334 589600 225418
rect 589000 225098 589182 225334
rect 589418 225098 589600 225334
rect 589000 189654 589600 225098
rect 589000 189418 589182 189654
rect 589418 189418 589600 189654
rect 589000 189334 589600 189418
rect 589000 189098 589182 189334
rect 589418 189098 589600 189334
rect 589000 153654 589600 189098
rect 589000 153418 589182 153654
rect 589418 153418 589600 153654
rect 589000 153334 589600 153418
rect 589000 153098 589182 153334
rect 589418 153098 589600 153334
rect 589000 117654 589600 153098
rect 589000 117418 589182 117654
rect 589418 117418 589600 117654
rect 589000 117334 589600 117418
rect 589000 117098 589182 117334
rect 589418 117098 589600 117334
rect 589000 81654 589600 117098
rect 589000 81418 589182 81654
rect 589418 81418 589600 81654
rect 589000 81334 589600 81418
rect 589000 81098 589182 81334
rect 589418 81098 589600 81334
rect 589000 45654 589600 81098
rect 589000 45418 589182 45654
rect 589418 45418 589600 45654
rect 589000 45334 589600 45418
rect 589000 45098 589182 45334
rect 589418 45098 589600 45334
rect 589000 9654 589600 45098
rect 589000 9418 589182 9654
rect 589418 9418 589600 9654
rect 589000 9334 589600 9418
rect 589000 9098 589182 9334
rect 589418 9098 589600 9334
rect 589000 -4026 589600 9098
rect 589000 -4262 589182 -4026
rect 589418 -4262 589600 -4026
rect 589000 -4346 589600 -4262
rect 589000 -4582 589182 -4346
rect 589418 -4582 589600 -4346
rect 589000 -4604 589600 -4582
rect 589920 675654 590520 708882
rect 589920 675418 590102 675654
rect 590338 675418 590520 675654
rect 589920 675334 590520 675418
rect 589920 675098 590102 675334
rect 590338 675098 590520 675334
rect 589920 639654 590520 675098
rect 589920 639418 590102 639654
rect 590338 639418 590520 639654
rect 589920 639334 590520 639418
rect 589920 639098 590102 639334
rect 590338 639098 590520 639334
rect 589920 603654 590520 639098
rect 589920 603418 590102 603654
rect 590338 603418 590520 603654
rect 589920 603334 590520 603418
rect 589920 603098 590102 603334
rect 590338 603098 590520 603334
rect 589920 567654 590520 603098
rect 589920 567418 590102 567654
rect 590338 567418 590520 567654
rect 589920 567334 590520 567418
rect 589920 567098 590102 567334
rect 590338 567098 590520 567334
rect 589920 531654 590520 567098
rect 589920 531418 590102 531654
rect 590338 531418 590520 531654
rect 589920 531334 590520 531418
rect 589920 531098 590102 531334
rect 590338 531098 590520 531334
rect 589920 495654 590520 531098
rect 589920 495418 590102 495654
rect 590338 495418 590520 495654
rect 589920 495334 590520 495418
rect 589920 495098 590102 495334
rect 590338 495098 590520 495334
rect 589920 459654 590520 495098
rect 589920 459418 590102 459654
rect 590338 459418 590520 459654
rect 589920 459334 590520 459418
rect 589920 459098 590102 459334
rect 590338 459098 590520 459334
rect 589920 423654 590520 459098
rect 589920 423418 590102 423654
rect 590338 423418 590520 423654
rect 589920 423334 590520 423418
rect 589920 423098 590102 423334
rect 590338 423098 590520 423334
rect 589920 387654 590520 423098
rect 589920 387418 590102 387654
rect 590338 387418 590520 387654
rect 589920 387334 590520 387418
rect 589920 387098 590102 387334
rect 590338 387098 590520 387334
rect 589920 351654 590520 387098
rect 589920 351418 590102 351654
rect 590338 351418 590520 351654
rect 589920 351334 590520 351418
rect 589920 351098 590102 351334
rect 590338 351098 590520 351334
rect 589920 315654 590520 351098
rect 589920 315418 590102 315654
rect 590338 315418 590520 315654
rect 589920 315334 590520 315418
rect 589920 315098 590102 315334
rect 590338 315098 590520 315334
rect 589920 279654 590520 315098
rect 589920 279418 590102 279654
rect 590338 279418 590520 279654
rect 589920 279334 590520 279418
rect 589920 279098 590102 279334
rect 590338 279098 590520 279334
rect 589920 243654 590520 279098
rect 589920 243418 590102 243654
rect 590338 243418 590520 243654
rect 589920 243334 590520 243418
rect 589920 243098 590102 243334
rect 590338 243098 590520 243334
rect 589920 207654 590520 243098
rect 589920 207418 590102 207654
rect 590338 207418 590520 207654
rect 589920 207334 590520 207418
rect 589920 207098 590102 207334
rect 590338 207098 590520 207334
rect 589920 171654 590520 207098
rect 589920 171418 590102 171654
rect 590338 171418 590520 171654
rect 589920 171334 590520 171418
rect 589920 171098 590102 171334
rect 590338 171098 590520 171334
rect 589920 135654 590520 171098
rect 589920 135418 590102 135654
rect 590338 135418 590520 135654
rect 589920 135334 590520 135418
rect 589920 135098 590102 135334
rect 590338 135098 590520 135334
rect 589920 99654 590520 135098
rect 589920 99418 590102 99654
rect 590338 99418 590520 99654
rect 589920 99334 590520 99418
rect 589920 99098 590102 99334
rect 590338 99098 590520 99334
rect 589920 63654 590520 99098
rect 589920 63418 590102 63654
rect 590338 63418 590520 63654
rect 589920 63334 590520 63418
rect 589920 63098 590102 63334
rect 590338 63098 590520 63334
rect 589920 27654 590520 63098
rect 589920 27418 590102 27654
rect 590338 27418 590520 27654
rect 589920 27334 590520 27418
rect 589920 27098 590102 27334
rect 590338 27098 590520 27334
rect 589920 -4946 590520 27098
rect 589920 -5182 590102 -4946
rect 590338 -5182 590520 -4946
rect 589920 -5266 590520 -5182
rect 589920 -5502 590102 -5266
rect 590338 -5502 590520 -5266
rect 589920 -5524 590520 -5502
rect 590840 697254 591440 709802
rect 590840 697018 591022 697254
rect 591258 697018 591440 697254
rect 590840 696934 591440 697018
rect 590840 696698 591022 696934
rect 591258 696698 591440 696934
rect 590840 661254 591440 696698
rect 590840 661018 591022 661254
rect 591258 661018 591440 661254
rect 590840 660934 591440 661018
rect 590840 660698 591022 660934
rect 591258 660698 591440 660934
rect 590840 625254 591440 660698
rect 590840 625018 591022 625254
rect 591258 625018 591440 625254
rect 590840 624934 591440 625018
rect 590840 624698 591022 624934
rect 591258 624698 591440 624934
rect 590840 589254 591440 624698
rect 590840 589018 591022 589254
rect 591258 589018 591440 589254
rect 590840 588934 591440 589018
rect 590840 588698 591022 588934
rect 591258 588698 591440 588934
rect 590840 553254 591440 588698
rect 590840 553018 591022 553254
rect 591258 553018 591440 553254
rect 590840 552934 591440 553018
rect 590840 552698 591022 552934
rect 591258 552698 591440 552934
rect 590840 517254 591440 552698
rect 590840 517018 591022 517254
rect 591258 517018 591440 517254
rect 590840 516934 591440 517018
rect 590840 516698 591022 516934
rect 591258 516698 591440 516934
rect 590840 481254 591440 516698
rect 590840 481018 591022 481254
rect 591258 481018 591440 481254
rect 590840 480934 591440 481018
rect 590840 480698 591022 480934
rect 591258 480698 591440 480934
rect 590840 445254 591440 480698
rect 590840 445018 591022 445254
rect 591258 445018 591440 445254
rect 590840 444934 591440 445018
rect 590840 444698 591022 444934
rect 591258 444698 591440 444934
rect 590840 409254 591440 444698
rect 590840 409018 591022 409254
rect 591258 409018 591440 409254
rect 590840 408934 591440 409018
rect 590840 408698 591022 408934
rect 591258 408698 591440 408934
rect 590840 373254 591440 408698
rect 590840 373018 591022 373254
rect 591258 373018 591440 373254
rect 590840 372934 591440 373018
rect 590840 372698 591022 372934
rect 591258 372698 591440 372934
rect 590840 337254 591440 372698
rect 590840 337018 591022 337254
rect 591258 337018 591440 337254
rect 590840 336934 591440 337018
rect 590840 336698 591022 336934
rect 591258 336698 591440 336934
rect 590840 301254 591440 336698
rect 590840 301018 591022 301254
rect 591258 301018 591440 301254
rect 590840 300934 591440 301018
rect 590840 300698 591022 300934
rect 591258 300698 591440 300934
rect 590840 265254 591440 300698
rect 590840 265018 591022 265254
rect 591258 265018 591440 265254
rect 590840 264934 591440 265018
rect 590840 264698 591022 264934
rect 591258 264698 591440 264934
rect 590840 229254 591440 264698
rect 590840 229018 591022 229254
rect 591258 229018 591440 229254
rect 590840 228934 591440 229018
rect 590840 228698 591022 228934
rect 591258 228698 591440 228934
rect 590840 193254 591440 228698
rect 590840 193018 591022 193254
rect 591258 193018 591440 193254
rect 590840 192934 591440 193018
rect 590840 192698 591022 192934
rect 591258 192698 591440 192934
rect 590840 157254 591440 192698
rect 590840 157018 591022 157254
rect 591258 157018 591440 157254
rect 590840 156934 591440 157018
rect 590840 156698 591022 156934
rect 591258 156698 591440 156934
rect 590840 121254 591440 156698
rect 590840 121018 591022 121254
rect 591258 121018 591440 121254
rect 590840 120934 591440 121018
rect 590840 120698 591022 120934
rect 591258 120698 591440 120934
rect 590840 85254 591440 120698
rect 590840 85018 591022 85254
rect 591258 85018 591440 85254
rect 590840 84934 591440 85018
rect 590840 84698 591022 84934
rect 591258 84698 591440 84934
rect 590840 49254 591440 84698
rect 590840 49018 591022 49254
rect 591258 49018 591440 49254
rect 590840 48934 591440 49018
rect 590840 48698 591022 48934
rect 591258 48698 591440 48934
rect 590840 13254 591440 48698
rect 590840 13018 591022 13254
rect 591258 13018 591440 13254
rect 590840 12934 591440 13018
rect 590840 12698 591022 12934
rect 591258 12698 591440 12934
rect 590840 -5866 591440 12698
rect 590840 -6102 591022 -5866
rect 591258 -6102 591440 -5866
rect 590840 -6186 591440 -6102
rect 590840 -6422 591022 -6186
rect 591258 -6422 591440 -6186
rect 590840 -6444 591440 -6422
rect 591760 679254 592360 710722
rect 591760 679018 591942 679254
rect 592178 679018 592360 679254
rect 591760 678934 592360 679018
rect 591760 678698 591942 678934
rect 592178 678698 592360 678934
rect 591760 643254 592360 678698
rect 591760 643018 591942 643254
rect 592178 643018 592360 643254
rect 591760 642934 592360 643018
rect 591760 642698 591942 642934
rect 592178 642698 592360 642934
rect 591760 607254 592360 642698
rect 591760 607018 591942 607254
rect 592178 607018 592360 607254
rect 591760 606934 592360 607018
rect 591760 606698 591942 606934
rect 592178 606698 592360 606934
rect 591760 571254 592360 606698
rect 591760 571018 591942 571254
rect 592178 571018 592360 571254
rect 591760 570934 592360 571018
rect 591760 570698 591942 570934
rect 592178 570698 592360 570934
rect 591760 535254 592360 570698
rect 591760 535018 591942 535254
rect 592178 535018 592360 535254
rect 591760 534934 592360 535018
rect 591760 534698 591942 534934
rect 592178 534698 592360 534934
rect 591760 499254 592360 534698
rect 591760 499018 591942 499254
rect 592178 499018 592360 499254
rect 591760 498934 592360 499018
rect 591760 498698 591942 498934
rect 592178 498698 592360 498934
rect 591760 463254 592360 498698
rect 591760 463018 591942 463254
rect 592178 463018 592360 463254
rect 591760 462934 592360 463018
rect 591760 462698 591942 462934
rect 592178 462698 592360 462934
rect 591760 427254 592360 462698
rect 591760 427018 591942 427254
rect 592178 427018 592360 427254
rect 591760 426934 592360 427018
rect 591760 426698 591942 426934
rect 592178 426698 592360 426934
rect 591760 391254 592360 426698
rect 591760 391018 591942 391254
rect 592178 391018 592360 391254
rect 591760 390934 592360 391018
rect 591760 390698 591942 390934
rect 592178 390698 592360 390934
rect 591760 355254 592360 390698
rect 591760 355018 591942 355254
rect 592178 355018 592360 355254
rect 591760 354934 592360 355018
rect 591760 354698 591942 354934
rect 592178 354698 592360 354934
rect 591760 319254 592360 354698
rect 591760 319018 591942 319254
rect 592178 319018 592360 319254
rect 591760 318934 592360 319018
rect 591760 318698 591942 318934
rect 592178 318698 592360 318934
rect 591760 283254 592360 318698
rect 591760 283018 591942 283254
rect 592178 283018 592360 283254
rect 591760 282934 592360 283018
rect 591760 282698 591942 282934
rect 592178 282698 592360 282934
rect 591760 247254 592360 282698
rect 591760 247018 591942 247254
rect 592178 247018 592360 247254
rect 591760 246934 592360 247018
rect 591760 246698 591942 246934
rect 592178 246698 592360 246934
rect 591760 211254 592360 246698
rect 591760 211018 591942 211254
rect 592178 211018 592360 211254
rect 591760 210934 592360 211018
rect 591760 210698 591942 210934
rect 592178 210698 592360 210934
rect 591760 175254 592360 210698
rect 591760 175018 591942 175254
rect 592178 175018 592360 175254
rect 591760 174934 592360 175018
rect 591760 174698 591942 174934
rect 592178 174698 592360 174934
rect 591760 139254 592360 174698
rect 591760 139018 591942 139254
rect 592178 139018 592360 139254
rect 591760 138934 592360 139018
rect 591760 138698 591942 138934
rect 592178 138698 592360 138934
rect 591760 103254 592360 138698
rect 591760 103018 591942 103254
rect 592178 103018 592360 103254
rect 591760 102934 592360 103018
rect 591760 102698 591942 102934
rect 592178 102698 592360 102934
rect 591760 67254 592360 102698
rect 591760 67018 591942 67254
rect 592178 67018 592360 67254
rect 591760 66934 592360 67018
rect 591760 66698 591942 66934
rect 592178 66698 592360 66934
rect 591760 31254 592360 66698
rect 591760 31018 591942 31254
rect 592178 31018 592360 31254
rect 591760 30934 592360 31018
rect 591760 30698 591942 30934
rect 592178 30698 592360 30934
rect 569604 -7022 569786 -6786
rect 570022 -7022 570204 -6786
rect 569604 -7106 570204 -7022
rect 569604 -7342 569786 -7106
rect 570022 -7342 570204 -7106
rect 569604 -7364 570204 -7342
rect 591760 -6786 592360 30698
rect 591760 -7022 591942 -6786
rect 592178 -7022 592360 -6786
rect 591760 -7106 592360 -7022
rect 591760 -7342 591942 -7106
rect 592178 -7342 592360 -7106
rect 591760 -7364 592360 -7342
<< via4 >>
rect -8254 711042 -8018 711278
rect -8254 710722 -8018 710958
rect -8254 679018 -8018 679254
rect -8254 678698 -8018 678934
rect -8254 643018 -8018 643254
rect -8254 642698 -8018 642934
rect -8254 607018 -8018 607254
rect -8254 606698 -8018 606934
rect -8254 571018 -8018 571254
rect -8254 570698 -8018 570934
rect -8254 535018 -8018 535254
rect -8254 534698 -8018 534934
rect -8254 499018 -8018 499254
rect -8254 498698 -8018 498934
rect -8254 463018 -8018 463254
rect -8254 462698 -8018 462934
rect -8254 427018 -8018 427254
rect -8254 426698 -8018 426934
rect -8254 391018 -8018 391254
rect -8254 390698 -8018 390934
rect -8254 355018 -8018 355254
rect -8254 354698 -8018 354934
rect -8254 319018 -8018 319254
rect -8254 318698 -8018 318934
rect -8254 283018 -8018 283254
rect -8254 282698 -8018 282934
rect -8254 247018 -8018 247254
rect -8254 246698 -8018 246934
rect -8254 211018 -8018 211254
rect -8254 210698 -8018 210934
rect -8254 175018 -8018 175254
rect -8254 174698 -8018 174934
rect -8254 139018 -8018 139254
rect -8254 138698 -8018 138934
rect -8254 103018 -8018 103254
rect -8254 102698 -8018 102934
rect -8254 67018 -8018 67254
rect -8254 66698 -8018 66934
rect -8254 31018 -8018 31254
rect -8254 30698 -8018 30934
rect -7334 710122 -7098 710358
rect -7334 709802 -7098 710038
rect 11786 710122 12022 710358
rect 11786 709802 12022 710038
rect -7334 697018 -7098 697254
rect -7334 696698 -7098 696934
rect -7334 661018 -7098 661254
rect -7334 660698 -7098 660934
rect -7334 625018 -7098 625254
rect -7334 624698 -7098 624934
rect -7334 589018 -7098 589254
rect -7334 588698 -7098 588934
rect -7334 553018 -7098 553254
rect -7334 552698 -7098 552934
rect -7334 517018 -7098 517254
rect -7334 516698 -7098 516934
rect -7334 481018 -7098 481254
rect -7334 480698 -7098 480934
rect -7334 445018 -7098 445254
rect -7334 444698 -7098 444934
rect -7334 409018 -7098 409254
rect -7334 408698 -7098 408934
rect -7334 373018 -7098 373254
rect -7334 372698 -7098 372934
rect -7334 337018 -7098 337254
rect -7334 336698 -7098 336934
rect -7334 301018 -7098 301254
rect -7334 300698 -7098 300934
rect -7334 265018 -7098 265254
rect -7334 264698 -7098 264934
rect -7334 229018 -7098 229254
rect -7334 228698 -7098 228934
rect -7334 193018 -7098 193254
rect -7334 192698 -7098 192934
rect -7334 157018 -7098 157254
rect -7334 156698 -7098 156934
rect -7334 121018 -7098 121254
rect -7334 120698 -7098 120934
rect -7334 85018 -7098 85254
rect -7334 84698 -7098 84934
rect -7334 49018 -7098 49254
rect -7334 48698 -7098 48934
rect -7334 13018 -7098 13254
rect -7334 12698 -7098 12934
rect -6414 709202 -6178 709438
rect -6414 708882 -6178 709118
rect -6414 675418 -6178 675654
rect -6414 675098 -6178 675334
rect -6414 639418 -6178 639654
rect -6414 639098 -6178 639334
rect -6414 603418 -6178 603654
rect -6414 603098 -6178 603334
rect -6414 567418 -6178 567654
rect -6414 567098 -6178 567334
rect -6414 531418 -6178 531654
rect -6414 531098 -6178 531334
rect -6414 495418 -6178 495654
rect -6414 495098 -6178 495334
rect -6414 459418 -6178 459654
rect -6414 459098 -6178 459334
rect -6414 423418 -6178 423654
rect -6414 423098 -6178 423334
rect -6414 387418 -6178 387654
rect -6414 387098 -6178 387334
rect -6414 351418 -6178 351654
rect -6414 351098 -6178 351334
rect -6414 315418 -6178 315654
rect -6414 315098 -6178 315334
rect -6414 279418 -6178 279654
rect -6414 279098 -6178 279334
rect -6414 243418 -6178 243654
rect -6414 243098 -6178 243334
rect -6414 207418 -6178 207654
rect -6414 207098 -6178 207334
rect -6414 171418 -6178 171654
rect -6414 171098 -6178 171334
rect -6414 135418 -6178 135654
rect -6414 135098 -6178 135334
rect -6414 99418 -6178 99654
rect -6414 99098 -6178 99334
rect -6414 63418 -6178 63654
rect -6414 63098 -6178 63334
rect -6414 27418 -6178 27654
rect -6414 27098 -6178 27334
rect -5494 708282 -5258 708518
rect -5494 707962 -5258 708198
rect 8186 708282 8422 708518
rect 8186 707962 8422 708198
rect -5494 693418 -5258 693654
rect -5494 693098 -5258 693334
rect -5494 657418 -5258 657654
rect -5494 657098 -5258 657334
rect -5494 621418 -5258 621654
rect -5494 621098 -5258 621334
rect -5494 585418 -5258 585654
rect -5494 585098 -5258 585334
rect -5494 549418 -5258 549654
rect -5494 549098 -5258 549334
rect -5494 513418 -5258 513654
rect -5494 513098 -5258 513334
rect -5494 477418 -5258 477654
rect -5494 477098 -5258 477334
rect -5494 441418 -5258 441654
rect -5494 441098 -5258 441334
rect -5494 405418 -5258 405654
rect -5494 405098 -5258 405334
rect -5494 369418 -5258 369654
rect -5494 369098 -5258 369334
rect -5494 333418 -5258 333654
rect -5494 333098 -5258 333334
rect -5494 297418 -5258 297654
rect -5494 297098 -5258 297334
rect -5494 261418 -5258 261654
rect -5494 261098 -5258 261334
rect -5494 225418 -5258 225654
rect -5494 225098 -5258 225334
rect -5494 189418 -5258 189654
rect -5494 189098 -5258 189334
rect -5494 153418 -5258 153654
rect -5494 153098 -5258 153334
rect -5494 117418 -5258 117654
rect -5494 117098 -5258 117334
rect -5494 81418 -5258 81654
rect -5494 81098 -5258 81334
rect -5494 45418 -5258 45654
rect -5494 45098 -5258 45334
rect -5494 9418 -5258 9654
rect -5494 9098 -5258 9334
rect -4574 707362 -4338 707598
rect -4574 707042 -4338 707278
rect -4574 671818 -4338 672054
rect -4574 671498 -4338 671734
rect -4574 635818 -4338 636054
rect -4574 635498 -4338 635734
rect -4574 599818 -4338 600054
rect -4574 599498 -4338 599734
rect -4574 563818 -4338 564054
rect -4574 563498 -4338 563734
rect -4574 527818 -4338 528054
rect -4574 527498 -4338 527734
rect -4574 491818 -4338 492054
rect -4574 491498 -4338 491734
rect -4574 455818 -4338 456054
rect -4574 455498 -4338 455734
rect -4574 419818 -4338 420054
rect -4574 419498 -4338 419734
rect -4574 383818 -4338 384054
rect -4574 383498 -4338 383734
rect -4574 347818 -4338 348054
rect -4574 347498 -4338 347734
rect -4574 311818 -4338 312054
rect -4574 311498 -4338 311734
rect -4574 275818 -4338 276054
rect -4574 275498 -4338 275734
rect -4574 239818 -4338 240054
rect -4574 239498 -4338 239734
rect -4574 203818 -4338 204054
rect -4574 203498 -4338 203734
rect -4574 167818 -4338 168054
rect -4574 167498 -4338 167734
rect -4574 131818 -4338 132054
rect -4574 131498 -4338 131734
rect -4574 95818 -4338 96054
rect -4574 95498 -4338 95734
rect -4574 59818 -4338 60054
rect -4574 59498 -4338 59734
rect -4574 23818 -4338 24054
rect -4574 23498 -4338 23734
rect -3654 706442 -3418 706678
rect -3654 706122 -3418 706358
rect 4586 706442 4822 706678
rect 4586 706122 4822 706358
rect -3654 689818 -3418 690054
rect -3654 689498 -3418 689734
rect -3654 653818 -3418 654054
rect -3654 653498 -3418 653734
rect -3654 617818 -3418 618054
rect -3654 617498 -3418 617734
rect -3654 581818 -3418 582054
rect -3654 581498 -3418 581734
rect -3654 545818 -3418 546054
rect -3654 545498 -3418 545734
rect -3654 509818 -3418 510054
rect -3654 509498 -3418 509734
rect -3654 473818 -3418 474054
rect -3654 473498 -3418 473734
rect -3654 437818 -3418 438054
rect -3654 437498 -3418 437734
rect -3654 401818 -3418 402054
rect -3654 401498 -3418 401734
rect -3654 365818 -3418 366054
rect -3654 365498 -3418 365734
rect -3654 329818 -3418 330054
rect -3654 329498 -3418 329734
rect -3654 293818 -3418 294054
rect -3654 293498 -3418 293734
rect -3654 257818 -3418 258054
rect -3654 257498 -3418 257734
rect -3654 221818 -3418 222054
rect -3654 221498 -3418 221734
rect -3654 185818 -3418 186054
rect -3654 185498 -3418 185734
rect -3654 149818 -3418 150054
rect -3654 149498 -3418 149734
rect -3654 113818 -3418 114054
rect -3654 113498 -3418 113734
rect -3654 77818 -3418 78054
rect -3654 77498 -3418 77734
rect -3654 41818 -3418 42054
rect -3654 41498 -3418 41734
rect -3654 5818 -3418 6054
rect -3654 5498 -3418 5734
rect -2734 705522 -2498 705758
rect -2734 705202 -2498 705438
rect -2734 668218 -2498 668454
rect -2734 667898 -2498 668134
rect -2734 632218 -2498 632454
rect -2734 631898 -2498 632134
rect -2734 596218 -2498 596454
rect -2734 595898 -2498 596134
rect -2734 560218 -2498 560454
rect -2734 559898 -2498 560134
rect -2734 524218 -2498 524454
rect -2734 523898 -2498 524134
rect -2734 488218 -2498 488454
rect -2734 487898 -2498 488134
rect -2734 452218 -2498 452454
rect -2734 451898 -2498 452134
rect -2734 416218 -2498 416454
rect -2734 415898 -2498 416134
rect -2734 380218 -2498 380454
rect -2734 379898 -2498 380134
rect -2734 344218 -2498 344454
rect -2734 343898 -2498 344134
rect -2734 308218 -2498 308454
rect -2734 307898 -2498 308134
rect -2734 272218 -2498 272454
rect -2734 271898 -2498 272134
rect -2734 236218 -2498 236454
rect -2734 235898 -2498 236134
rect -2734 200218 -2498 200454
rect -2734 199898 -2498 200134
rect -2734 164218 -2498 164454
rect -2734 163898 -2498 164134
rect -2734 128218 -2498 128454
rect -2734 127898 -2498 128134
rect -2734 92218 -2498 92454
rect -2734 91898 -2498 92134
rect -2734 56218 -2498 56454
rect -2734 55898 -2498 56134
rect -2734 20218 -2498 20454
rect -2734 19898 -2498 20134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 686218 -1578 686454
rect -1814 685898 -1578 686134
rect -1814 650218 -1578 650454
rect -1814 649898 -1578 650134
rect -1814 614218 -1578 614454
rect -1814 613898 -1578 614134
rect -1814 578218 -1578 578454
rect -1814 577898 -1578 578134
rect -1814 542218 -1578 542454
rect -1814 541898 -1578 542134
rect -1814 506218 -1578 506454
rect -1814 505898 -1578 506134
rect -1814 470218 -1578 470454
rect -1814 469898 -1578 470134
rect -1814 434218 -1578 434454
rect -1814 433898 -1578 434134
rect -1814 398218 -1578 398454
rect -1814 397898 -1578 398134
rect -1814 362218 -1578 362454
rect -1814 361898 -1578 362134
rect -1814 326218 -1578 326454
rect -1814 325898 -1578 326134
rect -1814 290218 -1578 290454
rect -1814 289898 -1578 290134
rect -1814 254218 -1578 254454
rect -1814 253898 -1578 254134
rect -1814 218218 -1578 218454
rect -1814 217898 -1578 218134
rect -1814 182218 -1578 182454
rect -1814 181898 -1578 182134
rect -1814 146218 -1578 146454
rect -1814 145898 -1578 146134
rect -1814 110218 -1578 110454
rect -1814 109898 -1578 110134
rect -1814 74218 -1578 74454
rect -1814 73898 -1578 74134
rect -1814 38218 -1578 38454
rect -1814 37898 -1578 38134
rect -1814 2218 -1578 2454
rect -1814 1898 -1578 2134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 986 686218 1222 686454
rect 986 685898 1222 686134
rect 986 650218 1222 650454
rect 986 649898 1222 650134
rect 986 614218 1222 614454
rect 986 613898 1222 614134
rect 986 578218 1222 578454
rect 986 577898 1222 578134
rect 986 542218 1222 542454
rect 986 541898 1222 542134
rect 986 506218 1222 506454
rect 986 505898 1222 506134
rect 986 470218 1222 470454
rect 986 469898 1222 470134
rect 986 434218 1222 434454
rect 986 433898 1222 434134
rect 986 398218 1222 398454
rect 986 397898 1222 398134
rect 986 362218 1222 362454
rect 986 361898 1222 362134
rect 986 326218 1222 326454
rect 986 325898 1222 326134
rect 986 290218 1222 290454
rect 986 289898 1222 290134
rect 986 254218 1222 254454
rect 986 253898 1222 254134
rect 986 218218 1222 218454
rect 986 217898 1222 218134
rect 986 182218 1222 182454
rect 986 181898 1222 182134
rect 986 146218 1222 146454
rect 986 145898 1222 146134
rect 986 110218 1222 110454
rect 986 109898 1222 110134
rect 986 74218 1222 74454
rect 986 73898 1222 74134
rect 986 38218 1222 38454
rect 986 37898 1222 38134
rect 986 2218 1222 2454
rect 986 1898 1222 2134
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2734 -1502 -2498 -1266
rect -2734 -1822 -2498 -1586
rect 4586 689818 4822 690054
rect 4586 689498 4822 689734
rect 4586 653818 4822 654054
rect 4586 653498 4822 653734
rect 4586 617818 4822 618054
rect 4586 617498 4822 617734
rect 4586 581818 4822 582054
rect 4586 581498 4822 581734
rect 4586 545818 4822 546054
rect 4586 545498 4822 545734
rect 4586 509818 4822 510054
rect 4586 509498 4822 509734
rect 4586 473818 4822 474054
rect 4586 473498 4822 473734
rect 4586 437818 4822 438054
rect 4586 437498 4822 437734
rect 4586 401818 4822 402054
rect 4586 401498 4822 401734
rect 4586 365818 4822 366054
rect 4586 365498 4822 365734
rect 4586 329818 4822 330054
rect 4586 329498 4822 329734
rect 4586 293818 4822 294054
rect 4586 293498 4822 293734
rect 4586 257818 4822 258054
rect 4586 257498 4822 257734
rect 4586 221818 4822 222054
rect 4586 221498 4822 221734
rect 4586 185818 4822 186054
rect 4586 185498 4822 185734
rect 4586 149818 4822 150054
rect 4586 149498 4822 149734
rect 4586 113818 4822 114054
rect 4586 113498 4822 113734
rect 4586 77818 4822 78054
rect 4586 77498 4822 77734
rect 4586 41818 4822 42054
rect 4586 41498 4822 41734
rect 4586 5818 4822 6054
rect 4586 5498 4822 5734
rect -3654 -2422 -3418 -2186
rect -3654 -2742 -3418 -2506
rect 4586 -2422 4822 -2186
rect 4586 -2742 4822 -2506
rect -4574 -3342 -4338 -3106
rect -4574 -3662 -4338 -3426
rect 8186 693418 8422 693654
rect 8186 693098 8422 693334
rect 8186 657418 8422 657654
rect 8186 657098 8422 657334
rect 8186 621418 8422 621654
rect 8186 621098 8422 621334
rect 8186 585418 8422 585654
rect 8186 585098 8422 585334
rect 8186 549418 8422 549654
rect 8186 549098 8422 549334
rect 8186 513418 8422 513654
rect 8186 513098 8422 513334
rect 8186 477418 8422 477654
rect 8186 477098 8422 477334
rect 8186 441418 8422 441654
rect 8186 441098 8422 441334
rect 8186 405418 8422 405654
rect 8186 405098 8422 405334
rect 8186 369418 8422 369654
rect 8186 369098 8422 369334
rect 8186 333418 8422 333654
rect 8186 333098 8422 333334
rect 8186 297418 8422 297654
rect 8186 297098 8422 297334
rect 8186 261418 8422 261654
rect 8186 261098 8422 261334
rect 8186 225418 8422 225654
rect 8186 225098 8422 225334
rect 8186 189418 8422 189654
rect 8186 189098 8422 189334
rect 8186 153418 8422 153654
rect 8186 153098 8422 153334
rect 8186 117418 8422 117654
rect 8186 117098 8422 117334
rect 8186 81418 8422 81654
rect 8186 81098 8422 81334
rect 8186 45418 8422 45654
rect 8186 45098 8422 45334
rect 8186 9418 8422 9654
rect 8186 9098 8422 9334
rect -5494 -4262 -5258 -4026
rect -5494 -4582 -5258 -4346
rect 8186 -4262 8422 -4026
rect 8186 -4582 8422 -4346
rect -6414 -5182 -6178 -4946
rect -6414 -5502 -6178 -5266
rect 29786 711042 30022 711278
rect 29786 710722 30022 710958
rect 26186 709202 26422 709438
rect 26186 708882 26422 709118
rect 22586 707362 22822 707598
rect 22586 707042 22822 707278
rect 11786 697018 12022 697254
rect 11786 696698 12022 696934
rect 11786 661018 12022 661254
rect 11786 660698 12022 660934
rect 11786 625018 12022 625254
rect 11786 624698 12022 624934
rect 11786 589018 12022 589254
rect 11786 588698 12022 588934
rect 11786 553018 12022 553254
rect 11786 552698 12022 552934
rect 11786 517018 12022 517254
rect 11786 516698 12022 516934
rect 11786 481018 12022 481254
rect 11786 480698 12022 480934
rect 11786 445018 12022 445254
rect 11786 444698 12022 444934
rect 11786 409018 12022 409254
rect 11786 408698 12022 408934
rect 11786 373018 12022 373254
rect 11786 372698 12022 372934
rect 11786 337018 12022 337254
rect 11786 336698 12022 336934
rect 11786 301018 12022 301254
rect 11786 300698 12022 300934
rect 11786 265018 12022 265254
rect 11786 264698 12022 264934
rect 11786 229018 12022 229254
rect 11786 228698 12022 228934
rect 11786 193018 12022 193254
rect 11786 192698 12022 192934
rect 11786 157018 12022 157254
rect 11786 156698 12022 156934
rect 11786 121018 12022 121254
rect 11786 120698 12022 120934
rect 11786 85018 12022 85254
rect 11786 84698 12022 84934
rect 11786 49018 12022 49254
rect 11786 48698 12022 48934
rect 11786 13018 12022 13254
rect 11786 12698 12022 12934
rect -7334 -6102 -7098 -5866
rect -7334 -6422 -7098 -6186
rect 18986 705522 19222 705758
rect 18986 705202 19222 705438
rect 18986 668218 19222 668454
rect 18986 667898 19222 668134
rect 18986 632218 19222 632454
rect 18986 631898 19222 632134
rect 18986 596218 19222 596454
rect 18986 595898 19222 596134
rect 18986 560218 19222 560454
rect 18986 559898 19222 560134
rect 18986 524218 19222 524454
rect 18986 523898 19222 524134
rect 18986 488218 19222 488454
rect 18986 487898 19222 488134
rect 18986 452218 19222 452454
rect 18986 451898 19222 452134
rect 18986 416218 19222 416454
rect 18986 415898 19222 416134
rect 18986 380218 19222 380454
rect 18986 379898 19222 380134
rect 18986 344218 19222 344454
rect 18986 343898 19222 344134
rect 18986 308218 19222 308454
rect 18986 307898 19222 308134
rect 18986 272218 19222 272454
rect 18986 271898 19222 272134
rect 18986 236218 19222 236454
rect 18986 235898 19222 236134
rect 18986 200218 19222 200454
rect 18986 199898 19222 200134
rect 18986 164218 19222 164454
rect 18986 163898 19222 164134
rect 18986 128218 19222 128454
rect 18986 127898 19222 128134
rect 18986 92218 19222 92454
rect 18986 91898 19222 92134
rect 18986 56218 19222 56454
rect 18986 55898 19222 56134
rect 18986 20218 19222 20454
rect 18986 19898 19222 20134
rect 18986 -1502 19222 -1266
rect 18986 -1822 19222 -1586
rect 22586 671818 22822 672054
rect 22586 671498 22822 671734
rect 22586 635818 22822 636054
rect 22586 635498 22822 635734
rect 22586 599818 22822 600054
rect 22586 599498 22822 599734
rect 22586 563818 22822 564054
rect 22586 563498 22822 563734
rect 22586 527818 22822 528054
rect 22586 527498 22822 527734
rect 22586 491818 22822 492054
rect 22586 491498 22822 491734
rect 22586 455818 22822 456054
rect 22586 455498 22822 455734
rect 22586 419818 22822 420054
rect 22586 419498 22822 419734
rect 22586 383818 22822 384054
rect 22586 383498 22822 383734
rect 22586 347818 22822 348054
rect 22586 347498 22822 347734
rect 22586 311818 22822 312054
rect 22586 311498 22822 311734
rect 22586 275818 22822 276054
rect 22586 275498 22822 275734
rect 22586 239818 22822 240054
rect 22586 239498 22822 239734
rect 22586 203818 22822 204054
rect 22586 203498 22822 203734
rect 22586 167818 22822 168054
rect 22586 167498 22822 167734
rect 22586 131818 22822 132054
rect 22586 131498 22822 131734
rect 22586 95818 22822 96054
rect 22586 95498 22822 95734
rect 22586 59818 22822 60054
rect 22586 59498 22822 59734
rect 22586 23818 22822 24054
rect 22586 23498 22822 23734
rect 22586 -3342 22822 -3106
rect 22586 -3662 22822 -3426
rect 26186 675418 26422 675654
rect 26186 675098 26422 675334
rect 26186 639418 26422 639654
rect 26186 639098 26422 639334
rect 26186 603418 26422 603654
rect 26186 603098 26422 603334
rect 26186 567418 26422 567654
rect 26186 567098 26422 567334
rect 26186 531418 26422 531654
rect 26186 531098 26422 531334
rect 26186 495418 26422 495654
rect 26186 495098 26422 495334
rect 26186 459418 26422 459654
rect 26186 459098 26422 459334
rect 26186 423418 26422 423654
rect 26186 423098 26422 423334
rect 26186 387418 26422 387654
rect 26186 387098 26422 387334
rect 26186 351418 26422 351654
rect 26186 351098 26422 351334
rect 26186 315418 26422 315654
rect 26186 315098 26422 315334
rect 26186 279418 26422 279654
rect 26186 279098 26422 279334
rect 26186 243418 26422 243654
rect 26186 243098 26422 243334
rect 26186 207418 26422 207654
rect 26186 207098 26422 207334
rect 26186 171418 26422 171654
rect 26186 171098 26422 171334
rect 26186 135418 26422 135654
rect 26186 135098 26422 135334
rect 26186 99418 26422 99654
rect 26186 99098 26422 99334
rect 26186 63418 26422 63654
rect 26186 63098 26422 63334
rect 26186 27418 26422 27654
rect 26186 27098 26422 27334
rect 26186 -5182 26422 -4946
rect 26186 -5502 26422 -5266
rect 47786 710122 48022 710358
rect 47786 709802 48022 710038
rect 44186 708282 44422 708518
rect 44186 707962 44422 708198
rect 40586 706442 40822 706678
rect 40586 706122 40822 706358
rect 29786 679018 30022 679254
rect 29786 678698 30022 678934
rect 29786 643018 30022 643254
rect 29786 642698 30022 642934
rect 29786 607018 30022 607254
rect 29786 606698 30022 606934
rect 29786 571018 30022 571254
rect 29786 570698 30022 570934
rect 29786 535018 30022 535254
rect 29786 534698 30022 534934
rect 29786 499018 30022 499254
rect 29786 498698 30022 498934
rect 29786 463018 30022 463254
rect 29786 462698 30022 462934
rect 29786 427018 30022 427254
rect 29786 426698 30022 426934
rect 29786 391018 30022 391254
rect 29786 390698 30022 390934
rect 29786 355018 30022 355254
rect 29786 354698 30022 354934
rect 29786 319018 30022 319254
rect 29786 318698 30022 318934
rect 29786 283018 30022 283254
rect 29786 282698 30022 282934
rect 29786 247018 30022 247254
rect 29786 246698 30022 246934
rect 29786 211018 30022 211254
rect 29786 210698 30022 210934
rect 29786 175018 30022 175254
rect 29786 174698 30022 174934
rect 29786 139018 30022 139254
rect 29786 138698 30022 138934
rect 29786 103018 30022 103254
rect 29786 102698 30022 102934
rect 29786 67018 30022 67254
rect 29786 66698 30022 66934
rect 29786 31018 30022 31254
rect 29786 30698 30022 30934
rect 11786 -6102 12022 -5866
rect 11786 -6422 12022 -6186
rect -8254 -7022 -8018 -6786
rect -8254 -7342 -8018 -7106
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect 36986 686218 37222 686454
rect 36986 685898 37222 686134
rect 36986 650218 37222 650454
rect 36986 649898 37222 650134
rect 36986 614218 37222 614454
rect 36986 613898 37222 614134
rect 36986 578218 37222 578454
rect 36986 577898 37222 578134
rect 36986 542218 37222 542454
rect 36986 541898 37222 542134
rect 36986 506218 37222 506454
rect 36986 505898 37222 506134
rect 36986 470218 37222 470454
rect 36986 469898 37222 470134
rect 36986 434218 37222 434454
rect 36986 433898 37222 434134
rect 36986 398218 37222 398454
rect 36986 397898 37222 398134
rect 36986 362218 37222 362454
rect 36986 361898 37222 362134
rect 36986 326218 37222 326454
rect 36986 325898 37222 326134
rect 36986 290218 37222 290454
rect 36986 289898 37222 290134
rect 36986 254218 37222 254454
rect 36986 253898 37222 254134
rect 36986 218218 37222 218454
rect 36986 217898 37222 218134
rect 36986 182218 37222 182454
rect 36986 181898 37222 182134
rect 36986 146218 37222 146454
rect 36986 145898 37222 146134
rect 36986 110218 37222 110454
rect 36986 109898 37222 110134
rect 36986 74218 37222 74454
rect 36986 73898 37222 74134
rect 36986 38218 37222 38454
rect 36986 37898 37222 38134
rect 36986 2218 37222 2454
rect 36986 1898 37222 2134
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 40586 689818 40822 690054
rect 40586 689498 40822 689734
rect 40586 653818 40822 654054
rect 40586 653498 40822 653734
rect 40586 617818 40822 618054
rect 40586 617498 40822 617734
rect 40586 581818 40822 582054
rect 40586 581498 40822 581734
rect 40586 545818 40822 546054
rect 40586 545498 40822 545734
rect 40586 509818 40822 510054
rect 40586 509498 40822 509734
rect 40586 473818 40822 474054
rect 40586 473498 40822 473734
rect 40586 437818 40822 438054
rect 40586 437498 40822 437734
rect 40586 401818 40822 402054
rect 40586 401498 40822 401734
rect 40586 365818 40822 366054
rect 40586 365498 40822 365734
rect 40586 329818 40822 330054
rect 40586 329498 40822 329734
rect 40586 293818 40822 294054
rect 40586 293498 40822 293734
rect 40586 257818 40822 258054
rect 40586 257498 40822 257734
rect 40586 221818 40822 222054
rect 40586 221498 40822 221734
rect 40586 185818 40822 186054
rect 40586 185498 40822 185734
rect 40586 149818 40822 150054
rect 40586 149498 40822 149734
rect 40586 113818 40822 114054
rect 40586 113498 40822 113734
rect 40586 77818 40822 78054
rect 40586 77498 40822 77734
rect 40586 41818 40822 42054
rect 40586 41498 40822 41734
rect 40586 5818 40822 6054
rect 40586 5498 40822 5734
rect 40586 -2422 40822 -2186
rect 40586 -2742 40822 -2506
rect 44186 693418 44422 693654
rect 44186 693098 44422 693334
rect 44186 657418 44422 657654
rect 44186 657098 44422 657334
rect 44186 621418 44422 621654
rect 44186 621098 44422 621334
rect 44186 585418 44422 585654
rect 44186 585098 44422 585334
rect 44186 549418 44422 549654
rect 44186 549098 44422 549334
rect 44186 513418 44422 513654
rect 44186 513098 44422 513334
rect 44186 477418 44422 477654
rect 44186 477098 44422 477334
rect 44186 441418 44422 441654
rect 44186 441098 44422 441334
rect 44186 405418 44422 405654
rect 44186 405098 44422 405334
rect 44186 369418 44422 369654
rect 44186 369098 44422 369334
rect 44186 333418 44422 333654
rect 44186 333098 44422 333334
rect 44186 297418 44422 297654
rect 44186 297098 44422 297334
rect 44186 261418 44422 261654
rect 44186 261098 44422 261334
rect 44186 225418 44422 225654
rect 44186 225098 44422 225334
rect 44186 189418 44422 189654
rect 44186 189098 44422 189334
rect 44186 153418 44422 153654
rect 44186 153098 44422 153334
rect 44186 117418 44422 117654
rect 44186 117098 44422 117334
rect 44186 81418 44422 81654
rect 44186 81098 44422 81334
rect 44186 45418 44422 45654
rect 44186 45098 44422 45334
rect 44186 9418 44422 9654
rect 44186 9098 44422 9334
rect 44186 -4262 44422 -4026
rect 44186 -4582 44422 -4346
rect 65786 711042 66022 711278
rect 65786 710722 66022 710958
rect 62186 709202 62422 709438
rect 62186 708882 62422 709118
rect 58586 707362 58822 707598
rect 58586 707042 58822 707278
rect 47786 697018 48022 697254
rect 47786 696698 48022 696934
rect 47786 661018 48022 661254
rect 47786 660698 48022 660934
rect 47786 625018 48022 625254
rect 47786 624698 48022 624934
rect 47786 589018 48022 589254
rect 47786 588698 48022 588934
rect 47786 553018 48022 553254
rect 47786 552698 48022 552934
rect 47786 517018 48022 517254
rect 47786 516698 48022 516934
rect 47786 481018 48022 481254
rect 47786 480698 48022 480934
rect 47786 445018 48022 445254
rect 47786 444698 48022 444934
rect 47786 409018 48022 409254
rect 47786 408698 48022 408934
rect 47786 373018 48022 373254
rect 47786 372698 48022 372934
rect 47786 337018 48022 337254
rect 47786 336698 48022 336934
rect 47786 301018 48022 301254
rect 47786 300698 48022 300934
rect 47786 265018 48022 265254
rect 47786 264698 48022 264934
rect 47786 229018 48022 229254
rect 47786 228698 48022 228934
rect 47786 193018 48022 193254
rect 47786 192698 48022 192934
rect 47786 157018 48022 157254
rect 47786 156698 48022 156934
rect 47786 121018 48022 121254
rect 47786 120698 48022 120934
rect 47786 85018 48022 85254
rect 47786 84698 48022 84934
rect 47786 49018 48022 49254
rect 47786 48698 48022 48934
rect 47786 13018 48022 13254
rect 47786 12698 48022 12934
rect 29786 -7022 30022 -6786
rect 29786 -7342 30022 -7106
rect 54986 705522 55222 705758
rect 54986 705202 55222 705438
rect 54986 668218 55222 668454
rect 54986 667898 55222 668134
rect 54986 632218 55222 632454
rect 54986 631898 55222 632134
rect 54986 596218 55222 596454
rect 54986 595898 55222 596134
rect 54986 560218 55222 560454
rect 54986 559898 55222 560134
rect 54986 524218 55222 524454
rect 54986 523898 55222 524134
rect 54986 488218 55222 488454
rect 54986 487898 55222 488134
rect 54986 452218 55222 452454
rect 54986 451898 55222 452134
rect 54986 416218 55222 416454
rect 54986 415898 55222 416134
rect 54986 380218 55222 380454
rect 54986 379898 55222 380134
rect 54986 344218 55222 344454
rect 54986 343898 55222 344134
rect 54986 308218 55222 308454
rect 54986 307898 55222 308134
rect 54986 272218 55222 272454
rect 54986 271898 55222 272134
rect 54986 236218 55222 236454
rect 54986 235898 55222 236134
rect 54986 200218 55222 200454
rect 54986 199898 55222 200134
rect 54986 164218 55222 164454
rect 54986 163898 55222 164134
rect 54986 128218 55222 128454
rect 54986 127898 55222 128134
rect 54986 92218 55222 92454
rect 54986 91898 55222 92134
rect 54986 56218 55222 56454
rect 54986 55898 55222 56134
rect 54986 20218 55222 20454
rect 54986 19898 55222 20134
rect 54986 -1502 55222 -1266
rect 54986 -1822 55222 -1586
rect 58586 671818 58822 672054
rect 58586 671498 58822 671734
rect 58586 635818 58822 636054
rect 58586 635498 58822 635734
rect 58586 599818 58822 600054
rect 58586 599498 58822 599734
rect 58586 563818 58822 564054
rect 58586 563498 58822 563734
rect 58586 527818 58822 528054
rect 58586 527498 58822 527734
rect 58586 491818 58822 492054
rect 58586 491498 58822 491734
rect 58586 455818 58822 456054
rect 58586 455498 58822 455734
rect 58586 419818 58822 420054
rect 58586 419498 58822 419734
rect 58586 383818 58822 384054
rect 58586 383498 58822 383734
rect 58586 347818 58822 348054
rect 58586 347498 58822 347734
rect 58586 311818 58822 312054
rect 58586 311498 58822 311734
rect 58586 275818 58822 276054
rect 58586 275498 58822 275734
rect 58586 239818 58822 240054
rect 58586 239498 58822 239734
rect 58586 203818 58822 204054
rect 58586 203498 58822 203734
rect 58586 167818 58822 168054
rect 58586 167498 58822 167734
rect 58586 131818 58822 132054
rect 58586 131498 58822 131734
rect 58586 95818 58822 96054
rect 58586 95498 58822 95734
rect 58586 59818 58822 60054
rect 58586 59498 58822 59734
rect 58586 23818 58822 24054
rect 58586 23498 58822 23734
rect 58586 -3342 58822 -3106
rect 58586 -3662 58822 -3426
rect 62186 675418 62422 675654
rect 62186 675098 62422 675334
rect 62186 639418 62422 639654
rect 62186 639098 62422 639334
rect 62186 603418 62422 603654
rect 62186 603098 62422 603334
rect 62186 567418 62422 567654
rect 62186 567098 62422 567334
rect 62186 531418 62422 531654
rect 62186 531098 62422 531334
rect 62186 495418 62422 495654
rect 62186 495098 62422 495334
rect 62186 459418 62422 459654
rect 62186 459098 62422 459334
rect 62186 423418 62422 423654
rect 62186 423098 62422 423334
rect 62186 387418 62422 387654
rect 62186 387098 62422 387334
rect 62186 351418 62422 351654
rect 62186 351098 62422 351334
rect 62186 315418 62422 315654
rect 62186 315098 62422 315334
rect 62186 279418 62422 279654
rect 62186 279098 62422 279334
rect 62186 243418 62422 243654
rect 62186 243098 62422 243334
rect 62186 207418 62422 207654
rect 62186 207098 62422 207334
rect 62186 171418 62422 171654
rect 62186 171098 62422 171334
rect 62186 135418 62422 135654
rect 62186 135098 62422 135334
rect 62186 99418 62422 99654
rect 62186 99098 62422 99334
rect 62186 63418 62422 63654
rect 62186 63098 62422 63334
rect 62186 27418 62422 27654
rect 62186 27098 62422 27334
rect 62186 -5182 62422 -4946
rect 62186 -5502 62422 -5266
rect 83786 710122 84022 710358
rect 83786 709802 84022 710038
rect 80186 708282 80422 708518
rect 80186 707962 80422 708198
rect 76586 706442 76822 706678
rect 76586 706122 76822 706358
rect 65786 679018 66022 679254
rect 65786 678698 66022 678934
rect 65786 643018 66022 643254
rect 65786 642698 66022 642934
rect 65786 607018 66022 607254
rect 65786 606698 66022 606934
rect 65786 571018 66022 571254
rect 65786 570698 66022 570934
rect 65786 535018 66022 535254
rect 65786 534698 66022 534934
rect 65786 499018 66022 499254
rect 65786 498698 66022 498934
rect 65786 463018 66022 463254
rect 65786 462698 66022 462934
rect 65786 427018 66022 427254
rect 65786 426698 66022 426934
rect 65786 391018 66022 391254
rect 65786 390698 66022 390934
rect 65786 355018 66022 355254
rect 65786 354698 66022 354934
rect 65786 319018 66022 319254
rect 65786 318698 66022 318934
rect 65786 283018 66022 283254
rect 65786 282698 66022 282934
rect 65786 247018 66022 247254
rect 65786 246698 66022 246934
rect 65786 211018 66022 211254
rect 65786 210698 66022 210934
rect 65786 175018 66022 175254
rect 65786 174698 66022 174934
rect 65786 139018 66022 139254
rect 65786 138698 66022 138934
rect 65786 103018 66022 103254
rect 65786 102698 66022 102934
rect 65786 67018 66022 67254
rect 65786 66698 66022 66934
rect 65786 31018 66022 31254
rect 65786 30698 66022 30934
rect 47786 -6102 48022 -5866
rect 47786 -6422 48022 -6186
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 72986 686218 73222 686454
rect 72986 685898 73222 686134
rect 72986 650218 73222 650454
rect 72986 649898 73222 650134
rect 72986 614218 73222 614454
rect 72986 613898 73222 614134
rect 72986 578218 73222 578454
rect 72986 577898 73222 578134
rect 72986 542218 73222 542454
rect 72986 541898 73222 542134
rect 72986 506218 73222 506454
rect 72986 505898 73222 506134
rect 72986 470218 73222 470454
rect 72986 469898 73222 470134
rect 72986 434218 73222 434454
rect 72986 433898 73222 434134
rect 72986 398218 73222 398454
rect 72986 397898 73222 398134
rect 72986 362218 73222 362454
rect 72986 361898 73222 362134
rect 72986 326218 73222 326454
rect 72986 325898 73222 326134
rect 72986 290218 73222 290454
rect 72986 289898 73222 290134
rect 72986 254218 73222 254454
rect 72986 253898 73222 254134
rect 72986 218218 73222 218454
rect 72986 217898 73222 218134
rect 72986 182218 73222 182454
rect 72986 181898 73222 182134
rect 72986 146218 73222 146454
rect 72986 145898 73222 146134
rect 72986 110218 73222 110454
rect 72986 109898 73222 110134
rect 72986 74218 73222 74454
rect 72986 73898 73222 74134
rect 72986 38218 73222 38454
rect 72986 37898 73222 38134
rect 72986 2218 73222 2454
rect 72986 1898 73222 2134
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 76586 689818 76822 690054
rect 76586 689498 76822 689734
rect 76586 653818 76822 654054
rect 76586 653498 76822 653734
rect 76586 617818 76822 618054
rect 76586 617498 76822 617734
rect 76586 581818 76822 582054
rect 76586 581498 76822 581734
rect 76586 545818 76822 546054
rect 76586 545498 76822 545734
rect 76586 509818 76822 510054
rect 76586 509498 76822 509734
rect 76586 473818 76822 474054
rect 76586 473498 76822 473734
rect 76586 437818 76822 438054
rect 76586 437498 76822 437734
rect 76586 401818 76822 402054
rect 76586 401498 76822 401734
rect 76586 365818 76822 366054
rect 76586 365498 76822 365734
rect 76586 329818 76822 330054
rect 76586 329498 76822 329734
rect 76586 293818 76822 294054
rect 76586 293498 76822 293734
rect 76586 257818 76822 258054
rect 76586 257498 76822 257734
rect 76586 221818 76822 222054
rect 76586 221498 76822 221734
rect 76586 185818 76822 186054
rect 76586 185498 76822 185734
rect 76586 149818 76822 150054
rect 76586 149498 76822 149734
rect 76586 113818 76822 114054
rect 76586 113498 76822 113734
rect 76586 77818 76822 78054
rect 76586 77498 76822 77734
rect 76586 41818 76822 42054
rect 76586 41498 76822 41734
rect 76586 5818 76822 6054
rect 76586 5498 76822 5734
rect 76586 -2422 76822 -2186
rect 76586 -2742 76822 -2506
rect 80186 693418 80422 693654
rect 80186 693098 80422 693334
rect 80186 657418 80422 657654
rect 80186 657098 80422 657334
rect 80186 621418 80422 621654
rect 80186 621098 80422 621334
rect 80186 585418 80422 585654
rect 80186 585098 80422 585334
rect 80186 549418 80422 549654
rect 80186 549098 80422 549334
rect 80186 513418 80422 513654
rect 80186 513098 80422 513334
rect 80186 477418 80422 477654
rect 80186 477098 80422 477334
rect 80186 441418 80422 441654
rect 80186 441098 80422 441334
rect 80186 405418 80422 405654
rect 80186 405098 80422 405334
rect 80186 369418 80422 369654
rect 80186 369098 80422 369334
rect 80186 333418 80422 333654
rect 80186 333098 80422 333334
rect 80186 297418 80422 297654
rect 80186 297098 80422 297334
rect 80186 261418 80422 261654
rect 80186 261098 80422 261334
rect 80186 225418 80422 225654
rect 80186 225098 80422 225334
rect 80186 189418 80422 189654
rect 80186 189098 80422 189334
rect 80186 153418 80422 153654
rect 80186 153098 80422 153334
rect 80186 117418 80422 117654
rect 80186 117098 80422 117334
rect 80186 81418 80422 81654
rect 80186 81098 80422 81334
rect 80186 45418 80422 45654
rect 80186 45098 80422 45334
rect 80186 9418 80422 9654
rect 80186 9098 80422 9334
rect 80186 -4262 80422 -4026
rect 80186 -4582 80422 -4346
rect 101786 711042 102022 711278
rect 101786 710722 102022 710958
rect 98186 709202 98422 709438
rect 98186 708882 98422 709118
rect 94586 707362 94822 707598
rect 94586 707042 94822 707278
rect 83786 697018 84022 697254
rect 83786 696698 84022 696934
rect 83786 661018 84022 661254
rect 83786 660698 84022 660934
rect 83786 625018 84022 625254
rect 83786 624698 84022 624934
rect 83786 589018 84022 589254
rect 83786 588698 84022 588934
rect 83786 553018 84022 553254
rect 83786 552698 84022 552934
rect 83786 517018 84022 517254
rect 83786 516698 84022 516934
rect 83786 481018 84022 481254
rect 83786 480698 84022 480934
rect 83786 445018 84022 445254
rect 83786 444698 84022 444934
rect 83786 409018 84022 409254
rect 83786 408698 84022 408934
rect 83786 373018 84022 373254
rect 83786 372698 84022 372934
rect 83786 337018 84022 337254
rect 83786 336698 84022 336934
rect 83786 301018 84022 301254
rect 83786 300698 84022 300934
rect 83786 265018 84022 265254
rect 83786 264698 84022 264934
rect 83786 229018 84022 229254
rect 83786 228698 84022 228934
rect 83786 193018 84022 193254
rect 83786 192698 84022 192934
rect 83786 157018 84022 157254
rect 83786 156698 84022 156934
rect 83786 121018 84022 121254
rect 83786 120698 84022 120934
rect 83786 85018 84022 85254
rect 83786 84698 84022 84934
rect 83786 49018 84022 49254
rect 83786 48698 84022 48934
rect 83786 13018 84022 13254
rect 83786 12698 84022 12934
rect 65786 -7022 66022 -6786
rect 65786 -7342 66022 -7106
rect 90986 705522 91222 705758
rect 90986 705202 91222 705438
rect 90986 668218 91222 668454
rect 90986 667898 91222 668134
rect 90986 632218 91222 632454
rect 90986 631898 91222 632134
rect 90986 596218 91222 596454
rect 90986 595898 91222 596134
rect 90986 560218 91222 560454
rect 90986 559898 91222 560134
rect 90986 524218 91222 524454
rect 90986 523898 91222 524134
rect 90986 488218 91222 488454
rect 90986 487898 91222 488134
rect 90986 452218 91222 452454
rect 90986 451898 91222 452134
rect 90986 416218 91222 416454
rect 90986 415898 91222 416134
rect 90986 380218 91222 380454
rect 90986 379898 91222 380134
rect 90986 344218 91222 344454
rect 90986 343898 91222 344134
rect 90986 308218 91222 308454
rect 90986 307898 91222 308134
rect 90986 272218 91222 272454
rect 90986 271898 91222 272134
rect 90986 236218 91222 236454
rect 90986 235898 91222 236134
rect 90986 200218 91222 200454
rect 90986 199898 91222 200134
rect 90986 164218 91222 164454
rect 90986 163898 91222 164134
rect 90986 128218 91222 128454
rect 90986 127898 91222 128134
rect 90986 92218 91222 92454
rect 90986 91898 91222 92134
rect 90986 56218 91222 56454
rect 90986 55898 91222 56134
rect 90986 20218 91222 20454
rect 90986 19898 91222 20134
rect 90986 -1502 91222 -1266
rect 90986 -1822 91222 -1586
rect 94586 671818 94822 672054
rect 94586 671498 94822 671734
rect 94586 635818 94822 636054
rect 94586 635498 94822 635734
rect 94586 599818 94822 600054
rect 94586 599498 94822 599734
rect 94586 563818 94822 564054
rect 94586 563498 94822 563734
rect 94586 527818 94822 528054
rect 94586 527498 94822 527734
rect 94586 491818 94822 492054
rect 94586 491498 94822 491734
rect 94586 455818 94822 456054
rect 94586 455498 94822 455734
rect 94586 419818 94822 420054
rect 94586 419498 94822 419734
rect 94586 383818 94822 384054
rect 94586 383498 94822 383734
rect 94586 347818 94822 348054
rect 94586 347498 94822 347734
rect 94586 311818 94822 312054
rect 94586 311498 94822 311734
rect 94586 275818 94822 276054
rect 94586 275498 94822 275734
rect 94586 239818 94822 240054
rect 94586 239498 94822 239734
rect 94586 203818 94822 204054
rect 94586 203498 94822 203734
rect 94586 167818 94822 168054
rect 94586 167498 94822 167734
rect 94586 131818 94822 132054
rect 94586 131498 94822 131734
rect 94586 95818 94822 96054
rect 94586 95498 94822 95734
rect 94586 59818 94822 60054
rect 94586 59498 94822 59734
rect 94586 23818 94822 24054
rect 94586 23498 94822 23734
rect 94586 -3342 94822 -3106
rect 94586 -3662 94822 -3426
rect 98186 675418 98422 675654
rect 98186 675098 98422 675334
rect 98186 639418 98422 639654
rect 98186 639098 98422 639334
rect 98186 603418 98422 603654
rect 98186 603098 98422 603334
rect 98186 567418 98422 567654
rect 98186 567098 98422 567334
rect 98186 531418 98422 531654
rect 98186 531098 98422 531334
rect 98186 495418 98422 495654
rect 98186 495098 98422 495334
rect 98186 459418 98422 459654
rect 98186 459098 98422 459334
rect 98186 423418 98422 423654
rect 98186 423098 98422 423334
rect 98186 387418 98422 387654
rect 98186 387098 98422 387334
rect 98186 351418 98422 351654
rect 98186 351098 98422 351334
rect 98186 315418 98422 315654
rect 98186 315098 98422 315334
rect 98186 279418 98422 279654
rect 98186 279098 98422 279334
rect 98186 243418 98422 243654
rect 98186 243098 98422 243334
rect 98186 207418 98422 207654
rect 98186 207098 98422 207334
rect 98186 171418 98422 171654
rect 98186 171098 98422 171334
rect 98186 135418 98422 135654
rect 98186 135098 98422 135334
rect 98186 99418 98422 99654
rect 98186 99098 98422 99334
rect 98186 63418 98422 63654
rect 98186 63098 98422 63334
rect 98186 27418 98422 27654
rect 98186 27098 98422 27334
rect 98186 -5182 98422 -4946
rect 98186 -5502 98422 -5266
rect 119786 710122 120022 710358
rect 119786 709802 120022 710038
rect 116186 708282 116422 708518
rect 116186 707962 116422 708198
rect 112586 706442 112822 706678
rect 112586 706122 112822 706358
rect 101786 679018 102022 679254
rect 101786 678698 102022 678934
rect 101786 643018 102022 643254
rect 101786 642698 102022 642934
rect 101786 607018 102022 607254
rect 101786 606698 102022 606934
rect 101786 571018 102022 571254
rect 101786 570698 102022 570934
rect 101786 535018 102022 535254
rect 101786 534698 102022 534934
rect 101786 499018 102022 499254
rect 101786 498698 102022 498934
rect 101786 463018 102022 463254
rect 101786 462698 102022 462934
rect 101786 427018 102022 427254
rect 101786 426698 102022 426934
rect 101786 391018 102022 391254
rect 101786 390698 102022 390934
rect 101786 355018 102022 355254
rect 101786 354698 102022 354934
rect 101786 319018 102022 319254
rect 101786 318698 102022 318934
rect 101786 283018 102022 283254
rect 101786 282698 102022 282934
rect 101786 247018 102022 247254
rect 101786 246698 102022 246934
rect 101786 211018 102022 211254
rect 101786 210698 102022 210934
rect 101786 175018 102022 175254
rect 101786 174698 102022 174934
rect 101786 139018 102022 139254
rect 101786 138698 102022 138934
rect 101786 103018 102022 103254
rect 101786 102698 102022 102934
rect 101786 67018 102022 67254
rect 101786 66698 102022 66934
rect 101786 31018 102022 31254
rect 101786 30698 102022 30934
rect 83786 -6102 84022 -5866
rect 83786 -6422 84022 -6186
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 108986 686218 109222 686454
rect 108986 685898 109222 686134
rect 108986 650218 109222 650454
rect 108986 649898 109222 650134
rect 108986 614218 109222 614454
rect 108986 613898 109222 614134
rect 108986 578218 109222 578454
rect 108986 577898 109222 578134
rect 108986 542218 109222 542454
rect 108986 541898 109222 542134
rect 108986 506218 109222 506454
rect 108986 505898 109222 506134
rect 108986 470218 109222 470454
rect 108986 469898 109222 470134
rect 108986 434218 109222 434454
rect 108986 433898 109222 434134
rect 108986 398218 109222 398454
rect 108986 397898 109222 398134
rect 108986 362218 109222 362454
rect 108986 361898 109222 362134
rect 108986 326218 109222 326454
rect 108986 325898 109222 326134
rect 108986 290218 109222 290454
rect 108986 289898 109222 290134
rect 108986 254218 109222 254454
rect 108986 253898 109222 254134
rect 108986 218218 109222 218454
rect 108986 217898 109222 218134
rect 108986 182218 109222 182454
rect 108986 181898 109222 182134
rect 108986 146218 109222 146454
rect 108986 145898 109222 146134
rect 108986 110218 109222 110454
rect 108986 109898 109222 110134
rect 108986 74218 109222 74454
rect 108986 73898 109222 74134
rect 108986 38218 109222 38454
rect 108986 37898 109222 38134
rect 108986 2218 109222 2454
rect 108986 1898 109222 2134
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 112586 689818 112822 690054
rect 112586 689498 112822 689734
rect 112586 653818 112822 654054
rect 112586 653498 112822 653734
rect 112586 617818 112822 618054
rect 112586 617498 112822 617734
rect 112586 581818 112822 582054
rect 112586 581498 112822 581734
rect 112586 545818 112822 546054
rect 112586 545498 112822 545734
rect 112586 509818 112822 510054
rect 112586 509498 112822 509734
rect 112586 473818 112822 474054
rect 112586 473498 112822 473734
rect 112586 437818 112822 438054
rect 112586 437498 112822 437734
rect 112586 401818 112822 402054
rect 112586 401498 112822 401734
rect 112586 365818 112822 366054
rect 112586 365498 112822 365734
rect 112586 329818 112822 330054
rect 112586 329498 112822 329734
rect 112586 293818 112822 294054
rect 112586 293498 112822 293734
rect 112586 257818 112822 258054
rect 112586 257498 112822 257734
rect 112586 221818 112822 222054
rect 112586 221498 112822 221734
rect 112586 185818 112822 186054
rect 112586 185498 112822 185734
rect 112586 149818 112822 150054
rect 112586 149498 112822 149734
rect 112586 113818 112822 114054
rect 112586 113498 112822 113734
rect 112586 77818 112822 78054
rect 112586 77498 112822 77734
rect 112586 41818 112822 42054
rect 112586 41498 112822 41734
rect 112586 5818 112822 6054
rect 112586 5498 112822 5734
rect 112586 -2422 112822 -2186
rect 112586 -2742 112822 -2506
rect 116186 693418 116422 693654
rect 116186 693098 116422 693334
rect 116186 657418 116422 657654
rect 116186 657098 116422 657334
rect 116186 621418 116422 621654
rect 116186 621098 116422 621334
rect 116186 585418 116422 585654
rect 116186 585098 116422 585334
rect 116186 549418 116422 549654
rect 116186 549098 116422 549334
rect 116186 513418 116422 513654
rect 116186 513098 116422 513334
rect 116186 477418 116422 477654
rect 116186 477098 116422 477334
rect 116186 441418 116422 441654
rect 116186 441098 116422 441334
rect 116186 405418 116422 405654
rect 116186 405098 116422 405334
rect 116186 369418 116422 369654
rect 116186 369098 116422 369334
rect 116186 333418 116422 333654
rect 116186 333098 116422 333334
rect 116186 297418 116422 297654
rect 116186 297098 116422 297334
rect 116186 261418 116422 261654
rect 116186 261098 116422 261334
rect 116186 225418 116422 225654
rect 116186 225098 116422 225334
rect 116186 189418 116422 189654
rect 116186 189098 116422 189334
rect 116186 153418 116422 153654
rect 116186 153098 116422 153334
rect 116186 117418 116422 117654
rect 116186 117098 116422 117334
rect 116186 81418 116422 81654
rect 116186 81098 116422 81334
rect 116186 45418 116422 45654
rect 116186 45098 116422 45334
rect 116186 9418 116422 9654
rect 116186 9098 116422 9334
rect 116186 -4262 116422 -4026
rect 116186 -4582 116422 -4346
rect 137786 711042 138022 711278
rect 137786 710722 138022 710958
rect 134186 709202 134422 709438
rect 134186 708882 134422 709118
rect 130586 707362 130822 707598
rect 130586 707042 130822 707278
rect 119786 697018 120022 697254
rect 119786 696698 120022 696934
rect 119786 661018 120022 661254
rect 119786 660698 120022 660934
rect 119786 625018 120022 625254
rect 119786 624698 120022 624934
rect 119786 589018 120022 589254
rect 119786 588698 120022 588934
rect 119786 553018 120022 553254
rect 119786 552698 120022 552934
rect 119786 517018 120022 517254
rect 119786 516698 120022 516934
rect 119786 481018 120022 481254
rect 119786 480698 120022 480934
rect 119786 445018 120022 445254
rect 119786 444698 120022 444934
rect 119786 409018 120022 409254
rect 119786 408698 120022 408934
rect 119786 373018 120022 373254
rect 119786 372698 120022 372934
rect 119786 337018 120022 337254
rect 119786 336698 120022 336934
rect 119786 301018 120022 301254
rect 119786 300698 120022 300934
rect 119786 265018 120022 265254
rect 119786 264698 120022 264934
rect 119786 229018 120022 229254
rect 119786 228698 120022 228934
rect 119786 193018 120022 193254
rect 119786 192698 120022 192934
rect 119786 157018 120022 157254
rect 119786 156698 120022 156934
rect 119786 121018 120022 121254
rect 119786 120698 120022 120934
rect 119786 85018 120022 85254
rect 119786 84698 120022 84934
rect 119786 49018 120022 49254
rect 119786 48698 120022 48934
rect 119786 13018 120022 13254
rect 119786 12698 120022 12934
rect 101786 -7022 102022 -6786
rect 101786 -7342 102022 -7106
rect 126986 705522 127222 705758
rect 126986 705202 127222 705438
rect 126986 668218 127222 668454
rect 126986 667898 127222 668134
rect 126986 632218 127222 632454
rect 126986 631898 127222 632134
rect 126986 596218 127222 596454
rect 126986 595898 127222 596134
rect 126986 560218 127222 560454
rect 126986 559898 127222 560134
rect 126986 524218 127222 524454
rect 126986 523898 127222 524134
rect 126986 488218 127222 488454
rect 126986 487898 127222 488134
rect 126986 452218 127222 452454
rect 126986 451898 127222 452134
rect 126986 416218 127222 416454
rect 126986 415898 127222 416134
rect 126986 380218 127222 380454
rect 126986 379898 127222 380134
rect 126986 344218 127222 344454
rect 126986 343898 127222 344134
rect 126986 308218 127222 308454
rect 126986 307898 127222 308134
rect 126986 272218 127222 272454
rect 126986 271898 127222 272134
rect 126986 236218 127222 236454
rect 126986 235898 127222 236134
rect 126986 200218 127222 200454
rect 126986 199898 127222 200134
rect 126986 164218 127222 164454
rect 126986 163898 127222 164134
rect 126986 128218 127222 128454
rect 126986 127898 127222 128134
rect 126986 92218 127222 92454
rect 126986 91898 127222 92134
rect 126986 56218 127222 56454
rect 126986 55898 127222 56134
rect 126986 20218 127222 20454
rect 126986 19898 127222 20134
rect 126986 -1502 127222 -1266
rect 126986 -1822 127222 -1586
rect 130586 671818 130822 672054
rect 130586 671498 130822 671734
rect 130586 635818 130822 636054
rect 130586 635498 130822 635734
rect 130586 599818 130822 600054
rect 130586 599498 130822 599734
rect 130586 563818 130822 564054
rect 130586 563498 130822 563734
rect 130586 527818 130822 528054
rect 130586 527498 130822 527734
rect 130586 491818 130822 492054
rect 130586 491498 130822 491734
rect 130586 455818 130822 456054
rect 130586 455498 130822 455734
rect 130586 419818 130822 420054
rect 130586 419498 130822 419734
rect 130586 383818 130822 384054
rect 130586 383498 130822 383734
rect 130586 347818 130822 348054
rect 130586 347498 130822 347734
rect 130586 311818 130822 312054
rect 130586 311498 130822 311734
rect 130586 275818 130822 276054
rect 130586 275498 130822 275734
rect 130586 239818 130822 240054
rect 130586 239498 130822 239734
rect 130586 203818 130822 204054
rect 130586 203498 130822 203734
rect 130586 167818 130822 168054
rect 130586 167498 130822 167734
rect 130586 131818 130822 132054
rect 130586 131498 130822 131734
rect 130586 95818 130822 96054
rect 130586 95498 130822 95734
rect 130586 59818 130822 60054
rect 130586 59498 130822 59734
rect 130586 23818 130822 24054
rect 130586 23498 130822 23734
rect 130586 -3342 130822 -3106
rect 130586 -3662 130822 -3426
rect 134186 675418 134422 675654
rect 134186 675098 134422 675334
rect 134186 639418 134422 639654
rect 134186 639098 134422 639334
rect 134186 603418 134422 603654
rect 134186 603098 134422 603334
rect 134186 567418 134422 567654
rect 134186 567098 134422 567334
rect 134186 531418 134422 531654
rect 134186 531098 134422 531334
rect 134186 495418 134422 495654
rect 134186 495098 134422 495334
rect 134186 459418 134422 459654
rect 134186 459098 134422 459334
rect 134186 423418 134422 423654
rect 134186 423098 134422 423334
rect 134186 387418 134422 387654
rect 134186 387098 134422 387334
rect 134186 351418 134422 351654
rect 134186 351098 134422 351334
rect 134186 315418 134422 315654
rect 134186 315098 134422 315334
rect 134186 279418 134422 279654
rect 134186 279098 134422 279334
rect 134186 243418 134422 243654
rect 134186 243098 134422 243334
rect 134186 207418 134422 207654
rect 134186 207098 134422 207334
rect 134186 171418 134422 171654
rect 134186 171098 134422 171334
rect 134186 135418 134422 135654
rect 134186 135098 134422 135334
rect 134186 99418 134422 99654
rect 134186 99098 134422 99334
rect 134186 63418 134422 63654
rect 134186 63098 134422 63334
rect 134186 27418 134422 27654
rect 134186 27098 134422 27334
rect 134186 -5182 134422 -4946
rect 134186 -5502 134422 -5266
rect 155786 710122 156022 710358
rect 155786 709802 156022 710038
rect 152186 708282 152422 708518
rect 152186 707962 152422 708198
rect 148586 706442 148822 706678
rect 148586 706122 148822 706358
rect 137786 679018 138022 679254
rect 137786 678698 138022 678934
rect 137786 643018 138022 643254
rect 137786 642698 138022 642934
rect 137786 607018 138022 607254
rect 137786 606698 138022 606934
rect 137786 571018 138022 571254
rect 137786 570698 138022 570934
rect 137786 535018 138022 535254
rect 137786 534698 138022 534934
rect 137786 499018 138022 499254
rect 137786 498698 138022 498934
rect 137786 463018 138022 463254
rect 137786 462698 138022 462934
rect 137786 427018 138022 427254
rect 137786 426698 138022 426934
rect 137786 391018 138022 391254
rect 137786 390698 138022 390934
rect 137786 355018 138022 355254
rect 137786 354698 138022 354934
rect 137786 319018 138022 319254
rect 137786 318698 138022 318934
rect 137786 283018 138022 283254
rect 137786 282698 138022 282934
rect 137786 247018 138022 247254
rect 137786 246698 138022 246934
rect 137786 211018 138022 211254
rect 137786 210698 138022 210934
rect 137786 175018 138022 175254
rect 137786 174698 138022 174934
rect 137786 139018 138022 139254
rect 137786 138698 138022 138934
rect 137786 103018 138022 103254
rect 137786 102698 138022 102934
rect 137786 67018 138022 67254
rect 137786 66698 138022 66934
rect 137786 31018 138022 31254
rect 137786 30698 138022 30934
rect 119786 -6102 120022 -5866
rect 119786 -6422 120022 -6186
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 144986 686218 145222 686454
rect 144986 685898 145222 686134
rect 144986 650218 145222 650454
rect 144986 649898 145222 650134
rect 144986 614218 145222 614454
rect 144986 613898 145222 614134
rect 144986 578218 145222 578454
rect 144986 577898 145222 578134
rect 144986 542218 145222 542454
rect 144986 541898 145222 542134
rect 144986 506218 145222 506454
rect 144986 505898 145222 506134
rect 144986 470218 145222 470454
rect 144986 469898 145222 470134
rect 144986 434218 145222 434454
rect 144986 433898 145222 434134
rect 144986 398218 145222 398454
rect 144986 397898 145222 398134
rect 144986 362218 145222 362454
rect 144986 361898 145222 362134
rect 144986 326218 145222 326454
rect 144986 325898 145222 326134
rect 144986 290218 145222 290454
rect 144986 289898 145222 290134
rect 144986 254218 145222 254454
rect 144986 253898 145222 254134
rect 144986 218218 145222 218454
rect 144986 217898 145222 218134
rect 144986 182218 145222 182454
rect 144986 181898 145222 182134
rect 144986 146218 145222 146454
rect 144986 145898 145222 146134
rect 144986 110218 145222 110454
rect 144986 109898 145222 110134
rect 144986 74218 145222 74454
rect 144986 73898 145222 74134
rect 144986 38218 145222 38454
rect 144986 37898 145222 38134
rect 144986 2218 145222 2454
rect 144986 1898 145222 2134
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 148586 689818 148822 690054
rect 148586 689498 148822 689734
rect 148586 653818 148822 654054
rect 148586 653498 148822 653734
rect 148586 617818 148822 618054
rect 148586 617498 148822 617734
rect 148586 581818 148822 582054
rect 148586 581498 148822 581734
rect 148586 545818 148822 546054
rect 148586 545498 148822 545734
rect 148586 509818 148822 510054
rect 148586 509498 148822 509734
rect 148586 473818 148822 474054
rect 148586 473498 148822 473734
rect 148586 437818 148822 438054
rect 148586 437498 148822 437734
rect 148586 401818 148822 402054
rect 148586 401498 148822 401734
rect 148586 365818 148822 366054
rect 148586 365498 148822 365734
rect 148586 329818 148822 330054
rect 148586 329498 148822 329734
rect 148586 293818 148822 294054
rect 148586 293498 148822 293734
rect 148586 257818 148822 258054
rect 148586 257498 148822 257734
rect 148586 221818 148822 222054
rect 148586 221498 148822 221734
rect 148586 185818 148822 186054
rect 148586 185498 148822 185734
rect 148586 149818 148822 150054
rect 148586 149498 148822 149734
rect 148586 113818 148822 114054
rect 148586 113498 148822 113734
rect 148586 77818 148822 78054
rect 148586 77498 148822 77734
rect 148586 41818 148822 42054
rect 148586 41498 148822 41734
rect 148586 5818 148822 6054
rect 148586 5498 148822 5734
rect 148586 -2422 148822 -2186
rect 148586 -2742 148822 -2506
rect 152186 693418 152422 693654
rect 152186 693098 152422 693334
rect 152186 657418 152422 657654
rect 152186 657098 152422 657334
rect 152186 621418 152422 621654
rect 152186 621098 152422 621334
rect 152186 585418 152422 585654
rect 152186 585098 152422 585334
rect 152186 549418 152422 549654
rect 152186 549098 152422 549334
rect 152186 513418 152422 513654
rect 152186 513098 152422 513334
rect 152186 477418 152422 477654
rect 152186 477098 152422 477334
rect 152186 441418 152422 441654
rect 152186 441098 152422 441334
rect 152186 405418 152422 405654
rect 152186 405098 152422 405334
rect 152186 369418 152422 369654
rect 152186 369098 152422 369334
rect 152186 333418 152422 333654
rect 152186 333098 152422 333334
rect 152186 297418 152422 297654
rect 152186 297098 152422 297334
rect 152186 261418 152422 261654
rect 152186 261098 152422 261334
rect 152186 225418 152422 225654
rect 152186 225098 152422 225334
rect 152186 189418 152422 189654
rect 152186 189098 152422 189334
rect 152186 153418 152422 153654
rect 152186 153098 152422 153334
rect 152186 117418 152422 117654
rect 152186 117098 152422 117334
rect 152186 81418 152422 81654
rect 152186 81098 152422 81334
rect 152186 45418 152422 45654
rect 152186 45098 152422 45334
rect 152186 9418 152422 9654
rect 152186 9098 152422 9334
rect 152186 -4262 152422 -4026
rect 152186 -4582 152422 -4346
rect 173786 711042 174022 711278
rect 173786 710722 174022 710958
rect 170186 709202 170422 709438
rect 170186 708882 170422 709118
rect 166586 707362 166822 707598
rect 166586 707042 166822 707278
rect 155786 697018 156022 697254
rect 155786 696698 156022 696934
rect 155786 661018 156022 661254
rect 155786 660698 156022 660934
rect 155786 625018 156022 625254
rect 155786 624698 156022 624934
rect 155786 589018 156022 589254
rect 155786 588698 156022 588934
rect 155786 553018 156022 553254
rect 155786 552698 156022 552934
rect 155786 517018 156022 517254
rect 155786 516698 156022 516934
rect 155786 481018 156022 481254
rect 155786 480698 156022 480934
rect 155786 445018 156022 445254
rect 155786 444698 156022 444934
rect 155786 409018 156022 409254
rect 155786 408698 156022 408934
rect 155786 373018 156022 373254
rect 155786 372698 156022 372934
rect 155786 337018 156022 337254
rect 155786 336698 156022 336934
rect 155786 301018 156022 301254
rect 155786 300698 156022 300934
rect 155786 265018 156022 265254
rect 155786 264698 156022 264934
rect 155786 229018 156022 229254
rect 155786 228698 156022 228934
rect 155786 193018 156022 193254
rect 155786 192698 156022 192934
rect 155786 157018 156022 157254
rect 155786 156698 156022 156934
rect 155786 121018 156022 121254
rect 155786 120698 156022 120934
rect 155786 85018 156022 85254
rect 155786 84698 156022 84934
rect 155786 49018 156022 49254
rect 155786 48698 156022 48934
rect 155786 13018 156022 13254
rect 155786 12698 156022 12934
rect 137786 -7022 138022 -6786
rect 137786 -7342 138022 -7106
rect 162986 705522 163222 705758
rect 162986 705202 163222 705438
rect 162986 668218 163222 668454
rect 162986 667898 163222 668134
rect 162986 632218 163222 632454
rect 162986 631898 163222 632134
rect 162986 596218 163222 596454
rect 162986 595898 163222 596134
rect 162986 560218 163222 560454
rect 162986 559898 163222 560134
rect 162986 524218 163222 524454
rect 162986 523898 163222 524134
rect 162986 488218 163222 488454
rect 162986 487898 163222 488134
rect 162986 452218 163222 452454
rect 162986 451898 163222 452134
rect 162986 416218 163222 416454
rect 162986 415898 163222 416134
rect 162986 380218 163222 380454
rect 162986 379898 163222 380134
rect 162986 344218 163222 344454
rect 162986 343898 163222 344134
rect 162986 308218 163222 308454
rect 162986 307898 163222 308134
rect 162986 272218 163222 272454
rect 162986 271898 163222 272134
rect 162986 236218 163222 236454
rect 162986 235898 163222 236134
rect 162986 200218 163222 200454
rect 162986 199898 163222 200134
rect 162986 164218 163222 164454
rect 162986 163898 163222 164134
rect 162986 128218 163222 128454
rect 162986 127898 163222 128134
rect 162986 92218 163222 92454
rect 162986 91898 163222 92134
rect 162986 56218 163222 56454
rect 162986 55898 163222 56134
rect 162986 20218 163222 20454
rect 162986 19898 163222 20134
rect 162986 -1502 163222 -1266
rect 162986 -1822 163222 -1586
rect 166586 671818 166822 672054
rect 166586 671498 166822 671734
rect 166586 635818 166822 636054
rect 166586 635498 166822 635734
rect 166586 599818 166822 600054
rect 166586 599498 166822 599734
rect 166586 563818 166822 564054
rect 166586 563498 166822 563734
rect 166586 527818 166822 528054
rect 166586 527498 166822 527734
rect 166586 491818 166822 492054
rect 166586 491498 166822 491734
rect 166586 455818 166822 456054
rect 166586 455498 166822 455734
rect 166586 419818 166822 420054
rect 166586 419498 166822 419734
rect 166586 383818 166822 384054
rect 166586 383498 166822 383734
rect 166586 347818 166822 348054
rect 166586 347498 166822 347734
rect 166586 311818 166822 312054
rect 166586 311498 166822 311734
rect 166586 275818 166822 276054
rect 166586 275498 166822 275734
rect 166586 239818 166822 240054
rect 166586 239498 166822 239734
rect 166586 203818 166822 204054
rect 166586 203498 166822 203734
rect 166586 167818 166822 168054
rect 166586 167498 166822 167734
rect 166586 131818 166822 132054
rect 166586 131498 166822 131734
rect 166586 95818 166822 96054
rect 166586 95498 166822 95734
rect 166586 59818 166822 60054
rect 166586 59498 166822 59734
rect 166586 23818 166822 24054
rect 166586 23498 166822 23734
rect 166586 -3342 166822 -3106
rect 166586 -3662 166822 -3426
rect 170186 675418 170422 675654
rect 170186 675098 170422 675334
rect 170186 639418 170422 639654
rect 170186 639098 170422 639334
rect 170186 603418 170422 603654
rect 170186 603098 170422 603334
rect 170186 567418 170422 567654
rect 170186 567098 170422 567334
rect 170186 531418 170422 531654
rect 170186 531098 170422 531334
rect 191786 710122 192022 710358
rect 191786 709802 192022 710038
rect 188186 708282 188422 708518
rect 188186 707962 188422 708198
rect 184586 706442 184822 706678
rect 184586 706122 184822 706358
rect 173786 679018 174022 679254
rect 173786 678698 174022 678934
rect 173786 643018 174022 643254
rect 173786 642698 174022 642934
rect 173786 607018 174022 607254
rect 173786 606698 174022 606934
rect 173786 571018 174022 571254
rect 173786 570698 174022 570934
rect 173786 535018 174022 535254
rect 173786 534698 174022 534934
rect 170186 495418 170422 495654
rect 170186 495098 170422 495334
rect 170186 459418 170422 459654
rect 170186 459098 170422 459334
rect 170186 423418 170422 423654
rect 170186 423098 170422 423334
rect 170186 387418 170422 387654
rect 170186 387098 170422 387334
rect 170186 351418 170422 351654
rect 170186 351098 170422 351334
rect 170186 315418 170422 315654
rect 170186 315098 170422 315334
rect 170186 279418 170422 279654
rect 170186 279098 170422 279334
rect 170186 243418 170422 243654
rect 170186 243098 170422 243334
rect 170186 207418 170422 207654
rect 170186 207098 170422 207334
rect 170186 171418 170422 171654
rect 170186 171098 170422 171334
rect 170186 135418 170422 135654
rect 170186 135098 170422 135334
rect 170186 99418 170422 99654
rect 170186 99098 170422 99334
rect 170186 63418 170422 63654
rect 170186 63098 170422 63334
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 180986 686218 181222 686454
rect 180986 685898 181222 686134
rect 180986 650218 181222 650454
rect 180986 649898 181222 650134
rect 180986 614218 181222 614454
rect 180986 613898 181222 614134
rect 180986 578218 181222 578454
rect 180986 577898 181222 578134
rect 180986 542218 181222 542454
rect 180986 541898 181222 542134
rect 173786 499018 174022 499254
rect 173786 498698 174022 498934
rect 173786 463018 174022 463254
rect 173786 462698 174022 462934
rect 173786 427018 174022 427254
rect 173786 426698 174022 426934
rect 173786 391018 174022 391254
rect 173786 390698 174022 390934
rect 173786 355018 174022 355254
rect 173786 354698 174022 354934
rect 173786 319018 174022 319254
rect 173786 318698 174022 318934
rect 173786 283018 174022 283254
rect 173786 282698 174022 282934
rect 173786 247018 174022 247254
rect 173786 246698 174022 246934
rect 173786 211018 174022 211254
rect 173786 210698 174022 210934
rect 173786 175018 174022 175254
rect 173786 174698 174022 174934
rect 173786 139018 174022 139254
rect 173786 138698 174022 138934
rect 173786 103018 174022 103254
rect 173786 102698 174022 102934
rect 173786 67018 174022 67254
rect 173786 66698 174022 66934
rect 170186 27418 170422 27654
rect 170186 27098 170422 27334
rect 170186 -5182 170422 -4946
rect 170186 -5502 170422 -5266
rect 173786 31018 174022 31254
rect 173786 30698 174022 30934
rect 155786 -6102 156022 -5866
rect 155786 -6422 156022 -6186
rect 184586 689818 184822 690054
rect 184586 689498 184822 689734
rect 184586 653818 184822 654054
rect 184586 653498 184822 653734
rect 184586 617818 184822 618054
rect 184586 617498 184822 617734
rect 184586 581818 184822 582054
rect 184586 581498 184822 581734
rect 184586 545818 184822 546054
rect 184586 545498 184822 545734
rect 180986 506218 181222 506454
rect 180986 505898 181222 506134
rect 180986 470218 181222 470454
rect 180986 469898 181222 470134
rect 180986 434218 181222 434454
rect 180986 433898 181222 434134
rect 180986 398218 181222 398454
rect 180986 397898 181222 398134
rect 180986 362218 181222 362454
rect 180986 361898 181222 362134
rect 180986 326218 181222 326454
rect 180986 325898 181222 326134
rect 180986 290218 181222 290454
rect 180986 289898 181222 290134
rect 180986 254218 181222 254454
rect 180986 253898 181222 254134
rect 180986 218218 181222 218454
rect 180986 217898 181222 218134
rect 180986 182218 181222 182454
rect 180986 181898 181222 182134
rect 180986 146218 181222 146454
rect 180986 145898 181222 146134
rect 180986 110218 181222 110454
rect 180986 109898 181222 110134
rect 180986 74218 181222 74454
rect 180986 73898 181222 74134
rect 180986 38218 181222 38454
rect 180986 37898 181222 38134
rect 180986 2218 181222 2454
rect 180986 1898 181222 2134
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 184586 509818 184822 510054
rect 184586 509498 184822 509734
rect 184586 473818 184822 474054
rect 184586 473498 184822 473734
rect 184586 437818 184822 438054
rect 184586 437498 184822 437734
rect 184586 401818 184822 402054
rect 184586 401498 184822 401734
rect 184586 365818 184822 366054
rect 184586 365498 184822 365734
rect 184586 329818 184822 330054
rect 184586 329498 184822 329734
rect 184586 293818 184822 294054
rect 184586 293498 184822 293734
rect 184586 257818 184822 258054
rect 184586 257498 184822 257734
rect 184586 221818 184822 222054
rect 184586 221498 184822 221734
rect 184586 185818 184822 186054
rect 184586 185498 184822 185734
rect 184586 149818 184822 150054
rect 184586 149498 184822 149734
rect 184586 113818 184822 114054
rect 184586 113498 184822 113734
rect 184586 77818 184822 78054
rect 184586 77498 184822 77734
rect 184586 41818 184822 42054
rect 184586 41498 184822 41734
rect 184586 5818 184822 6054
rect 184586 5498 184822 5734
rect 184586 -2422 184822 -2186
rect 184586 -2742 184822 -2506
rect 188186 693418 188422 693654
rect 188186 693098 188422 693334
rect 188186 657418 188422 657654
rect 188186 657098 188422 657334
rect 188186 621418 188422 621654
rect 188186 621098 188422 621334
rect 188186 585418 188422 585654
rect 188186 585098 188422 585334
rect 188186 549418 188422 549654
rect 188186 549098 188422 549334
rect 188186 513418 188422 513654
rect 188186 513098 188422 513334
rect 188186 477418 188422 477654
rect 188186 477098 188422 477334
rect 188186 441418 188422 441654
rect 188186 441098 188422 441334
rect 188186 405418 188422 405654
rect 188186 405098 188422 405334
rect 188186 369418 188422 369654
rect 188186 369098 188422 369334
rect 188186 333418 188422 333654
rect 188186 333098 188422 333334
rect 188186 297418 188422 297654
rect 188186 297098 188422 297334
rect 188186 261418 188422 261654
rect 188186 261098 188422 261334
rect 188186 225418 188422 225654
rect 188186 225098 188422 225334
rect 188186 189418 188422 189654
rect 188186 189098 188422 189334
rect 188186 153418 188422 153654
rect 188186 153098 188422 153334
rect 188186 117418 188422 117654
rect 188186 117098 188422 117334
rect 188186 81418 188422 81654
rect 188186 81098 188422 81334
rect 188186 45418 188422 45654
rect 188186 45098 188422 45334
rect 188186 9418 188422 9654
rect 188186 9098 188422 9334
rect 188186 -4262 188422 -4026
rect 188186 -4582 188422 -4346
rect 209786 711042 210022 711278
rect 209786 710722 210022 710958
rect 206186 709202 206422 709438
rect 206186 708882 206422 709118
rect 202586 707362 202822 707598
rect 202586 707042 202822 707278
rect 191786 697018 192022 697254
rect 191786 696698 192022 696934
rect 191786 661018 192022 661254
rect 191786 660698 192022 660934
rect 191786 625018 192022 625254
rect 191786 624698 192022 624934
rect 191786 589018 192022 589254
rect 191786 588698 192022 588934
rect 191786 553018 192022 553254
rect 191786 552698 192022 552934
rect 198986 705522 199222 705758
rect 198986 705202 199222 705438
rect 198986 668218 199222 668454
rect 198986 667898 199222 668134
rect 198986 632218 199222 632454
rect 198986 631898 199222 632134
rect 198986 596218 199222 596454
rect 198986 595898 199222 596134
rect 198986 560218 199222 560454
rect 198986 559898 199222 560134
rect 198986 524218 199222 524454
rect 198986 523898 199222 524134
rect 191786 517018 192022 517254
rect 191786 516698 192022 516934
rect 191786 481018 192022 481254
rect 191786 480698 192022 480934
rect 191786 445018 192022 445254
rect 191786 444698 192022 444934
rect 191786 409018 192022 409254
rect 191786 408698 192022 408934
rect 191786 373018 192022 373254
rect 191786 372698 192022 372934
rect 191786 337018 192022 337254
rect 191786 336698 192022 336934
rect 191786 301018 192022 301254
rect 191786 300698 192022 300934
rect 191786 265018 192022 265254
rect 191786 264698 192022 264934
rect 191786 229018 192022 229254
rect 191786 228698 192022 228934
rect 191786 193018 192022 193254
rect 191786 192698 192022 192934
rect 191786 157018 192022 157254
rect 191786 156698 192022 156934
rect 202586 671818 202822 672054
rect 202586 671498 202822 671734
rect 202586 635818 202822 636054
rect 202586 635498 202822 635734
rect 202586 599818 202822 600054
rect 202586 599498 202822 599734
rect 202586 563818 202822 564054
rect 202586 563498 202822 563734
rect 202586 527818 202822 528054
rect 202586 527498 202822 527734
rect 198986 488218 199222 488454
rect 198986 487898 199222 488134
rect 198986 452218 199222 452454
rect 198986 451898 199222 452134
rect 198986 416218 199222 416454
rect 198986 415898 199222 416134
rect 198986 380218 199222 380454
rect 198986 379898 199222 380134
rect 198986 344218 199222 344454
rect 198986 343898 199222 344134
rect 198986 308218 199222 308454
rect 198986 307898 199222 308134
rect 198986 272218 199222 272454
rect 198986 271898 199222 272134
rect 198986 236218 199222 236454
rect 198986 235898 199222 236134
rect 198986 200218 199222 200454
rect 198986 199898 199222 200134
rect 198986 164218 199222 164454
rect 198986 163898 199222 164134
rect 191786 121018 192022 121254
rect 191786 120698 192022 120934
rect 191786 85018 192022 85254
rect 191786 84698 192022 84934
rect 198986 128218 199222 128454
rect 198986 127898 199222 128134
rect 198986 92218 199222 92454
rect 198986 91898 199222 92134
rect 191786 49018 192022 49254
rect 191786 48698 192022 48934
rect 191786 13018 192022 13254
rect 191786 12698 192022 12934
rect 173786 -7022 174022 -6786
rect 173786 -7342 174022 -7106
rect 198986 56218 199222 56454
rect 198986 55898 199222 56134
rect 198986 20218 199222 20454
rect 198986 19898 199222 20134
rect 198986 -1502 199222 -1266
rect 198986 -1822 199222 -1586
rect 206186 675418 206422 675654
rect 206186 675098 206422 675334
rect 206186 639418 206422 639654
rect 206186 639098 206422 639334
rect 206186 603418 206422 603654
rect 206186 603098 206422 603334
rect 206186 567418 206422 567654
rect 206186 567098 206422 567334
rect 206186 531418 206422 531654
rect 206186 531098 206422 531334
rect 202586 491818 202822 492054
rect 202586 491498 202822 491734
rect 202586 455818 202822 456054
rect 202586 455498 202822 455734
rect 202586 419818 202822 420054
rect 202586 419498 202822 419734
rect 202586 383818 202822 384054
rect 202586 383498 202822 383734
rect 202586 347818 202822 348054
rect 202586 347498 202822 347734
rect 202586 311818 202822 312054
rect 202586 311498 202822 311734
rect 202586 275818 202822 276054
rect 202586 275498 202822 275734
rect 202586 239818 202822 240054
rect 202586 239498 202822 239734
rect 202586 203818 202822 204054
rect 202586 203498 202822 203734
rect 202586 167818 202822 168054
rect 202586 167498 202822 167734
rect 202586 131818 202822 132054
rect 202586 131498 202822 131734
rect 202586 95818 202822 96054
rect 202586 95498 202822 95734
rect 202586 59818 202822 60054
rect 202586 59498 202822 59734
rect 202586 23818 202822 24054
rect 202586 23498 202822 23734
rect 202586 -3342 202822 -3106
rect 202586 -3662 202822 -3426
rect 206186 495418 206422 495654
rect 206186 495098 206422 495334
rect 206186 459418 206422 459654
rect 206186 459098 206422 459334
rect 206186 423418 206422 423654
rect 206186 423098 206422 423334
rect 206186 387418 206422 387654
rect 206186 387098 206422 387334
rect 206186 351418 206422 351654
rect 206186 351098 206422 351334
rect 206186 315418 206422 315654
rect 206186 315098 206422 315334
rect 206186 279418 206422 279654
rect 206186 279098 206422 279334
rect 206186 243418 206422 243654
rect 206186 243098 206422 243334
rect 206186 207418 206422 207654
rect 206186 207098 206422 207334
rect 206186 171418 206422 171654
rect 206186 171098 206422 171334
rect 206186 135418 206422 135654
rect 206186 135098 206422 135334
rect 206186 99418 206422 99654
rect 206186 99098 206422 99334
rect 206186 63418 206422 63654
rect 206186 63098 206422 63334
rect 206186 27418 206422 27654
rect 206186 27098 206422 27334
rect 206186 -5182 206422 -4946
rect 206186 -5502 206422 -5266
rect 227786 710122 228022 710358
rect 227786 709802 228022 710038
rect 224186 708282 224422 708518
rect 224186 707962 224422 708198
rect 220586 706442 220822 706678
rect 220586 706122 220822 706358
rect 209786 679018 210022 679254
rect 209786 678698 210022 678934
rect 209786 643018 210022 643254
rect 209786 642698 210022 642934
rect 209786 607018 210022 607254
rect 209786 606698 210022 606934
rect 209786 571018 210022 571254
rect 209786 570698 210022 570934
rect 209786 535018 210022 535254
rect 209786 534698 210022 534934
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 216986 686218 217222 686454
rect 216986 685898 217222 686134
rect 216986 650218 217222 650454
rect 216986 649898 217222 650134
rect 216986 614218 217222 614454
rect 216986 613898 217222 614134
rect 216986 578218 217222 578454
rect 216986 577898 217222 578134
rect 216986 542218 217222 542454
rect 216986 541898 217222 542134
rect 210286 517924 210372 517938
rect 210372 517924 210436 517938
rect 210436 517924 210522 517938
rect 210286 517702 210522 517924
rect 209786 499018 210022 499254
rect 209786 498698 210022 498934
rect 209786 463018 210022 463254
rect 209786 462698 210022 462934
rect 209786 427018 210022 427254
rect 209786 426698 210022 426934
rect 209786 391018 210022 391254
rect 209786 390698 210022 390934
rect 209786 355018 210022 355254
rect 209786 354698 210022 354934
rect 209786 319018 210022 319254
rect 209786 318698 210022 318934
rect 209786 283018 210022 283254
rect 209786 282698 210022 282934
rect 209786 247018 210022 247254
rect 209786 246698 210022 246934
rect 209786 211018 210022 211254
rect 209786 210698 210022 210934
rect 209786 175018 210022 175254
rect 209786 174698 210022 174934
rect 209786 139018 210022 139254
rect 209786 138698 210022 138934
rect 209786 103018 210022 103254
rect 209786 102698 210022 102934
rect 209786 67018 210022 67254
rect 209786 66698 210022 66934
rect 209786 31018 210022 31254
rect 209786 30698 210022 30934
rect 191786 -6102 192022 -5866
rect 191786 -6422 192022 -6186
rect 220586 689818 220822 690054
rect 220586 689498 220822 689734
rect 220586 653818 220822 654054
rect 220586 653498 220822 653734
rect 220586 617818 220822 618054
rect 220586 617498 220822 617734
rect 220586 581818 220822 582054
rect 220586 581498 220822 581734
rect 220586 545818 220822 546054
rect 220586 545498 220822 545734
rect 219118 517924 219204 517938
rect 219204 517924 219268 517938
rect 219268 517924 219354 517938
rect 219118 517702 219354 517924
rect 216986 506218 217222 506454
rect 216986 505898 217222 506134
rect 216986 470218 217222 470454
rect 216986 469898 217222 470134
rect 216986 434218 217222 434454
rect 216986 433898 217222 434134
rect 216986 398218 217222 398454
rect 216986 397898 217222 398134
rect 216986 362218 217222 362454
rect 216986 361898 217222 362134
rect 216986 326218 217222 326454
rect 216986 325898 217222 326134
rect 216986 290218 217222 290454
rect 216986 289898 217222 290134
rect 216986 254218 217222 254454
rect 216986 253898 217222 254134
rect 216986 218218 217222 218454
rect 216986 217898 217222 218134
rect 216986 182218 217222 182454
rect 216986 181898 217222 182134
rect 216986 146218 217222 146454
rect 216986 145898 217222 146134
rect 216986 110218 217222 110454
rect 216986 109898 217222 110134
rect 216986 74218 217222 74454
rect 216986 73898 217222 74134
rect 216986 38218 217222 38454
rect 216986 37898 217222 38134
rect 216986 2218 217222 2454
rect 216986 1898 217222 2134
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 220586 509818 220822 510054
rect 220586 509498 220822 509734
rect 220586 473818 220822 474054
rect 220586 473498 220822 473734
rect 220586 437818 220822 438054
rect 220586 437498 220822 437734
rect 220586 401818 220822 402054
rect 220586 401498 220822 401734
rect 220586 365818 220822 366054
rect 220586 365498 220822 365734
rect 220586 329818 220822 330054
rect 220586 329498 220822 329734
rect 220586 293818 220822 294054
rect 220586 293498 220822 293734
rect 220586 257818 220822 258054
rect 220586 257498 220822 257734
rect 220586 221818 220822 222054
rect 220586 221498 220822 221734
rect 220586 185818 220822 186054
rect 220586 185498 220822 185734
rect 220586 149818 220822 150054
rect 220586 149498 220822 149734
rect 220586 113818 220822 114054
rect 220586 113498 220822 113734
rect 220586 77818 220822 78054
rect 220586 77498 220822 77734
rect 220586 41818 220822 42054
rect 220586 41498 220822 41734
rect 220586 5818 220822 6054
rect 220586 5498 220822 5734
rect 220586 -2422 220822 -2186
rect 220586 -2742 220822 -2506
rect 224186 693418 224422 693654
rect 224186 693098 224422 693334
rect 224186 657418 224422 657654
rect 224186 657098 224422 657334
rect 224186 621418 224422 621654
rect 224186 621098 224422 621334
rect 224186 585418 224422 585654
rect 224186 585098 224422 585334
rect 224186 549418 224422 549654
rect 224186 549098 224422 549334
rect 224186 513418 224422 513654
rect 224186 513098 224422 513334
rect 224186 477418 224422 477654
rect 224186 477098 224422 477334
rect 224186 441418 224422 441654
rect 224186 441098 224422 441334
rect 224186 405418 224422 405654
rect 224186 405098 224422 405334
rect 224186 369418 224422 369654
rect 224186 369098 224422 369334
rect 224186 333418 224422 333654
rect 224186 333098 224422 333334
rect 224186 297418 224422 297654
rect 224186 297098 224422 297334
rect 224186 261418 224422 261654
rect 224186 261098 224422 261334
rect 224186 225418 224422 225654
rect 224186 225098 224422 225334
rect 224186 189418 224422 189654
rect 224186 189098 224422 189334
rect 224186 153418 224422 153654
rect 224186 153098 224422 153334
rect 224186 117418 224422 117654
rect 224186 117098 224422 117334
rect 224186 81418 224422 81654
rect 224186 81098 224422 81334
rect 224186 45418 224422 45654
rect 224186 45098 224422 45334
rect 224186 9418 224422 9654
rect 224186 9098 224422 9334
rect 224186 -4262 224422 -4026
rect 224186 -4582 224422 -4346
rect 245786 711042 246022 711278
rect 245786 710722 246022 710958
rect 242186 709202 242422 709438
rect 242186 708882 242422 709118
rect 238586 707362 238822 707598
rect 238586 707042 238822 707278
rect 227786 697018 228022 697254
rect 227786 696698 228022 696934
rect 227786 661018 228022 661254
rect 227786 660698 228022 660934
rect 227786 625018 228022 625254
rect 227786 624698 228022 624934
rect 227786 589018 228022 589254
rect 227786 588698 228022 588934
rect 227786 553018 228022 553254
rect 227786 552698 228022 552934
rect 234986 705522 235222 705758
rect 234986 705202 235222 705438
rect 234986 668218 235222 668454
rect 234986 667898 235222 668134
rect 234986 632218 235222 632454
rect 234986 631898 235222 632134
rect 234986 596218 235222 596454
rect 234986 595898 235222 596134
rect 234986 560218 235222 560454
rect 234986 559898 235222 560134
rect 234986 524218 235222 524454
rect 234986 523898 235222 524134
rect 234390 517924 234476 517938
rect 234476 517924 234540 517938
rect 234540 517924 234626 517938
rect 234390 517702 234626 517924
rect 227786 517018 228022 517254
rect 227786 516698 228022 516934
rect 227786 481018 228022 481254
rect 227786 480698 228022 480934
rect 227786 445018 228022 445254
rect 227786 444698 228022 444934
rect 227786 409018 228022 409254
rect 227786 408698 228022 408934
rect 227786 373018 228022 373254
rect 227786 372698 228022 372934
rect 227786 337018 228022 337254
rect 227786 336698 228022 336934
rect 227786 301018 228022 301254
rect 227786 300698 228022 300934
rect 227786 265018 228022 265254
rect 227786 264698 228022 264934
rect 227786 229018 228022 229254
rect 227786 228698 228022 228934
rect 227786 193018 228022 193254
rect 227786 192698 228022 192934
rect 227786 157018 228022 157254
rect 227786 156698 228022 156934
rect 227786 121018 228022 121254
rect 227786 120698 228022 120934
rect 227786 85018 228022 85254
rect 227786 84698 228022 84934
rect 227786 49018 228022 49254
rect 227786 48698 228022 48934
rect 227786 13018 228022 13254
rect 227786 12698 228022 12934
rect 209786 -7022 210022 -6786
rect 209786 -7342 210022 -7106
rect 238586 671818 238822 672054
rect 238586 671498 238822 671734
rect 238586 635818 238822 636054
rect 238586 635498 238822 635734
rect 238586 599818 238822 600054
rect 238586 599498 238822 599734
rect 238586 563818 238822 564054
rect 238586 563498 238822 563734
rect 238586 527818 238822 528054
rect 238586 527498 238822 527734
rect 234986 488218 235222 488454
rect 234986 487898 235222 488134
rect 234986 452218 235222 452454
rect 234986 451898 235222 452134
rect 234986 416218 235222 416454
rect 234986 415898 235222 416134
rect 234986 380218 235222 380454
rect 234986 379898 235222 380134
rect 234986 344218 235222 344454
rect 234986 343898 235222 344134
rect 234986 308218 235222 308454
rect 234986 307898 235222 308134
rect 234986 272218 235222 272454
rect 234986 271898 235222 272134
rect 234986 236218 235222 236454
rect 234986 235898 235222 236134
rect 234986 200218 235222 200454
rect 234986 199898 235222 200134
rect 234986 164218 235222 164454
rect 234986 163898 235222 164134
rect 234986 128218 235222 128454
rect 234986 127898 235222 128134
rect 234986 92218 235222 92454
rect 234986 91898 235222 92134
rect 234986 56218 235222 56454
rect 234986 55898 235222 56134
rect 234986 20218 235222 20454
rect 234986 19898 235222 20134
rect 234986 -1502 235222 -1266
rect 234986 -1822 235222 -1586
rect 242186 675418 242422 675654
rect 242186 675098 242422 675334
rect 242186 639418 242422 639654
rect 242186 639098 242422 639334
rect 242186 603418 242422 603654
rect 242186 603098 242422 603334
rect 242186 567418 242422 567654
rect 242186 567098 242422 567334
rect 242186 531418 242422 531654
rect 242186 531098 242422 531334
rect 238586 491818 238822 492054
rect 238586 491498 238822 491734
rect 238586 455818 238822 456054
rect 238586 455498 238822 455734
rect 238586 419818 238822 420054
rect 238586 419498 238822 419734
rect 238586 383818 238822 384054
rect 238586 383498 238822 383734
rect 238586 347818 238822 348054
rect 238586 347498 238822 347734
rect 238586 311818 238822 312054
rect 238586 311498 238822 311734
rect 238586 275818 238822 276054
rect 238586 275498 238822 275734
rect 238586 239818 238822 240054
rect 238586 239498 238822 239734
rect 238586 203818 238822 204054
rect 238586 203498 238822 203734
rect 238586 167818 238822 168054
rect 238586 167498 238822 167734
rect 238586 131818 238822 132054
rect 238586 131498 238822 131734
rect 238586 95818 238822 96054
rect 238586 95498 238822 95734
rect 238586 59818 238822 60054
rect 238586 59498 238822 59734
rect 238586 23818 238822 24054
rect 238586 23498 238822 23734
rect 238586 -3342 238822 -3106
rect 238586 -3662 238822 -3426
rect 263786 710122 264022 710358
rect 263786 709802 264022 710038
rect 260186 708282 260422 708518
rect 260186 707962 260422 708198
rect 256586 706442 256822 706678
rect 256586 706122 256822 706358
rect 245786 679018 246022 679254
rect 245786 678698 246022 678934
rect 245786 643018 246022 643254
rect 245786 642698 246022 642934
rect 245786 607018 246022 607254
rect 245786 606698 246022 606934
rect 245786 571018 246022 571254
rect 245786 570698 246022 570934
rect 245786 535018 246022 535254
rect 245786 534698 246022 534934
rect 243590 517924 243676 517938
rect 243676 517924 243740 517938
rect 243740 517924 243826 517938
rect 243590 517702 243826 517924
rect 244694 517702 244930 517938
rect 242186 495418 242422 495654
rect 242186 495098 242422 495334
rect 242186 459418 242422 459654
rect 242186 459098 242422 459334
rect 242186 423418 242422 423654
rect 242186 423098 242422 423334
rect 242186 387418 242422 387654
rect 242186 387098 242422 387334
rect 242186 351418 242422 351654
rect 242186 351098 242422 351334
rect 242186 315418 242422 315654
rect 242186 315098 242422 315334
rect 242186 279418 242422 279654
rect 242186 279098 242422 279334
rect 242186 243418 242422 243654
rect 242186 243098 242422 243334
rect 242186 207418 242422 207654
rect 242186 207098 242422 207334
rect 242186 171418 242422 171654
rect 242186 171098 242422 171334
rect 242186 135418 242422 135654
rect 242186 135098 242422 135334
rect 242186 99418 242422 99654
rect 242186 99098 242422 99334
rect 242186 63418 242422 63654
rect 242186 63098 242422 63334
rect 242186 27418 242422 27654
rect 242186 27098 242422 27334
rect 242186 -5182 242422 -4946
rect 242186 -5502 242422 -5266
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 252986 686218 253222 686454
rect 252986 685898 253222 686134
rect 252986 650218 253222 650454
rect 252986 649898 253222 650134
rect 252986 614218 253222 614454
rect 252986 613898 253222 614134
rect 252986 578218 253222 578454
rect 252986 577898 253222 578134
rect 252986 542218 253222 542454
rect 252986 541898 253222 542134
rect 245786 499018 246022 499254
rect 245786 498698 246022 498934
rect 245786 463018 246022 463254
rect 245786 462698 246022 462934
rect 245786 427018 246022 427254
rect 245786 426698 246022 426934
rect 245786 391018 246022 391254
rect 245786 390698 246022 390934
rect 245786 355018 246022 355254
rect 245786 354698 246022 354934
rect 245786 319018 246022 319254
rect 245786 318698 246022 318934
rect 245786 283018 246022 283254
rect 245786 282698 246022 282934
rect 245786 247018 246022 247254
rect 245786 246698 246022 246934
rect 245786 211018 246022 211254
rect 245786 210698 246022 210934
rect 245786 175018 246022 175254
rect 245786 174698 246022 174934
rect 245786 139018 246022 139254
rect 245786 138698 246022 138934
rect 245786 103018 246022 103254
rect 245786 102698 246022 102934
rect 245786 67018 246022 67254
rect 245786 66698 246022 66934
rect 245786 31018 246022 31254
rect 245786 30698 246022 30934
rect 227786 -6102 228022 -5866
rect 227786 -6422 228022 -6186
rect 256586 689818 256822 690054
rect 256586 689498 256822 689734
rect 256586 653818 256822 654054
rect 256586 653498 256822 653734
rect 256586 617818 256822 618054
rect 256586 617498 256822 617734
rect 256586 581818 256822 582054
rect 256586 581498 256822 581734
rect 256586 545818 256822 546054
rect 256586 545498 256822 545734
rect 254078 517924 254164 517938
rect 254164 517924 254228 517938
rect 254228 517924 254314 517938
rect 254078 517702 254314 517924
rect 252986 506218 253222 506454
rect 252986 505898 253222 506134
rect 252986 470218 253222 470454
rect 252986 469898 253222 470134
rect 252986 434218 253222 434454
rect 252986 433898 253222 434134
rect 252986 398218 253222 398454
rect 252986 397898 253222 398134
rect 252986 362218 253222 362454
rect 252986 361898 253222 362134
rect 252986 326218 253222 326454
rect 252986 325898 253222 326134
rect 252986 290218 253222 290454
rect 252986 289898 253222 290134
rect 252986 254218 253222 254454
rect 252986 253898 253222 254134
rect 252986 218218 253222 218454
rect 252986 217898 253222 218134
rect 252986 182218 253222 182454
rect 252986 181898 253222 182134
rect 252986 146218 253222 146454
rect 252986 145898 253222 146134
rect 252986 110218 253222 110454
rect 252986 109898 253222 110134
rect 252986 74218 253222 74454
rect 252986 73898 253222 74134
rect 252986 38218 253222 38454
rect 252986 37898 253222 38134
rect 252986 2218 253222 2454
rect 252986 1898 253222 2134
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 256586 509818 256822 510054
rect 256586 509498 256822 509734
rect 256586 473818 256822 474054
rect 256586 473498 256822 473734
rect 256586 437818 256822 438054
rect 256586 437498 256822 437734
rect 256586 401818 256822 402054
rect 256586 401498 256822 401734
rect 256586 365818 256822 366054
rect 256586 365498 256822 365734
rect 256586 329818 256822 330054
rect 256586 329498 256822 329734
rect 256586 293818 256822 294054
rect 256586 293498 256822 293734
rect 256586 257818 256822 258054
rect 256586 257498 256822 257734
rect 256586 221818 256822 222054
rect 256586 221498 256822 221734
rect 256586 185818 256822 186054
rect 256586 185498 256822 185734
rect 256586 149818 256822 150054
rect 256586 149498 256822 149734
rect 256586 113818 256822 114054
rect 256586 113498 256822 113734
rect 256586 77818 256822 78054
rect 256586 77498 256822 77734
rect 256586 41818 256822 42054
rect 256586 41498 256822 41734
rect 256586 5818 256822 6054
rect 256586 5498 256822 5734
rect 256586 -2422 256822 -2186
rect 256586 -2742 256822 -2506
rect 260186 693418 260422 693654
rect 260186 693098 260422 693334
rect 260186 657418 260422 657654
rect 260186 657098 260422 657334
rect 260186 621418 260422 621654
rect 260186 621098 260422 621334
rect 260186 585418 260422 585654
rect 260186 585098 260422 585334
rect 260186 549418 260422 549654
rect 260186 549098 260422 549334
rect 281786 711042 282022 711278
rect 281786 710722 282022 710958
rect 278186 709202 278422 709438
rect 278186 708882 278422 709118
rect 274586 707362 274822 707598
rect 274586 707042 274822 707278
rect 263786 697018 264022 697254
rect 263786 696698 264022 696934
rect 263786 661018 264022 661254
rect 263786 660698 264022 660934
rect 270986 705522 271222 705758
rect 270986 705202 271222 705438
rect 270986 668218 271222 668454
rect 270986 667898 271222 668134
rect 263786 625018 264022 625254
rect 263786 624698 264022 624934
rect 263786 589018 264022 589254
rect 263786 588698 264022 588934
rect 263786 553018 264022 553254
rect 263786 552698 264022 552934
rect 260186 513418 260422 513654
rect 260186 513098 260422 513334
rect 260186 477418 260422 477654
rect 260186 477098 260422 477334
rect 260186 441418 260422 441654
rect 260186 441098 260422 441334
rect 260186 405418 260422 405654
rect 260186 405098 260422 405334
rect 260186 369418 260422 369654
rect 260186 369098 260422 369334
rect 260186 333418 260422 333654
rect 260186 333098 260422 333334
rect 260186 297418 260422 297654
rect 260186 297098 260422 297334
rect 260186 261418 260422 261654
rect 260186 261098 260422 261334
rect 260186 225418 260422 225654
rect 260186 225098 260422 225334
rect 260186 189418 260422 189654
rect 260186 189098 260422 189334
rect 260186 153418 260422 153654
rect 260186 153098 260422 153334
rect 260186 117418 260422 117654
rect 260186 117098 260422 117334
rect 260186 81418 260422 81654
rect 260186 81098 260422 81334
rect 260186 45418 260422 45654
rect 260186 45098 260422 45334
rect 260186 9418 260422 9654
rect 260186 9098 260422 9334
rect 260186 -4262 260422 -4026
rect 260186 -4582 260422 -4346
rect 270986 632218 271222 632454
rect 270986 631898 271222 632134
rect 270986 596218 271222 596454
rect 270986 595898 271222 596134
rect 270986 560218 271222 560454
rect 270986 559898 271222 560134
rect 270986 524218 271222 524454
rect 270986 523898 271222 524134
rect 264382 517924 264468 517938
rect 264468 517924 264532 517938
rect 264532 517924 264618 517938
rect 264382 517702 264618 517924
rect 263786 517018 264022 517254
rect 263786 516698 264022 516934
rect 263786 481018 264022 481254
rect 263786 480698 264022 480934
rect 263786 445018 264022 445254
rect 263786 444698 264022 444934
rect 263786 409018 264022 409254
rect 263786 408698 264022 408934
rect 263786 373018 264022 373254
rect 263786 372698 264022 372934
rect 263786 337018 264022 337254
rect 263786 336698 264022 336934
rect 263786 301018 264022 301254
rect 263786 300698 264022 300934
rect 263786 265018 264022 265254
rect 263786 264698 264022 264934
rect 263786 229018 264022 229254
rect 263786 228698 264022 228934
rect 263786 193018 264022 193254
rect 263786 192698 264022 192934
rect 263786 157018 264022 157254
rect 263786 156698 264022 156934
rect 263786 121018 264022 121254
rect 263786 120698 264022 120934
rect 263786 85018 264022 85254
rect 263786 84698 264022 84934
rect 263786 49018 264022 49254
rect 263786 48698 264022 48934
rect 263786 13018 264022 13254
rect 263786 12698 264022 12934
rect 245786 -7022 246022 -6786
rect 245786 -7342 246022 -7106
rect 274586 671818 274822 672054
rect 274586 671498 274822 671734
rect 274586 635818 274822 636054
rect 274586 635498 274822 635734
rect 274586 599818 274822 600054
rect 274586 599498 274822 599734
rect 274586 563818 274822 564054
rect 274586 563498 274822 563734
rect 274586 527818 274822 528054
rect 274586 527498 274822 527734
rect 273398 517924 273484 517938
rect 273484 517924 273548 517938
rect 273548 517924 273634 517938
rect 273398 517702 273634 517924
rect 270986 488218 271222 488454
rect 270986 487898 271222 488134
rect 270986 452218 271222 452454
rect 270986 451898 271222 452134
rect 270986 416218 271222 416454
rect 270986 415898 271222 416134
rect 270986 380218 271222 380454
rect 270986 379898 271222 380134
rect 270986 344218 271222 344454
rect 270986 343898 271222 344134
rect 270986 308218 271222 308454
rect 270986 307898 271222 308134
rect 270986 272218 271222 272454
rect 270986 271898 271222 272134
rect 270986 236218 271222 236454
rect 270986 235898 271222 236134
rect 270986 200218 271222 200454
rect 270986 199898 271222 200134
rect 270986 164218 271222 164454
rect 270986 163898 271222 164134
rect 270986 128218 271222 128454
rect 270986 127898 271222 128134
rect 270986 92218 271222 92454
rect 270986 91898 271222 92134
rect 270986 56218 271222 56454
rect 270986 55898 271222 56134
rect 270986 20218 271222 20454
rect 270986 19898 271222 20134
rect 270986 -1502 271222 -1266
rect 270986 -1822 271222 -1586
rect 274586 491818 274822 492054
rect 274586 491498 274822 491734
rect 274586 455818 274822 456054
rect 274586 455498 274822 455734
rect 274586 419818 274822 420054
rect 274586 419498 274822 419734
rect 274586 383818 274822 384054
rect 274586 383498 274822 383734
rect 274586 347818 274822 348054
rect 274586 347498 274822 347734
rect 274586 311818 274822 312054
rect 274586 311498 274822 311734
rect 274586 275818 274822 276054
rect 274586 275498 274822 275734
rect 274586 239818 274822 240054
rect 274586 239498 274822 239734
rect 278186 675418 278422 675654
rect 278186 675098 278422 675334
rect 278186 639418 278422 639654
rect 278186 639098 278422 639334
rect 278186 603418 278422 603654
rect 278186 603098 278422 603334
rect 278186 567418 278422 567654
rect 278186 567098 278422 567334
rect 278186 531418 278422 531654
rect 278186 531098 278422 531334
rect 299786 710122 300022 710358
rect 299786 709802 300022 710038
rect 296186 708282 296422 708518
rect 296186 707962 296422 708198
rect 292586 706442 292822 706678
rect 292586 706122 292822 706358
rect 281786 679018 282022 679254
rect 281786 678698 282022 678934
rect 281786 643018 282022 643254
rect 281786 642698 282022 642934
rect 281786 607018 282022 607254
rect 281786 606698 282022 606934
rect 281786 571018 282022 571254
rect 281786 570698 282022 570934
rect 281786 535018 282022 535254
rect 281786 534698 282022 534934
rect 278186 495418 278422 495654
rect 278186 495098 278422 495334
rect 278186 459418 278422 459654
rect 278186 459098 278422 459334
rect 278186 423418 278422 423654
rect 278186 423098 278422 423334
rect 278186 387418 278422 387654
rect 278186 387098 278422 387334
rect 278186 351418 278422 351654
rect 278186 351098 278422 351334
rect 278186 315418 278422 315654
rect 278186 315098 278422 315334
rect 278186 279418 278422 279654
rect 278186 279098 278422 279334
rect 278186 243418 278422 243654
rect 278186 243098 278422 243334
rect 274586 203818 274822 204054
rect 274586 203498 274822 203734
rect 274586 167818 274822 168054
rect 274586 167498 274822 167734
rect 278186 207418 278422 207654
rect 278186 207098 278422 207334
rect 278186 171418 278422 171654
rect 278186 171098 278422 171334
rect 274586 131818 274822 132054
rect 274586 131498 274822 131734
rect 274586 95818 274822 96054
rect 274586 95498 274822 95734
rect 274586 59818 274822 60054
rect 274586 59498 274822 59734
rect 274586 23818 274822 24054
rect 274586 23498 274822 23734
rect 274586 -3342 274822 -3106
rect 274586 -3662 274822 -3426
rect 278186 135418 278422 135654
rect 278186 135098 278422 135334
rect 278186 99418 278422 99654
rect 278186 99098 278422 99334
rect 278186 63418 278422 63654
rect 278186 63098 278422 63334
rect 278186 27418 278422 27654
rect 278186 27098 278422 27334
rect 278186 -5182 278422 -4946
rect 278186 -5502 278422 -5266
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 288986 686218 289222 686454
rect 288986 685898 289222 686134
rect 288986 650218 289222 650454
rect 288986 649898 289222 650134
rect 288986 614218 289222 614454
rect 288986 613898 289222 614134
rect 288986 578218 289222 578454
rect 288986 577898 289222 578134
rect 288986 542218 289222 542454
rect 288986 541898 289222 542134
rect 283334 517702 283570 517938
rect 281786 499018 282022 499254
rect 281786 498698 282022 498934
rect 281786 463018 282022 463254
rect 281786 462698 282022 462934
rect 281786 427018 282022 427254
rect 281786 426698 282022 426934
rect 281786 391018 282022 391254
rect 281786 390698 282022 390934
rect 281786 355018 282022 355254
rect 281786 354698 282022 354934
rect 281786 319018 282022 319254
rect 281786 318698 282022 318934
rect 281786 283018 282022 283254
rect 281786 282698 282022 282934
rect 281786 247018 282022 247254
rect 281786 246698 282022 246934
rect 281786 211018 282022 211254
rect 281786 210698 282022 210934
rect 281786 175018 282022 175254
rect 281786 174698 282022 174934
rect 281786 139018 282022 139254
rect 281786 138698 282022 138934
rect 288986 506218 289222 506454
rect 288986 505898 289222 506134
rect 288986 470218 289222 470454
rect 288986 469898 289222 470134
rect 288986 434218 289222 434454
rect 288986 433898 289222 434134
rect 288986 398218 289222 398454
rect 288986 397898 289222 398134
rect 288986 362218 289222 362454
rect 288986 361898 289222 362134
rect 288986 326218 289222 326454
rect 288986 325898 289222 326134
rect 288986 290218 289222 290454
rect 288986 289898 289222 290134
rect 288986 254218 289222 254454
rect 288986 253898 289222 254134
rect 288986 218218 289222 218454
rect 288986 217898 289222 218134
rect 288986 182218 289222 182454
rect 288986 181898 289222 182134
rect 288986 146218 289222 146454
rect 288986 145898 289222 146134
rect 288986 110218 289222 110454
rect 288986 109898 289222 110134
rect 281786 103018 282022 103254
rect 281786 102698 282022 102934
rect 281786 67018 282022 67254
rect 281786 66698 282022 66934
rect 281786 31018 282022 31254
rect 281786 30698 282022 30934
rect 263786 -6102 264022 -5866
rect 263786 -6422 264022 -6186
rect 288986 74218 289222 74454
rect 288986 73898 289222 74134
rect 288986 38218 289222 38454
rect 288986 37898 289222 38134
rect 288986 2218 289222 2454
rect 288986 1898 289222 2134
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 292586 689818 292822 690054
rect 292586 689498 292822 689734
rect 292586 653818 292822 654054
rect 292586 653498 292822 653734
rect 292586 617818 292822 618054
rect 292586 617498 292822 617734
rect 292586 581818 292822 582054
rect 292586 581498 292822 581734
rect 292586 545818 292822 546054
rect 292586 545498 292822 545734
rect 296186 693418 296422 693654
rect 296186 693098 296422 693334
rect 296186 657418 296422 657654
rect 296186 657098 296422 657334
rect 296186 621418 296422 621654
rect 296186 621098 296422 621334
rect 296186 585418 296422 585654
rect 296186 585098 296422 585334
rect 296186 549418 296422 549654
rect 296186 549098 296422 549334
rect 292586 509818 292822 510054
rect 292586 509498 292822 509734
rect 292586 473818 292822 474054
rect 292586 473498 292822 473734
rect 292586 437818 292822 438054
rect 292586 437498 292822 437734
rect 292586 401818 292822 402054
rect 292586 401498 292822 401734
rect 292586 365818 292822 366054
rect 292586 365498 292822 365734
rect 292586 329818 292822 330054
rect 292586 329498 292822 329734
rect 292586 293818 292822 294054
rect 292586 293498 292822 293734
rect 292586 257818 292822 258054
rect 292586 257498 292822 257734
rect 292586 221818 292822 222054
rect 292586 221498 292822 221734
rect 292586 185818 292822 186054
rect 292586 185498 292822 185734
rect 292586 149818 292822 150054
rect 292586 149498 292822 149734
rect 292586 113818 292822 114054
rect 292586 113498 292822 113734
rect 292586 77818 292822 78054
rect 292586 77498 292822 77734
rect 292586 41818 292822 42054
rect 292586 41498 292822 41734
rect 292586 5818 292822 6054
rect 292586 5498 292822 5734
rect 292586 -2422 292822 -2186
rect 292586 -2742 292822 -2506
rect 317786 711042 318022 711278
rect 317786 710722 318022 710958
rect 314186 709202 314422 709438
rect 314186 708882 314422 709118
rect 310586 707362 310822 707598
rect 310586 707042 310822 707278
rect 299786 697018 300022 697254
rect 299786 696698 300022 696934
rect 299786 661018 300022 661254
rect 299786 660698 300022 660934
rect 299786 625018 300022 625254
rect 299786 624698 300022 624934
rect 299786 589018 300022 589254
rect 299786 588698 300022 588934
rect 299786 553018 300022 553254
rect 299786 552698 300022 552934
rect 296186 513418 296422 513654
rect 296186 513098 296422 513334
rect 296186 477418 296422 477654
rect 296186 477098 296422 477334
rect 296186 441418 296422 441654
rect 296186 441098 296422 441334
rect 296186 405418 296422 405654
rect 296186 405098 296422 405334
rect 296186 369418 296422 369654
rect 296186 369098 296422 369334
rect 296186 333418 296422 333654
rect 296186 333098 296422 333334
rect 296186 297418 296422 297654
rect 296186 297098 296422 297334
rect 296186 261418 296422 261654
rect 296186 261098 296422 261334
rect 296186 225418 296422 225654
rect 296186 225098 296422 225334
rect 296186 189418 296422 189654
rect 296186 189098 296422 189334
rect 296186 153418 296422 153654
rect 296186 153098 296422 153334
rect 296186 117418 296422 117654
rect 296186 117098 296422 117334
rect 296186 81418 296422 81654
rect 296186 81098 296422 81334
rect 296186 45418 296422 45654
rect 296186 45098 296422 45334
rect 296186 9418 296422 9654
rect 296186 9098 296422 9334
rect 296186 -4262 296422 -4026
rect 296186 -4582 296422 -4346
rect 306986 705522 307222 705758
rect 306986 705202 307222 705438
rect 306986 668218 307222 668454
rect 306986 667898 307222 668134
rect 306986 632218 307222 632454
rect 306986 631898 307222 632134
rect 306986 596218 307222 596454
rect 306986 595898 307222 596134
rect 306986 560218 307222 560454
rect 306986 559898 307222 560134
rect 306986 524218 307222 524454
rect 306986 523898 307222 524134
rect 302654 517702 302890 517938
rect 299786 517018 300022 517254
rect 299786 516698 300022 516934
rect 299786 481018 300022 481254
rect 299786 480698 300022 480934
rect 299786 445018 300022 445254
rect 299786 444698 300022 444934
rect 299786 409018 300022 409254
rect 299786 408698 300022 408934
rect 299786 373018 300022 373254
rect 299786 372698 300022 372934
rect 299786 337018 300022 337254
rect 299786 336698 300022 336934
rect 299786 301018 300022 301254
rect 299786 300698 300022 300934
rect 299786 265018 300022 265254
rect 299786 264698 300022 264934
rect 299786 229018 300022 229254
rect 299786 228698 300022 228934
rect 299786 193018 300022 193254
rect 299786 192698 300022 192934
rect 299786 157018 300022 157254
rect 299786 156698 300022 156934
rect 299786 121018 300022 121254
rect 299786 120698 300022 120934
rect 299786 85018 300022 85254
rect 299786 84698 300022 84934
rect 299786 49018 300022 49254
rect 299786 48698 300022 48934
rect 299786 13018 300022 13254
rect 299786 12698 300022 12934
rect 281786 -7022 282022 -6786
rect 281786 -7342 282022 -7106
rect 310586 671818 310822 672054
rect 310586 671498 310822 671734
rect 310586 635818 310822 636054
rect 310586 635498 310822 635734
rect 310586 599818 310822 600054
rect 310586 599498 310822 599734
rect 310586 563818 310822 564054
rect 310586 563498 310822 563734
rect 310586 527818 310822 528054
rect 310586 527498 310822 527734
rect 306986 488218 307222 488454
rect 306986 487898 307222 488134
rect 306986 452218 307222 452454
rect 306986 451898 307222 452134
rect 306986 416218 307222 416454
rect 306986 415898 307222 416134
rect 306986 380218 307222 380454
rect 306986 379898 307222 380134
rect 306986 344218 307222 344454
rect 306986 343898 307222 344134
rect 306986 308218 307222 308454
rect 306986 307898 307222 308134
rect 306986 272218 307222 272454
rect 306986 271898 307222 272134
rect 306986 236218 307222 236454
rect 306986 235898 307222 236134
rect 306986 200218 307222 200454
rect 306986 199898 307222 200134
rect 306986 164218 307222 164454
rect 306986 163898 307222 164134
rect 306986 128218 307222 128454
rect 306986 127898 307222 128134
rect 306986 92218 307222 92454
rect 306986 91898 307222 92134
rect 306986 56218 307222 56454
rect 306986 55898 307222 56134
rect 314186 675418 314422 675654
rect 314186 675098 314422 675334
rect 314186 639418 314422 639654
rect 314186 639098 314422 639334
rect 314186 603418 314422 603654
rect 314186 603098 314422 603334
rect 314186 567418 314422 567654
rect 314186 567098 314422 567334
rect 314186 531418 314422 531654
rect 314186 531098 314422 531334
rect 310586 491818 310822 492054
rect 310586 491498 310822 491734
rect 310586 455818 310822 456054
rect 310586 455498 310822 455734
rect 310586 419818 310822 420054
rect 310586 419498 310822 419734
rect 310586 383818 310822 384054
rect 310586 383498 310822 383734
rect 310586 347818 310822 348054
rect 310586 347498 310822 347734
rect 310586 311818 310822 312054
rect 310586 311498 310822 311734
rect 310586 275818 310822 276054
rect 310586 275498 310822 275734
rect 310586 239818 310822 240054
rect 310586 239498 310822 239734
rect 310586 203818 310822 204054
rect 310586 203498 310822 203734
rect 310586 167818 310822 168054
rect 310586 167498 310822 167734
rect 310586 131818 310822 132054
rect 310586 131498 310822 131734
rect 310586 95818 310822 96054
rect 310586 95498 310822 95734
rect 310586 59818 310822 60054
rect 310586 59498 310822 59734
rect 306986 20218 307222 20454
rect 306986 19898 307222 20134
rect 306986 -1502 307222 -1266
rect 306986 -1822 307222 -1586
rect 310586 23818 310822 24054
rect 310586 23498 310822 23734
rect 310586 -3342 310822 -3106
rect 310586 -3662 310822 -3426
rect 314186 495418 314422 495654
rect 314186 495098 314422 495334
rect 314186 459418 314422 459654
rect 314186 459098 314422 459334
rect 314186 423418 314422 423654
rect 314186 423098 314422 423334
rect 314186 387418 314422 387654
rect 314186 387098 314422 387334
rect 314186 351418 314422 351654
rect 314186 351098 314422 351334
rect 314186 315418 314422 315654
rect 314186 315098 314422 315334
rect 314186 279418 314422 279654
rect 314186 279098 314422 279334
rect 314186 243418 314422 243654
rect 314186 243098 314422 243334
rect 314186 207418 314422 207654
rect 314186 207098 314422 207334
rect 314186 171418 314422 171654
rect 314186 171098 314422 171334
rect 314186 135418 314422 135654
rect 314186 135098 314422 135334
rect 314186 99418 314422 99654
rect 314186 99098 314422 99334
rect 314186 63418 314422 63654
rect 314186 63098 314422 63334
rect 314186 27418 314422 27654
rect 314186 27098 314422 27334
rect 314186 -5182 314422 -4946
rect 314186 -5502 314422 -5266
rect 335786 710122 336022 710358
rect 335786 709802 336022 710038
rect 332186 708282 332422 708518
rect 332186 707962 332422 708198
rect 328586 706442 328822 706678
rect 328586 706122 328822 706358
rect 317786 679018 318022 679254
rect 317786 678698 318022 678934
rect 317786 643018 318022 643254
rect 317786 642698 318022 642934
rect 317786 607018 318022 607254
rect 317786 606698 318022 606934
rect 317786 571018 318022 571254
rect 317786 570698 318022 570934
rect 317786 535018 318022 535254
rect 317786 534698 318022 534934
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 324986 686218 325222 686454
rect 324986 685898 325222 686134
rect 324986 650218 325222 650454
rect 324986 649898 325222 650134
rect 324986 614218 325222 614454
rect 324986 613898 325222 614134
rect 324986 578218 325222 578454
rect 324986 577898 325222 578134
rect 324986 542218 325222 542454
rect 324986 541898 325222 542134
rect 317786 499018 318022 499254
rect 317786 498698 318022 498934
rect 317786 463018 318022 463254
rect 317786 462698 318022 462934
rect 317786 427018 318022 427254
rect 317786 426698 318022 426934
rect 317786 391018 318022 391254
rect 317786 390698 318022 390934
rect 317786 355018 318022 355254
rect 317786 354698 318022 354934
rect 317786 319018 318022 319254
rect 317786 318698 318022 318934
rect 317786 283018 318022 283254
rect 317786 282698 318022 282934
rect 317786 247018 318022 247254
rect 317786 246698 318022 246934
rect 317786 211018 318022 211254
rect 317786 210698 318022 210934
rect 317786 175018 318022 175254
rect 317786 174698 318022 174934
rect 324986 506218 325222 506454
rect 324986 505898 325222 506134
rect 324986 470218 325222 470454
rect 324986 469898 325222 470134
rect 324986 434218 325222 434454
rect 324986 433898 325222 434134
rect 324986 398218 325222 398454
rect 324986 397898 325222 398134
rect 324986 362218 325222 362454
rect 324986 361898 325222 362134
rect 324986 326218 325222 326454
rect 324986 325898 325222 326134
rect 324986 290218 325222 290454
rect 324986 289898 325222 290134
rect 324986 254218 325222 254454
rect 324986 253898 325222 254134
rect 324986 218218 325222 218454
rect 324986 217898 325222 218134
rect 324986 182218 325222 182454
rect 324986 181898 325222 182134
rect 324986 146218 325222 146454
rect 324986 145898 325222 146134
rect 317786 139018 318022 139254
rect 317786 138698 318022 138934
rect 317786 103018 318022 103254
rect 317786 102698 318022 102934
rect 317786 67018 318022 67254
rect 317786 66698 318022 66934
rect 317786 31018 318022 31254
rect 317786 30698 318022 30934
rect 299786 -6102 300022 -5866
rect 299786 -6422 300022 -6186
rect 324986 110218 325222 110454
rect 324986 109898 325222 110134
rect 324986 74218 325222 74454
rect 324986 73898 325222 74134
rect 328586 689818 328822 690054
rect 328586 689498 328822 689734
rect 328586 653818 328822 654054
rect 328586 653498 328822 653734
rect 328586 617818 328822 618054
rect 328586 617498 328822 617734
rect 328586 581818 328822 582054
rect 328586 581498 328822 581734
rect 328586 545818 328822 546054
rect 328586 545498 328822 545734
rect 328586 509818 328822 510054
rect 328586 509498 328822 509734
rect 328586 473818 328822 474054
rect 328586 473498 328822 473734
rect 328586 437818 328822 438054
rect 328586 437498 328822 437734
rect 328586 401818 328822 402054
rect 328586 401498 328822 401734
rect 328586 365818 328822 366054
rect 328586 365498 328822 365734
rect 328586 329818 328822 330054
rect 328586 329498 328822 329734
rect 328586 293818 328822 294054
rect 328586 293498 328822 293734
rect 328586 257818 328822 258054
rect 328586 257498 328822 257734
rect 328586 221818 328822 222054
rect 328586 221498 328822 221734
rect 328586 185818 328822 186054
rect 328586 185498 328822 185734
rect 328586 149818 328822 150054
rect 328586 149498 328822 149734
rect 332186 693418 332422 693654
rect 332186 693098 332422 693334
rect 332186 657418 332422 657654
rect 332186 657098 332422 657334
rect 332186 621418 332422 621654
rect 332186 621098 332422 621334
rect 332186 585418 332422 585654
rect 332186 585098 332422 585334
rect 332186 549418 332422 549654
rect 332186 549098 332422 549334
rect 353786 711042 354022 711278
rect 353786 710722 354022 710958
rect 350186 709202 350422 709438
rect 350186 708882 350422 709118
rect 346586 707362 346822 707598
rect 346586 707042 346822 707278
rect 335786 697018 336022 697254
rect 335786 696698 336022 696934
rect 335786 661018 336022 661254
rect 335786 660698 336022 660934
rect 335786 625018 336022 625254
rect 335786 624698 336022 624934
rect 335786 589018 336022 589254
rect 335786 588698 336022 588934
rect 335786 553018 336022 553254
rect 335786 552698 336022 552934
rect 335222 517702 335458 517938
rect 332186 513418 332422 513654
rect 332186 513098 332422 513334
rect 332186 477418 332422 477654
rect 332186 477098 332422 477334
rect 332186 441418 332422 441654
rect 332186 441098 332422 441334
rect 332186 405418 332422 405654
rect 332186 405098 332422 405334
rect 332186 369418 332422 369654
rect 332186 369098 332422 369334
rect 332186 333418 332422 333654
rect 332186 333098 332422 333334
rect 332186 297418 332422 297654
rect 332186 297098 332422 297334
rect 332186 261418 332422 261654
rect 332186 261098 332422 261334
rect 332186 225418 332422 225654
rect 332186 225098 332422 225334
rect 332186 189418 332422 189654
rect 332186 189098 332422 189334
rect 332186 153418 332422 153654
rect 332186 153098 332422 153334
rect 328586 113818 328822 114054
rect 328586 113498 328822 113734
rect 332186 117418 332422 117654
rect 332186 117098 332422 117334
rect 328586 77818 328822 78054
rect 328586 77498 328822 77734
rect 332186 81418 332422 81654
rect 332186 81098 332422 81334
rect 328586 41818 328822 42054
rect 328586 41498 328822 41734
rect 324986 38218 325222 38454
rect 324986 37898 325222 38134
rect 324986 2218 325222 2454
rect 324986 1898 325222 2134
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 328586 5818 328822 6054
rect 328586 5498 328822 5734
rect 328586 -2422 328822 -2186
rect 328586 -2742 328822 -2506
rect 332186 45418 332422 45654
rect 332186 45098 332422 45334
rect 332186 9418 332422 9654
rect 332186 9098 332422 9334
rect 332186 -4262 332422 -4026
rect 332186 -4582 332422 -4346
rect 342986 705522 343222 705758
rect 342986 705202 343222 705438
rect 342986 668218 343222 668454
rect 342986 667898 343222 668134
rect 342986 632218 343222 632454
rect 342986 631898 343222 632134
rect 342986 596218 343222 596454
rect 342986 595898 343222 596134
rect 342986 560218 343222 560454
rect 342986 559898 343222 560134
rect 342986 524218 343222 524454
rect 342986 523898 343222 524134
rect 336326 517702 336562 517938
rect 335786 517018 336022 517254
rect 335786 516698 336022 516934
rect 335786 481018 336022 481254
rect 335786 480698 336022 480934
rect 335786 445018 336022 445254
rect 335786 444698 336022 444934
rect 335786 409018 336022 409254
rect 335786 408698 336022 408934
rect 335786 373018 336022 373254
rect 335786 372698 336022 372934
rect 335786 337018 336022 337254
rect 335786 336698 336022 336934
rect 335786 301018 336022 301254
rect 335786 300698 336022 300934
rect 335786 265018 336022 265254
rect 335786 264698 336022 264934
rect 335786 229018 336022 229254
rect 335786 228698 336022 228934
rect 335786 193018 336022 193254
rect 335786 192698 336022 192934
rect 335786 157018 336022 157254
rect 335786 156698 336022 156934
rect 335786 121018 336022 121254
rect 335786 120698 336022 120934
rect 335786 85018 336022 85254
rect 335786 84698 336022 84934
rect 335786 49018 336022 49254
rect 335786 48698 336022 48934
rect 342986 488218 343222 488454
rect 342986 487898 343222 488134
rect 342986 452218 343222 452454
rect 342986 451898 343222 452134
rect 342986 416218 343222 416454
rect 342986 415898 343222 416134
rect 342986 380218 343222 380454
rect 342986 379898 343222 380134
rect 342986 344218 343222 344454
rect 342986 343898 343222 344134
rect 342986 308218 343222 308454
rect 342986 307898 343222 308134
rect 342986 272218 343222 272454
rect 342986 271898 343222 272134
rect 342986 236218 343222 236454
rect 342986 235898 343222 236134
rect 342986 200218 343222 200454
rect 342986 199898 343222 200134
rect 342986 164218 343222 164454
rect 342986 163898 343222 164134
rect 342986 128218 343222 128454
rect 342986 127898 343222 128134
rect 342986 92218 343222 92454
rect 342986 91898 343222 92134
rect 342986 56218 343222 56454
rect 342986 55898 343222 56134
rect 335786 13018 336022 13254
rect 335786 12698 336022 12934
rect 317786 -7022 318022 -6786
rect 317786 -7342 318022 -7106
rect 342986 20218 343222 20454
rect 342986 19898 343222 20134
rect 342986 -1502 343222 -1266
rect 342986 -1822 343222 -1586
rect 346586 671818 346822 672054
rect 346586 671498 346822 671734
rect 346586 635818 346822 636054
rect 346586 635498 346822 635734
rect 346586 599818 346822 600054
rect 346586 599498 346822 599734
rect 346586 563818 346822 564054
rect 346586 563498 346822 563734
rect 346586 527818 346822 528054
rect 346586 527498 346822 527734
rect 346586 491818 346822 492054
rect 346586 491498 346822 491734
rect 346586 455818 346822 456054
rect 346586 455498 346822 455734
rect 346586 419818 346822 420054
rect 346586 419498 346822 419734
rect 346586 383818 346822 384054
rect 346586 383498 346822 383734
rect 346586 347818 346822 348054
rect 346586 347498 346822 347734
rect 346586 311818 346822 312054
rect 346586 311498 346822 311734
rect 346586 275818 346822 276054
rect 346586 275498 346822 275734
rect 346586 239818 346822 240054
rect 346586 239498 346822 239734
rect 346586 203818 346822 204054
rect 346586 203498 346822 203734
rect 346586 167818 346822 168054
rect 346586 167498 346822 167734
rect 346586 131818 346822 132054
rect 346586 131498 346822 131734
rect 346586 95818 346822 96054
rect 346586 95498 346822 95734
rect 346586 59818 346822 60054
rect 346586 59498 346822 59734
rect 346586 23818 346822 24054
rect 346586 23498 346822 23734
rect 346586 -3342 346822 -3106
rect 346586 -3662 346822 -3426
rect 350186 675418 350422 675654
rect 350186 675098 350422 675334
rect 350186 639418 350422 639654
rect 350186 639098 350422 639334
rect 350186 603418 350422 603654
rect 350186 603098 350422 603334
rect 350186 567418 350422 567654
rect 350186 567098 350422 567334
rect 350186 531418 350422 531654
rect 350186 531098 350422 531334
rect 350186 495418 350422 495654
rect 350186 495098 350422 495334
rect 350186 459418 350422 459654
rect 350186 459098 350422 459334
rect 350186 423418 350422 423654
rect 350186 423098 350422 423334
rect 350186 387418 350422 387654
rect 350186 387098 350422 387334
rect 350186 351418 350422 351654
rect 350186 351098 350422 351334
rect 350186 315418 350422 315654
rect 350186 315098 350422 315334
rect 350186 279418 350422 279654
rect 350186 279098 350422 279334
rect 350186 243418 350422 243654
rect 350186 243098 350422 243334
rect 350186 207418 350422 207654
rect 350186 207098 350422 207334
rect 350186 171418 350422 171654
rect 350186 171098 350422 171334
rect 350186 135418 350422 135654
rect 350186 135098 350422 135334
rect 350186 99418 350422 99654
rect 350186 99098 350422 99334
rect 350186 63418 350422 63654
rect 350186 63098 350422 63334
rect 350186 27418 350422 27654
rect 350186 27098 350422 27334
rect 350186 -5182 350422 -4946
rect 350186 -5502 350422 -5266
rect 371786 710122 372022 710358
rect 371786 709802 372022 710038
rect 368186 708282 368422 708518
rect 368186 707962 368422 708198
rect 364586 706442 364822 706678
rect 364586 706122 364822 706358
rect 353786 679018 354022 679254
rect 353786 678698 354022 678934
rect 353786 643018 354022 643254
rect 353786 642698 354022 642934
rect 353786 607018 354022 607254
rect 353786 606698 354022 606934
rect 353786 571018 354022 571254
rect 353786 570698 354022 570934
rect 353786 535018 354022 535254
rect 353786 534698 354022 534934
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 360986 686218 361222 686454
rect 360986 685898 361222 686134
rect 360986 650218 361222 650454
rect 360986 649898 361222 650134
rect 360986 614218 361222 614454
rect 360986 613898 361222 614134
rect 360986 578218 361222 578454
rect 360986 577898 361222 578134
rect 360986 542218 361222 542454
rect 360986 541898 361222 542134
rect 353786 499018 354022 499254
rect 353786 498698 354022 498934
rect 353786 463018 354022 463254
rect 353786 462698 354022 462934
rect 353786 427018 354022 427254
rect 353786 426698 354022 426934
rect 353786 391018 354022 391254
rect 353786 390698 354022 390934
rect 353786 355018 354022 355254
rect 353786 354698 354022 354934
rect 353786 319018 354022 319254
rect 353786 318698 354022 318934
rect 353786 283018 354022 283254
rect 353786 282698 354022 282934
rect 353786 247018 354022 247254
rect 353786 246698 354022 246934
rect 353786 211018 354022 211254
rect 353786 210698 354022 210934
rect 353786 175018 354022 175254
rect 353786 174698 354022 174934
rect 353786 139018 354022 139254
rect 353786 138698 354022 138934
rect 353786 103018 354022 103254
rect 353786 102698 354022 102934
rect 353786 67018 354022 67254
rect 353786 66698 354022 66934
rect 364586 689818 364822 690054
rect 364586 689498 364822 689734
rect 364586 653818 364822 654054
rect 364586 653498 364822 653734
rect 364586 617818 364822 618054
rect 364586 617498 364822 617734
rect 364586 581818 364822 582054
rect 364586 581498 364822 581734
rect 364586 545818 364822 546054
rect 364586 545498 364822 545734
rect 360986 506218 361222 506454
rect 360986 505898 361222 506134
rect 360986 470218 361222 470454
rect 360986 469898 361222 470134
rect 360986 434218 361222 434454
rect 360986 433898 361222 434134
rect 360986 398218 361222 398454
rect 360986 397898 361222 398134
rect 360986 362218 361222 362454
rect 360986 361898 361222 362134
rect 360986 326218 361222 326454
rect 360986 325898 361222 326134
rect 360986 290218 361222 290454
rect 360986 289898 361222 290134
rect 360986 254218 361222 254454
rect 360986 253898 361222 254134
rect 360986 218218 361222 218454
rect 360986 217898 361222 218134
rect 360986 182218 361222 182454
rect 360986 181898 361222 182134
rect 360986 146218 361222 146454
rect 360986 145898 361222 146134
rect 360986 110218 361222 110454
rect 360986 109898 361222 110134
rect 360986 74218 361222 74454
rect 360986 73898 361222 74134
rect 353786 31018 354022 31254
rect 353786 30698 354022 30934
rect 335786 -6102 336022 -5866
rect 335786 -6422 336022 -6186
rect 360986 38218 361222 38454
rect 360986 37898 361222 38134
rect 368186 693418 368422 693654
rect 368186 693098 368422 693334
rect 368186 657418 368422 657654
rect 368186 657098 368422 657334
rect 368186 621418 368422 621654
rect 368186 621098 368422 621334
rect 368186 585418 368422 585654
rect 368186 585098 368422 585334
rect 368186 549418 368422 549654
rect 368186 549098 368422 549334
rect 364586 509818 364822 510054
rect 364586 509498 364822 509734
rect 364586 473818 364822 474054
rect 364586 473498 364822 473734
rect 364586 437818 364822 438054
rect 364586 437498 364822 437734
rect 364586 401818 364822 402054
rect 364586 401498 364822 401734
rect 364586 365818 364822 366054
rect 364586 365498 364822 365734
rect 364586 329818 364822 330054
rect 364586 329498 364822 329734
rect 364586 293818 364822 294054
rect 364586 293498 364822 293734
rect 364586 257818 364822 258054
rect 364586 257498 364822 257734
rect 364586 221818 364822 222054
rect 364586 221498 364822 221734
rect 389786 711042 390022 711278
rect 389786 710722 390022 710958
rect 386186 709202 386422 709438
rect 386186 708882 386422 709118
rect 382586 707362 382822 707598
rect 382586 707042 382822 707278
rect 371786 697018 372022 697254
rect 371786 696698 372022 696934
rect 371786 661018 372022 661254
rect 371786 660698 372022 660934
rect 371786 625018 372022 625254
rect 371786 624698 372022 624934
rect 371786 589018 372022 589254
rect 371786 588698 372022 588934
rect 371786 553018 372022 553254
rect 371786 552698 372022 552934
rect 368186 513418 368422 513654
rect 368186 513098 368422 513334
rect 368186 477418 368422 477654
rect 368186 477098 368422 477334
rect 368186 441418 368422 441654
rect 368186 441098 368422 441334
rect 368186 405418 368422 405654
rect 368186 405098 368422 405334
rect 368186 369418 368422 369654
rect 368186 369098 368422 369334
rect 368186 333418 368422 333654
rect 368186 333098 368422 333334
rect 371786 517018 372022 517254
rect 371786 516698 372022 516934
rect 371786 481018 372022 481254
rect 371786 480698 372022 480934
rect 371786 445018 372022 445254
rect 371786 444698 372022 444934
rect 371786 409018 372022 409254
rect 371786 408698 372022 408934
rect 371786 373018 372022 373254
rect 371786 372698 372022 372934
rect 371786 337018 372022 337254
rect 371786 336698 372022 336934
rect 368186 297418 368422 297654
rect 368186 297098 368422 297334
rect 368186 261418 368422 261654
rect 368186 261098 368422 261334
rect 368186 225418 368422 225654
rect 368186 225098 368422 225334
rect 364586 185818 364822 186054
rect 364586 185498 364822 185734
rect 364586 149818 364822 150054
rect 364586 149498 364822 149734
rect 364586 113818 364822 114054
rect 364586 113498 364822 113734
rect 364586 77818 364822 78054
rect 364586 77498 364822 77734
rect 364586 41818 364822 42054
rect 364586 41498 364822 41734
rect 360986 2218 361222 2454
rect 360986 1898 361222 2134
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 364586 5818 364822 6054
rect 364586 5498 364822 5734
rect 364586 -2422 364822 -2186
rect 364586 -2742 364822 -2506
rect 368186 189418 368422 189654
rect 368186 189098 368422 189334
rect 368186 153418 368422 153654
rect 368186 153098 368422 153334
rect 368186 117418 368422 117654
rect 368186 117098 368422 117334
rect 368186 81418 368422 81654
rect 368186 81098 368422 81334
rect 368186 45418 368422 45654
rect 368186 45098 368422 45334
rect 368186 9418 368422 9654
rect 368186 9098 368422 9334
rect 368186 -4262 368422 -4026
rect 368186 -4582 368422 -4346
rect 371786 301018 372022 301254
rect 371786 300698 372022 300934
rect 371786 265018 372022 265254
rect 371786 264698 372022 264934
rect 371786 229018 372022 229254
rect 371786 228698 372022 228934
rect 371786 193018 372022 193254
rect 371786 192698 372022 192934
rect 371786 157018 372022 157254
rect 371786 156698 372022 156934
rect 371786 121018 372022 121254
rect 371786 120698 372022 120934
rect 371786 85018 372022 85254
rect 371786 84698 372022 84934
rect 371786 49018 372022 49254
rect 371786 48698 372022 48934
rect 371786 13018 372022 13254
rect 371786 12698 372022 12934
rect 353786 -7022 354022 -6786
rect 353786 -7342 354022 -7106
rect 378986 705522 379222 705758
rect 378986 705202 379222 705438
rect 378986 668218 379222 668454
rect 378986 667898 379222 668134
rect 378986 632218 379222 632454
rect 378986 631898 379222 632134
rect 378986 596218 379222 596454
rect 378986 595898 379222 596134
rect 378986 560218 379222 560454
rect 378986 559898 379222 560134
rect 378986 524218 379222 524454
rect 378986 523898 379222 524134
rect 378986 488218 379222 488454
rect 378986 487898 379222 488134
rect 378986 452218 379222 452454
rect 378986 451898 379222 452134
rect 378986 416218 379222 416454
rect 378986 415898 379222 416134
rect 378986 380218 379222 380454
rect 378986 379898 379222 380134
rect 378986 344218 379222 344454
rect 378986 343898 379222 344134
rect 378986 308218 379222 308454
rect 378986 307898 379222 308134
rect 378986 272218 379222 272454
rect 378986 271898 379222 272134
rect 378986 236218 379222 236454
rect 378986 235898 379222 236134
rect 378986 200218 379222 200454
rect 378986 199898 379222 200134
rect 378986 164218 379222 164454
rect 378986 163898 379222 164134
rect 378986 128218 379222 128454
rect 378986 127898 379222 128134
rect 378986 92218 379222 92454
rect 378986 91898 379222 92134
rect 378986 56218 379222 56454
rect 378986 55898 379222 56134
rect 378986 20218 379222 20454
rect 378986 19898 379222 20134
rect 378986 -1502 379222 -1266
rect 378986 -1822 379222 -1586
rect 382586 671818 382822 672054
rect 382586 671498 382822 671734
rect 382586 635818 382822 636054
rect 382586 635498 382822 635734
rect 382586 599818 382822 600054
rect 382586 599498 382822 599734
rect 382586 563818 382822 564054
rect 382586 563498 382822 563734
rect 382586 527818 382822 528054
rect 382586 527498 382822 527734
rect 382586 491818 382822 492054
rect 382586 491498 382822 491734
rect 386186 675418 386422 675654
rect 386186 675098 386422 675334
rect 386186 639418 386422 639654
rect 386186 639098 386422 639334
rect 386186 603418 386422 603654
rect 386186 603098 386422 603334
rect 386186 567418 386422 567654
rect 386186 567098 386422 567334
rect 386186 531418 386422 531654
rect 386186 531098 386422 531334
rect 386186 495418 386422 495654
rect 386186 495098 386422 495334
rect 382586 455818 382822 456054
rect 382586 455498 382822 455734
rect 382586 419818 382822 420054
rect 382586 419498 382822 419734
rect 382586 383818 382822 384054
rect 382586 383498 382822 383734
rect 382586 347818 382822 348054
rect 382586 347498 382822 347734
rect 382586 311818 382822 312054
rect 382586 311498 382822 311734
rect 382586 275818 382822 276054
rect 382586 275498 382822 275734
rect 382586 239818 382822 240054
rect 382586 239498 382822 239734
rect 382586 203818 382822 204054
rect 382586 203498 382822 203734
rect 382586 167818 382822 168054
rect 382586 167498 382822 167734
rect 382586 131818 382822 132054
rect 382586 131498 382822 131734
rect 382586 95818 382822 96054
rect 382586 95498 382822 95734
rect 382586 59818 382822 60054
rect 382586 59498 382822 59734
rect 386186 459418 386422 459654
rect 386186 459098 386422 459334
rect 386186 423418 386422 423654
rect 386186 423098 386422 423334
rect 386186 387418 386422 387654
rect 386186 387098 386422 387334
rect 386186 351418 386422 351654
rect 386186 351098 386422 351334
rect 386186 315418 386422 315654
rect 386186 315098 386422 315334
rect 386186 279418 386422 279654
rect 386186 279098 386422 279334
rect 386186 243418 386422 243654
rect 386186 243098 386422 243334
rect 386186 207418 386422 207654
rect 386186 207098 386422 207334
rect 386186 171418 386422 171654
rect 386186 171098 386422 171334
rect 386186 135418 386422 135654
rect 386186 135098 386422 135334
rect 386186 99418 386422 99654
rect 386186 99098 386422 99334
rect 386186 63418 386422 63654
rect 386186 63098 386422 63334
rect 382586 23818 382822 24054
rect 382586 23498 382822 23734
rect 382586 -3342 382822 -3106
rect 382586 -3662 382822 -3426
rect 386186 27418 386422 27654
rect 386186 27098 386422 27334
rect 386186 -5182 386422 -4946
rect 386186 -5502 386422 -5266
rect 407786 710122 408022 710358
rect 407786 709802 408022 710038
rect 404186 708282 404422 708518
rect 404186 707962 404422 708198
rect 400586 706442 400822 706678
rect 400586 706122 400822 706358
rect 389786 679018 390022 679254
rect 389786 678698 390022 678934
rect 389786 643018 390022 643254
rect 389786 642698 390022 642934
rect 389786 607018 390022 607254
rect 389786 606698 390022 606934
rect 389786 571018 390022 571254
rect 389786 570698 390022 570934
rect 389786 535018 390022 535254
rect 389786 534698 390022 534934
rect 389786 499018 390022 499254
rect 389786 498698 390022 498934
rect 389786 463018 390022 463254
rect 389786 462698 390022 462934
rect 389786 427018 390022 427254
rect 389786 426698 390022 426934
rect 389786 391018 390022 391254
rect 389786 390698 390022 390934
rect 389786 355018 390022 355254
rect 389786 354698 390022 354934
rect 389786 319018 390022 319254
rect 389786 318698 390022 318934
rect 389786 283018 390022 283254
rect 389786 282698 390022 282934
rect 389786 247018 390022 247254
rect 389786 246698 390022 246934
rect 389786 211018 390022 211254
rect 389786 210698 390022 210934
rect 389786 175018 390022 175254
rect 389786 174698 390022 174934
rect 389786 139018 390022 139254
rect 389786 138698 390022 138934
rect 389786 103018 390022 103254
rect 389786 102698 390022 102934
rect 389786 67018 390022 67254
rect 389786 66698 390022 66934
rect 389786 31018 390022 31254
rect 389786 30698 390022 30934
rect 371786 -6102 372022 -5866
rect 371786 -6422 372022 -6186
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 396986 686218 397222 686454
rect 396986 685898 397222 686134
rect 396986 650218 397222 650454
rect 396986 649898 397222 650134
rect 396986 614218 397222 614454
rect 396986 613898 397222 614134
rect 396986 578218 397222 578454
rect 396986 577898 397222 578134
rect 396986 542218 397222 542454
rect 396986 541898 397222 542134
rect 396986 506218 397222 506454
rect 396986 505898 397222 506134
rect 396986 470218 397222 470454
rect 396986 469898 397222 470134
rect 396986 434218 397222 434454
rect 396986 433898 397222 434134
rect 396986 398218 397222 398454
rect 396986 397898 397222 398134
rect 396986 362218 397222 362454
rect 396986 361898 397222 362134
rect 396986 326218 397222 326454
rect 396986 325898 397222 326134
rect 396986 290218 397222 290454
rect 396986 289898 397222 290134
rect 396986 254218 397222 254454
rect 396986 253898 397222 254134
rect 396986 218218 397222 218454
rect 396986 217898 397222 218134
rect 396986 182218 397222 182454
rect 396986 181898 397222 182134
rect 396986 146218 397222 146454
rect 396986 145898 397222 146134
rect 396986 110218 397222 110454
rect 396986 109898 397222 110134
rect 396986 74218 397222 74454
rect 396986 73898 397222 74134
rect 396986 38218 397222 38454
rect 396986 37898 397222 38134
rect 396986 2218 397222 2454
rect 396986 1898 397222 2134
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 400586 689818 400822 690054
rect 400586 689498 400822 689734
rect 400586 653818 400822 654054
rect 400586 653498 400822 653734
rect 400586 617818 400822 618054
rect 400586 617498 400822 617734
rect 400586 581818 400822 582054
rect 400586 581498 400822 581734
rect 400586 545818 400822 546054
rect 400586 545498 400822 545734
rect 400586 509818 400822 510054
rect 400586 509498 400822 509734
rect 400586 473818 400822 474054
rect 400586 473498 400822 473734
rect 400586 437818 400822 438054
rect 400586 437498 400822 437734
rect 400586 401818 400822 402054
rect 400586 401498 400822 401734
rect 400586 365818 400822 366054
rect 400586 365498 400822 365734
rect 400586 329818 400822 330054
rect 400586 329498 400822 329734
rect 400586 293818 400822 294054
rect 400586 293498 400822 293734
rect 400586 257818 400822 258054
rect 400586 257498 400822 257734
rect 400586 221818 400822 222054
rect 400586 221498 400822 221734
rect 400586 185818 400822 186054
rect 400586 185498 400822 185734
rect 400586 149818 400822 150054
rect 400586 149498 400822 149734
rect 400586 113818 400822 114054
rect 400586 113498 400822 113734
rect 400586 77818 400822 78054
rect 400586 77498 400822 77734
rect 400586 41818 400822 42054
rect 400586 41498 400822 41734
rect 400586 5818 400822 6054
rect 400586 5498 400822 5734
rect 400586 -2422 400822 -2186
rect 400586 -2742 400822 -2506
rect 404186 693418 404422 693654
rect 404186 693098 404422 693334
rect 404186 657418 404422 657654
rect 404186 657098 404422 657334
rect 404186 621418 404422 621654
rect 404186 621098 404422 621334
rect 404186 585418 404422 585654
rect 404186 585098 404422 585334
rect 404186 549418 404422 549654
rect 404186 549098 404422 549334
rect 404186 513418 404422 513654
rect 404186 513098 404422 513334
rect 404186 477418 404422 477654
rect 404186 477098 404422 477334
rect 404186 441418 404422 441654
rect 404186 441098 404422 441334
rect 404186 405418 404422 405654
rect 404186 405098 404422 405334
rect 404186 369418 404422 369654
rect 404186 369098 404422 369334
rect 404186 333418 404422 333654
rect 404186 333098 404422 333334
rect 404186 297418 404422 297654
rect 404186 297098 404422 297334
rect 404186 261418 404422 261654
rect 404186 261098 404422 261334
rect 404186 225418 404422 225654
rect 404186 225098 404422 225334
rect 404186 189418 404422 189654
rect 404186 189098 404422 189334
rect 404186 153418 404422 153654
rect 404186 153098 404422 153334
rect 404186 117418 404422 117654
rect 404186 117098 404422 117334
rect 404186 81418 404422 81654
rect 404186 81098 404422 81334
rect 404186 45418 404422 45654
rect 404186 45098 404422 45334
rect 404186 9418 404422 9654
rect 404186 9098 404422 9334
rect 404186 -4262 404422 -4026
rect 404186 -4582 404422 -4346
rect 425786 711042 426022 711278
rect 425786 710722 426022 710958
rect 422186 709202 422422 709438
rect 422186 708882 422422 709118
rect 418586 707362 418822 707598
rect 418586 707042 418822 707278
rect 407786 697018 408022 697254
rect 407786 696698 408022 696934
rect 407786 661018 408022 661254
rect 407786 660698 408022 660934
rect 407786 625018 408022 625254
rect 407786 624698 408022 624934
rect 407786 589018 408022 589254
rect 407786 588698 408022 588934
rect 407786 553018 408022 553254
rect 407786 552698 408022 552934
rect 407786 517018 408022 517254
rect 407786 516698 408022 516934
rect 407786 481018 408022 481254
rect 407786 480698 408022 480934
rect 407786 445018 408022 445254
rect 407786 444698 408022 444934
rect 407786 409018 408022 409254
rect 407786 408698 408022 408934
rect 407786 373018 408022 373254
rect 407786 372698 408022 372934
rect 407786 337018 408022 337254
rect 407786 336698 408022 336934
rect 407786 301018 408022 301254
rect 407786 300698 408022 300934
rect 407786 265018 408022 265254
rect 407786 264698 408022 264934
rect 407786 229018 408022 229254
rect 407786 228698 408022 228934
rect 407786 193018 408022 193254
rect 407786 192698 408022 192934
rect 407786 157018 408022 157254
rect 407786 156698 408022 156934
rect 407786 121018 408022 121254
rect 407786 120698 408022 120934
rect 407786 85018 408022 85254
rect 407786 84698 408022 84934
rect 407786 49018 408022 49254
rect 407786 48698 408022 48934
rect 407786 13018 408022 13254
rect 407786 12698 408022 12934
rect 389786 -7022 390022 -6786
rect 389786 -7342 390022 -7106
rect 414986 705522 415222 705758
rect 414986 705202 415222 705438
rect 414986 668218 415222 668454
rect 414986 667898 415222 668134
rect 414986 632218 415222 632454
rect 414986 631898 415222 632134
rect 414986 596218 415222 596454
rect 414986 595898 415222 596134
rect 414986 560218 415222 560454
rect 414986 559898 415222 560134
rect 414986 524218 415222 524454
rect 414986 523898 415222 524134
rect 414986 488218 415222 488454
rect 414986 487898 415222 488134
rect 414986 452218 415222 452454
rect 414986 451898 415222 452134
rect 414986 416218 415222 416454
rect 414986 415898 415222 416134
rect 414986 380218 415222 380454
rect 414986 379898 415222 380134
rect 414986 344218 415222 344454
rect 414986 343898 415222 344134
rect 414986 308218 415222 308454
rect 414986 307898 415222 308134
rect 414986 272218 415222 272454
rect 414986 271898 415222 272134
rect 414986 236218 415222 236454
rect 414986 235898 415222 236134
rect 414986 200218 415222 200454
rect 414986 199898 415222 200134
rect 414986 164218 415222 164454
rect 414986 163898 415222 164134
rect 414986 128218 415222 128454
rect 414986 127898 415222 128134
rect 414986 92218 415222 92454
rect 414986 91898 415222 92134
rect 414986 56218 415222 56454
rect 414986 55898 415222 56134
rect 414986 20218 415222 20454
rect 414986 19898 415222 20134
rect 414986 -1502 415222 -1266
rect 414986 -1822 415222 -1586
rect 418586 671818 418822 672054
rect 418586 671498 418822 671734
rect 418586 635818 418822 636054
rect 418586 635498 418822 635734
rect 418586 599818 418822 600054
rect 418586 599498 418822 599734
rect 418586 563818 418822 564054
rect 418586 563498 418822 563734
rect 418586 527818 418822 528054
rect 418586 527498 418822 527734
rect 418586 491818 418822 492054
rect 418586 491498 418822 491734
rect 418586 455818 418822 456054
rect 418586 455498 418822 455734
rect 418586 419818 418822 420054
rect 418586 419498 418822 419734
rect 418586 383818 418822 384054
rect 418586 383498 418822 383734
rect 418586 347818 418822 348054
rect 418586 347498 418822 347734
rect 418586 311818 418822 312054
rect 418586 311498 418822 311734
rect 418586 275818 418822 276054
rect 418586 275498 418822 275734
rect 418586 239818 418822 240054
rect 418586 239498 418822 239734
rect 418586 203818 418822 204054
rect 418586 203498 418822 203734
rect 418586 167818 418822 168054
rect 418586 167498 418822 167734
rect 418586 131818 418822 132054
rect 418586 131498 418822 131734
rect 418586 95818 418822 96054
rect 418586 95498 418822 95734
rect 418586 59818 418822 60054
rect 418586 59498 418822 59734
rect 418586 23818 418822 24054
rect 418586 23498 418822 23734
rect 418586 -3342 418822 -3106
rect 418586 -3662 418822 -3426
rect 422186 675418 422422 675654
rect 422186 675098 422422 675334
rect 422186 639418 422422 639654
rect 422186 639098 422422 639334
rect 422186 603418 422422 603654
rect 422186 603098 422422 603334
rect 422186 567418 422422 567654
rect 422186 567098 422422 567334
rect 422186 531418 422422 531654
rect 422186 531098 422422 531334
rect 422186 495418 422422 495654
rect 422186 495098 422422 495334
rect 422186 459418 422422 459654
rect 422186 459098 422422 459334
rect 422186 423418 422422 423654
rect 422186 423098 422422 423334
rect 422186 387418 422422 387654
rect 422186 387098 422422 387334
rect 422186 351418 422422 351654
rect 422186 351098 422422 351334
rect 422186 315418 422422 315654
rect 422186 315098 422422 315334
rect 422186 279418 422422 279654
rect 422186 279098 422422 279334
rect 422186 243418 422422 243654
rect 422186 243098 422422 243334
rect 422186 207418 422422 207654
rect 422186 207098 422422 207334
rect 422186 171418 422422 171654
rect 422186 171098 422422 171334
rect 422186 135418 422422 135654
rect 422186 135098 422422 135334
rect 422186 99418 422422 99654
rect 422186 99098 422422 99334
rect 422186 63418 422422 63654
rect 422186 63098 422422 63334
rect 422186 27418 422422 27654
rect 422186 27098 422422 27334
rect 422186 -5182 422422 -4946
rect 422186 -5502 422422 -5266
rect 443786 710122 444022 710358
rect 443786 709802 444022 710038
rect 440186 708282 440422 708518
rect 440186 707962 440422 708198
rect 436586 706442 436822 706678
rect 436586 706122 436822 706358
rect 425786 679018 426022 679254
rect 425786 678698 426022 678934
rect 425786 643018 426022 643254
rect 425786 642698 426022 642934
rect 425786 607018 426022 607254
rect 425786 606698 426022 606934
rect 425786 571018 426022 571254
rect 425786 570698 426022 570934
rect 425786 535018 426022 535254
rect 425786 534698 426022 534934
rect 425786 499018 426022 499254
rect 425786 498698 426022 498934
rect 425786 463018 426022 463254
rect 425786 462698 426022 462934
rect 425786 427018 426022 427254
rect 425786 426698 426022 426934
rect 425786 391018 426022 391254
rect 425786 390698 426022 390934
rect 425786 355018 426022 355254
rect 425786 354698 426022 354934
rect 425786 319018 426022 319254
rect 425786 318698 426022 318934
rect 425786 283018 426022 283254
rect 425786 282698 426022 282934
rect 425786 247018 426022 247254
rect 425786 246698 426022 246934
rect 425786 211018 426022 211254
rect 425786 210698 426022 210934
rect 425786 175018 426022 175254
rect 425786 174698 426022 174934
rect 425786 139018 426022 139254
rect 425786 138698 426022 138934
rect 425786 103018 426022 103254
rect 425786 102698 426022 102934
rect 425786 67018 426022 67254
rect 425786 66698 426022 66934
rect 425786 31018 426022 31254
rect 425786 30698 426022 30934
rect 407786 -6102 408022 -5866
rect 407786 -6422 408022 -6186
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 432986 686218 433222 686454
rect 432986 685898 433222 686134
rect 432986 650218 433222 650454
rect 432986 649898 433222 650134
rect 432986 614218 433222 614454
rect 432986 613898 433222 614134
rect 432986 578218 433222 578454
rect 432986 577898 433222 578134
rect 432986 542218 433222 542454
rect 432986 541898 433222 542134
rect 432986 506218 433222 506454
rect 432986 505898 433222 506134
rect 432986 470218 433222 470454
rect 432986 469898 433222 470134
rect 432986 434218 433222 434454
rect 432986 433898 433222 434134
rect 432986 398218 433222 398454
rect 432986 397898 433222 398134
rect 432986 362218 433222 362454
rect 432986 361898 433222 362134
rect 432986 326218 433222 326454
rect 432986 325898 433222 326134
rect 432986 290218 433222 290454
rect 432986 289898 433222 290134
rect 432986 254218 433222 254454
rect 432986 253898 433222 254134
rect 432986 218218 433222 218454
rect 432986 217898 433222 218134
rect 432986 182218 433222 182454
rect 432986 181898 433222 182134
rect 432986 146218 433222 146454
rect 432986 145898 433222 146134
rect 432986 110218 433222 110454
rect 432986 109898 433222 110134
rect 432986 74218 433222 74454
rect 432986 73898 433222 74134
rect 432986 38218 433222 38454
rect 432986 37898 433222 38134
rect 432986 2218 433222 2454
rect 432986 1898 433222 2134
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 436586 689818 436822 690054
rect 436586 689498 436822 689734
rect 436586 653818 436822 654054
rect 436586 653498 436822 653734
rect 436586 617818 436822 618054
rect 436586 617498 436822 617734
rect 436586 581818 436822 582054
rect 436586 581498 436822 581734
rect 436586 545818 436822 546054
rect 436586 545498 436822 545734
rect 436586 509818 436822 510054
rect 436586 509498 436822 509734
rect 436586 473818 436822 474054
rect 436586 473498 436822 473734
rect 436586 437818 436822 438054
rect 436586 437498 436822 437734
rect 436586 401818 436822 402054
rect 436586 401498 436822 401734
rect 436586 365818 436822 366054
rect 436586 365498 436822 365734
rect 436586 329818 436822 330054
rect 436586 329498 436822 329734
rect 436586 293818 436822 294054
rect 436586 293498 436822 293734
rect 436586 257818 436822 258054
rect 436586 257498 436822 257734
rect 436586 221818 436822 222054
rect 436586 221498 436822 221734
rect 436586 185818 436822 186054
rect 436586 185498 436822 185734
rect 436586 149818 436822 150054
rect 436586 149498 436822 149734
rect 436586 113818 436822 114054
rect 436586 113498 436822 113734
rect 436586 77818 436822 78054
rect 436586 77498 436822 77734
rect 436586 41818 436822 42054
rect 436586 41498 436822 41734
rect 436586 5818 436822 6054
rect 436586 5498 436822 5734
rect 436586 -2422 436822 -2186
rect 436586 -2742 436822 -2506
rect 440186 693418 440422 693654
rect 440186 693098 440422 693334
rect 440186 657418 440422 657654
rect 440186 657098 440422 657334
rect 440186 621418 440422 621654
rect 440186 621098 440422 621334
rect 440186 585418 440422 585654
rect 440186 585098 440422 585334
rect 440186 549418 440422 549654
rect 440186 549098 440422 549334
rect 440186 513418 440422 513654
rect 440186 513098 440422 513334
rect 440186 477418 440422 477654
rect 440186 477098 440422 477334
rect 440186 441418 440422 441654
rect 440186 441098 440422 441334
rect 440186 405418 440422 405654
rect 440186 405098 440422 405334
rect 440186 369418 440422 369654
rect 440186 369098 440422 369334
rect 440186 333418 440422 333654
rect 440186 333098 440422 333334
rect 440186 297418 440422 297654
rect 440186 297098 440422 297334
rect 440186 261418 440422 261654
rect 440186 261098 440422 261334
rect 440186 225418 440422 225654
rect 440186 225098 440422 225334
rect 440186 189418 440422 189654
rect 440186 189098 440422 189334
rect 440186 153418 440422 153654
rect 440186 153098 440422 153334
rect 440186 117418 440422 117654
rect 440186 117098 440422 117334
rect 440186 81418 440422 81654
rect 440186 81098 440422 81334
rect 440186 45418 440422 45654
rect 440186 45098 440422 45334
rect 440186 9418 440422 9654
rect 440186 9098 440422 9334
rect 440186 -4262 440422 -4026
rect 440186 -4582 440422 -4346
rect 461786 711042 462022 711278
rect 461786 710722 462022 710958
rect 458186 709202 458422 709438
rect 458186 708882 458422 709118
rect 454586 707362 454822 707598
rect 454586 707042 454822 707278
rect 443786 697018 444022 697254
rect 443786 696698 444022 696934
rect 443786 661018 444022 661254
rect 443786 660698 444022 660934
rect 443786 625018 444022 625254
rect 443786 624698 444022 624934
rect 443786 589018 444022 589254
rect 443786 588698 444022 588934
rect 443786 553018 444022 553254
rect 443786 552698 444022 552934
rect 443786 517018 444022 517254
rect 443786 516698 444022 516934
rect 443786 481018 444022 481254
rect 443786 480698 444022 480934
rect 443786 445018 444022 445254
rect 443786 444698 444022 444934
rect 443786 409018 444022 409254
rect 443786 408698 444022 408934
rect 443786 373018 444022 373254
rect 443786 372698 444022 372934
rect 443786 337018 444022 337254
rect 443786 336698 444022 336934
rect 443786 301018 444022 301254
rect 443786 300698 444022 300934
rect 443786 265018 444022 265254
rect 443786 264698 444022 264934
rect 443786 229018 444022 229254
rect 443786 228698 444022 228934
rect 443786 193018 444022 193254
rect 443786 192698 444022 192934
rect 443786 157018 444022 157254
rect 443786 156698 444022 156934
rect 443786 121018 444022 121254
rect 443786 120698 444022 120934
rect 443786 85018 444022 85254
rect 443786 84698 444022 84934
rect 443786 49018 444022 49254
rect 443786 48698 444022 48934
rect 443786 13018 444022 13254
rect 443786 12698 444022 12934
rect 425786 -7022 426022 -6786
rect 425786 -7342 426022 -7106
rect 450986 705522 451222 705758
rect 450986 705202 451222 705438
rect 450986 668218 451222 668454
rect 450986 667898 451222 668134
rect 450986 632218 451222 632454
rect 450986 631898 451222 632134
rect 450986 596218 451222 596454
rect 450986 595898 451222 596134
rect 450986 560218 451222 560454
rect 450986 559898 451222 560134
rect 450986 524218 451222 524454
rect 450986 523898 451222 524134
rect 450986 488218 451222 488454
rect 450986 487898 451222 488134
rect 450986 452218 451222 452454
rect 450986 451898 451222 452134
rect 450986 416218 451222 416454
rect 450986 415898 451222 416134
rect 450986 380218 451222 380454
rect 450986 379898 451222 380134
rect 450986 344218 451222 344454
rect 450986 343898 451222 344134
rect 450986 308218 451222 308454
rect 450986 307898 451222 308134
rect 450986 272218 451222 272454
rect 450986 271898 451222 272134
rect 450986 236218 451222 236454
rect 450986 235898 451222 236134
rect 450986 200218 451222 200454
rect 450986 199898 451222 200134
rect 450986 164218 451222 164454
rect 450986 163898 451222 164134
rect 450986 128218 451222 128454
rect 450986 127898 451222 128134
rect 450986 92218 451222 92454
rect 450986 91898 451222 92134
rect 450986 56218 451222 56454
rect 450986 55898 451222 56134
rect 450986 20218 451222 20454
rect 450986 19898 451222 20134
rect 450986 -1502 451222 -1266
rect 450986 -1822 451222 -1586
rect 454586 671818 454822 672054
rect 454586 671498 454822 671734
rect 454586 635818 454822 636054
rect 454586 635498 454822 635734
rect 454586 599818 454822 600054
rect 454586 599498 454822 599734
rect 454586 563818 454822 564054
rect 454586 563498 454822 563734
rect 454586 527818 454822 528054
rect 454586 527498 454822 527734
rect 454586 491818 454822 492054
rect 454586 491498 454822 491734
rect 454586 455818 454822 456054
rect 454586 455498 454822 455734
rect 454586 419818 454822 420054
rect 454586 419498 454822 419734
rect 454586 383818 454822 384054
rect 454586 383498 454822 383734
rect 454586 347818 454822 348054
rect 454586 347498 454822 347734
rect 454586 311818 454822 312054
rect 454586 311498 454822 311734
rect 454586 275818 454822 276054
rect 454586 275498 454822 275734
rect 454586 239818 454822 240054
rect 454586 239498 454822 239734
rect 454586 203818 454822 204054
rect 454586 203498 454822 203734
rect 454586 167818 454822 168054
rect 454586 167498 454822 167734
rect 454586 131818 454822 132054
rect 454586 131498 454822 131734
rect 454586 95818 454822 96054
rect 454586 95498 454822 95734
rect 454586 59818 454822 60054
rect 454586 59498 454822 59734
rect 454586 23818 454822 24054
rect 454586 23498 454822 23734
rect 454586 -3342 454822 -3106
rect 454586 -3662 454822 -3426
rect 458186 675418 458422 675654
rect 458186 675098 458422 675334
rect 458186 639418 458422 639654
rect 458186 639098 458422 639334
rect 458186 603418 458422 603654
rect 458186 603098 458422 603334
rect 458186 567418 458422 567654
rect 458186 567098 458422 567334
rect 458186 531418 458422 531654
rect 458186 531098 458422 531334
rect 458186 495418 458422 495654
rect 458186 495098 458422 495334
rect 458186 459418 458422 459654
rect 458186 459098 458422 459334
rect 458186 423418 458422 423654
rect 458186 423098 458422 423334
rect 458186 387418 458422 387654
rect 458186 387098 458422 387334
rect 458186 351418 458422 351654
rect 458186 351098 458422 351334
rect 458186 315418 458422 315654
rect 458186 315098 458422 315334
rect 458186 279418 458422 279654
rect 458186 279098 458422 279334
rect 458186 243418 458422 243654
rect 458186 243098 458422 243334
rect 458186 207418 458422 207654
rect 458186 207098 458422 207334
rect 458186 171418 458422 171654
rect 458186 171098 458422 171334
rect 458186 135418 458422 135654
rect 458186 135098 458422 135334
rect 458186 99418 458422 99654
rect 458186 99098 458422 99334
rect 458186 63418 458422 63654
rect 458186 63098 458422 63334
rect 458186 27418 458422 27654
rect 458186 27098 458422 27334
rect 458186 -5182 458422 -4946
rect 458186 -5502 458422 -5266
rect 479786 710122 480022 710358
rect 479786 709802 480022 710038
rect 476186 708282 476422 708518
rect 476186 707962 476422 708198
rect 472586 706442 472822 706678
rect 472586 706122 472822 706358
rect 461786 679018 462022 679254
rect 461786 678698 462022 678934
rect 461786 643018 462022 643254
rect 461786 642698 462022 642934
rect 461786 607018 462022 607254
rect 461786 606698 462022 606934
rect 461786 571018 462022 571254
rect 461786 570698 462022 570934
rect 461786 535018 462022 535254
rect 461786 534698 462022 534934
rect 461786 499018 462022 499254
rect 461786 498698 462022 498934
rect 461786 463018 462022 463254
rect 461786 462698 462022 462934
rect 461786 427018 462022 427254
rect 461786 426698 462022 426934
rect 461786 391018 462022 391254
rect 461786 390698 462022 390934
rect 461786 355018 462022 355254
rect 461786 354698 462022 354934
rect 461786 319018 462022 319254
rect 461786 318698 462022 318934
rect 461786 283018 462022 283254
rect 461786 282698 462022 282934
rect 461786 247018 462022 247254
rect 461786 246698 462022 246934
rect 461786 211018 462022 211254
rect 461786 210698 462022 210934
rect 461786 175018 462022 175254
rect 461786 174698 462022 174934
rect 461786 139018 462022 139254
rect 461786 138698 462022 138934
rect 461786 103018 462022 103254
rect 461786 102698 462022 102934
rect 461786 67018 462022 67254
rect 461786 66698 462022 66934
rect 461786 31018 462022 31254
rect 461786 30698 462022 30934
rect 443786 -6102 444022 -5866
rect 443786 -6422 444022 -6186
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 468986 686218 469222 686454
rect 468986 685898 469222 686134
rect 468986 650218 469222 650454
rect 468986 649898 469222 650134
rect 468986 614218 469222 614454
rect 468986 613898 469222 614134
rect 468986 578218 469222 578454
rect 468986 577898 469222 578134
rect 468986 542218 469222 542454
rect 468986 541898 469222 542134
rect 468986 506218 469222 506454
rect 468986 505898 469222 506134
rect 468986 470218 469222 470454
rect 468986 469898 469222 470134
rect 468986 434218 469222 434454
rect 468986 433898 469222 434134
rect 468986 398218 469222 398454
rect 468986 397898 469222 398134
rect 468986 362218 469222 362454
rect 468986 361898 469222 362134
rect 468986 326218 469222 326454
rect 468986 325898 469222 326134
rect 468986 290218 469222 290454
rect 468986 289898 469222 290134
rect 468986 254218 469222 254454
rect 468986 253898 469222 254134
rect 468986 218218 469222 218454
rect 468986 217898 469222 218134
rect 468986 182218 469222 182454
rect 468986 181898 469222 182134
rect 468986 146218 469222 146454
rect 468986 145898 469222 146134
rect 468986 110218 469222 110454
rect 468986 109898 469222 110134
rect 468986 74218 469222 74454
rect 468986 73898 469222 74134
rect 468986 38218 469222 38454
rect 468986 37898 469222 38134
rect 468986 2218 469222 2454
rect 468986 1898 469222 2134
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 472586 689818 472822 690054
rect 472586 689498 472822 689734
rect 472586 653818 472822 654054
rect 472586 653498 472822 653734
rect 472586 617818 472822 618054
rect 472586 617498 472822 617734
rect 472586 581818 472822 582054
rect 472586 581498 472822 581734
rect 472586 545818 472822 546054
rect 472586 545498 472822 545734
rect 472586 509818 472822 510054
rect 472586 509498 472822 509734
rect 472586 473818 472822 474054
rect 472586 473498 472822 473734
rect 472586 437818 472822 438054
rect 472586 437498 472822 437734
rect 472586 401818 472822 402054
rect 472586 401498 472822 401734
rect 472586 365818 472822 366054
rect 472586 365498 472822 365734
rect 472586 329818 472822 330054
rect 472586 329498 472822 329734
rect 472586 293818 472822 294054
rect 472586 293498 472822 293734
rect 472586 257818 472822 258054
rect 472586 257498 472822 257734
rect 472586 221818 472822 222054
rect 472586 221498 472822 221734
rect 472586 185818 472822 186054
rect 472586 185498 472822 185734
rect 472586 149818 472822 150054
rect 472586 149498 472822 149734
rect 472586 113818 472822 114054
rect 472586 113498 472822 113734
rect 472586 77818 472822 78054
rect 472586 77498 472822 77734
rect 472586 41818 472822 42054
rect 472586 41498 472822 41734
rect 472586 5818 472822 6054
rect 472586 5498 472822 5734
rect 472586 -2422 472822 -2186
rect 472586 -2742 472822 -2506
rect 476186 693418 476422 693654
rect 476186 693098 476422 693334
rect 476186 657418 476422 657654
rect 476186 657098 476422 657334
rect 476186 621418 476422 621654
rect 476186 621098 476422 621334
rect 476186 585418 476422 585654
rect 476186 585098 476422 585334
rect 476186 549418 476422 549654
rect 476186 549098 476422 549334
rect 476186 513418 476422 513654
rect 476186 513098 476422 513334
rect 476186 477418 476422 477654
rect 476186 477098 476422 477334
rect 476186 441418 476422 441654
rect 476186 441098 476422 441334
rect 476186 405418 476422 405654
rect 476186 405098 476422 405334
rect 476186 369418 476422 369654
rect 476186 369098 476422 369334
rect 476186 333418 476422 333654
rect 476186 333098 476422 333334
rect 476186 297418 476422 297654
rect 476186 297098 476422 297334
rect 476186 261418 476422 261654
rect 476186 261098 476422 261334
rect 476186 225418 476422 225654
rect 476186 225098 476422 225334
rect 476186 189418 476422 189654
rect 476186 189098 476422 189334
rect 476186 153418 476422 153654
rect 476186 153098 476422 153334
rect 476186 117418 476422 117654
rect 476186 117098 476422 117334
rect 476186 81418 476422 81654
rect 476186 81098 476422 81334
rect 476186 45418 476422 45654
rect 476186 45098 476422 45334
rect 476186 9418 476422 9654
rect 476186 9098 476422 9334
rect 476186 -4262 476422 -4026
rect 476186 -4582 476422 -4346
rect 497786 711042 498022 711278
rect 497786 710722 498022 710958
rect 494186 709202 494422 709438
rect 494186 708882 494422 709118
rect 490586 707362 490822 707598
rect 490586 707042 490822 707278
rect 479786 697018 480022 697254
rect 479786 696698 480022 696934
rect 479786 661018 480022 661254
rect 479786 660698 480022 660934
rect 479786 625018 480022 625254
rect 479786 624698 480022 624934
rect 479786 589018 480022 589254
rect 479786 588698 480022 588934
rect 479786 553018 480022 553254
rect 479786 552698 480022 552934
rect 479786 517018 480022 517254
rect 479786 516698 480022 516934
rect 479786 481018 480022 481254
rect 479786 480698 480022 480934
rect 479786 445018 480022 445254
rect 479786 444698 480022 444934
rect 479786 409018 480022 409254
rect 479786 408698 480022 408934
rect 479786 373018 480022 373254
rect 479786 372698 480022 372934
rect 479786 337018 480022 337254
rect 479786 336698 480022 336934
rect 479786 301018 480022 301254
rect 479786 300698 480022 300934
rect 479786 265018 480022 265254
rect 479786 264698 480022 264934
rect 479786 229018 480022 229254
rect 479786 228698 480022 228934
rect 479786 193018 480022 193254
rect 479786 192698 480022 192934
rect 479786 157018 480022 157254
rect 479786 156698 480022 156934
rect 479786 121018 480022 121254
rect 479786 120698 480022 120934
rect 479786 85018 480022 85254
rect 479786 84698 480022 84934
rect 479786 49018 480022 49254
rect 479786 48698 480022 48934
rect 479786 13018 480022 13254
rect 479786 12698 480022 12934
rect 461786 -7022 462022 -6786
rect 461786 -7342 462022 -7106
rect 486986 705522 487222 705758
rect 486986 705202 487222 705438
rect 486986 668218 487222 668454
rect 486986 667898 487222 668134
rect 486986 632218 487222 632454
rect 486986 631898 487222 632134
rect 486986 596218 487222 596454
rect 486986 595898 487222 596134
rect 486986 560218 487222 560454
rect 486986 559898 487222 560134
rect 486986 524218 487222 524454
rect 486986 523898 487222 524134
rect 486986 488218 487222 488454
rect 486986 487898 487222 488134
rect 486986 452218 487222 452454
rect 486986 451898 487222 452134
rect 486986 416218 487222 416454
rect 486986 415898 487222 416134
rect 486986 380218 487222 380454
rect 486986 379898 487222 380134
rect 486986 344218 487222 344454
rect 486986 343898 487222 344134
rect 486986 308218 487222 308454
rect 486986 307898 487222 308134
rect 486986 272218 487222 272454
rect 486986 271898 487222 272134
rect 486986 236218 487222 236454
rect 486986 235898 487222 236134
rect 486986 200218 487222 200454
rect 486986 199898 487222 200134
rect 486986 164218 487222 164454
rect 486986 163898 487222 164134
rect 486986 128218 487222 128454
rect 486986 127898 487222 128134
rect 486986 92218 487222 92454
rect 486986 91898 487222 92134
rect 486986 56218 487222 56454
rect 486986 55898 487222 56134
rect 486986 20218 487222 20454
rect 486986 19898 487222 20134
rect 486986 -1502 487222 -1266
rect 486986 -1822 487222 -1586
rect 490586 671818 490822 672054
rect 490586 671498 490822 671734
rect 490586 635818 490822 636054
rect 490586 635498 490822 635734
rect 490586 599818 490822 600054
rect 490586 599498 490822 599734
rect 490586 563818 490822 564054
rect 490586 563498 490822 563734
rect 490586 527818 490822 528054
rect 490586 527498 490822 527734
rect 490586 491818 490822 492054
rect 490586 491498 490822 491734
rect 490586 455818 490822 456054
rect 490586 455498 490822 455734
rect 490586 419818 490822 420054
rect 490586 419498 490822 419734
rect 490586 383818 490822 384054
rect 490586 383498 490822 383734
rect 490586 347818 490822 348054
rect 490586 347498 490822 347734
rect 490586 311818 490822 312054
rect 490586 311498 490822 311734
rect 490586 275818 490822 276054
rect 490586 275498 490822 275734
rect 490586 239818 490822 240054
rect 490586 239498 490822 239734
rect 490586 203818 490822 204054
rect 490586 203498 490822 203734
rect 490586 167818 490822 168054
rect 490586 167498 490822 167734
rect 490586 131818 490822 132054
rect 490586 131498 490822 131734
rect 490586 95818 490822 96054
rect 490586 95498 490822 95734
rect 490586 59818 490822 60054
rect 490586 59498 490822 59734
rect 490586 23818 490822 24054
rect 490586 23498 490822 23734
rect 490586 -3342 490822 -3106
rect 490586 -3662 490822 -3426
rect 494186 675418 494422 675654
rect 494186 675098 494422 675334
rect 494186 639418 494422 639654
rect 494186 639098 494422 639334
rect 494186 603418 494422 603654
rect 494186 603098 494422 603334
rect 494186 567418 494422 567654
rect 494186 567098 494422 567334
rect 494186 531418 494422 531654
rect 494186 531098 494422 531334
rect 494186 495418 494422 495654
rect 494186 495098 494422 495334
rect 494186 459418 494422 459654
rect 494186 459098 494422 459334
rect 494186 423418 494422 423654
rect 494186 423098 494422 423334
rect 494186 387418 494422 387654
rect 494186 387098 494422 387334
rect 494186 351418 494422 351654
rect 494186 351098 494422 351334
rect 494186 315418 494422 315654
rect 494186 315098 494422 315334
rect 494186 279418 494422 279654
rect 494186 279098 494422 279334
rect 494186 243418 494422 243654
rect 494186 243098 494422 243334
rect 494186 207418 494422 207654
rect 494186 207098 494422 207334
rect 494186 171418 494422 171654
rect 494186 171098 494422 171334
rect 494186 135418 494422 135654
rect 494186 135098 494422 135334
rect 494186 99418 494422 99654
rect 494186 99098 494422 99334
rect 494186 63418 494422 63654
rect 494186 63098 494422 63334
rect 494186 27418 494422 27654
rect 494186 27098 494422 27334
rect 494186 -5182 494422 -4946
rect 494186 -5502 494422 -5266
rect 515786 710122 516022 710358
rect 515786 709802 516022 710038
rect 512186 708282 512422 708518
rect 512186 707962 512422 708198
rect 508586 706442 508822 706678
rect 508586 706122 508822 706358
rect 497786 679018 498022 679254
rect 497786 678698 498022 678934
rect 497786 643018 498022 643254
rect 497786 642698 498022 642934
rect 497786 607018 498022 607254
rect 497786 606698 498022 606934
rect 497786 571018 498022 571254
rect 497786 570698 498022 570934
rect 497786 535018 498022 535254
rect 497786 534698 498022 534934
rect 497786 499018 498022 499254
rect 497786 498698 498022 498934
rect 497786 463018 498022 463254
rect 497786 462698 498022 462934
rect 497786 427018 498022 427254
rect 497786 426698 498022 426934
rect 497786 391018 498022 391254
rect 497786 390698 498022 390934
rect 497786 355018 498022 355254
rect 497786 354698 498022 354934
rect 497786 319018 498022 319254
rect 497786 318698 498022 318934
rect 497786 283018 498022 283254
rect 497786 282698 498022 282934
rect 497786 247018 498022 247254
rect 497786 246698 498022 246934
rect 497786 211018 498022 211254
rect 497786 210698 498022 210934
rect 497786 175018 498022 175254
rect 497786 174698 498022 174934
rect 497786 139018 498022 139254
rect 497786 138698 498022 138934
rect 497786 103018 498022 103254
rect 497786 102698 498022 102934
rect 497786 67018 498022 67254
rect 497786 66698 498022 66934
rect 497786 31018 498022 31254
rect 497786 30698 498022 30934
rect 479786 -6102 480022 -5866
rect 479786 -6422 480022 -6186
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 504986 686218 505222 686454
rect 504986 685898 505222 686134
rect 504986 650218 505222 650454
rect 504986 649898 505222 650134
rect 504986 614218 505222 614454
rect 504986 613898 505222 614134
rect 504986 578218 505222 578454
rect 504986 577898 505222 578134
rect 504986 542218 505222 542454
rect 504986 541898 505222 542134
rect 504986 506218 505222 506454
rect 504986 505898 505222 506134
rect 504986 470218 505222 470454
rect 504986 469898 505222 470134
rect 504986 434218 505222 434454
rect 504986 433898 505222 434134
rect 504986 398218 505222 398454
rect 504986 397898 505222 398134
rect 504986 362218 505222 362454
rect 504986 361898 505222 362134
rect 504986 326218 505222 326454
rect 504986 325898 505222 326134
rect 504986 290218 505222 290454
rect 504986 289898 505222 290134
rect 504986 254218 505222 254454
rect 504986 253898 505222 254134
rect 504986 218218 505222 218454
rect 504986 217898 505222 218134
rect 504986 182218 505222 182454
rect 504986 181898 505222 182134
rect 504986 146218 505222 146454
rect 504986 145898 505222 146134
rect 504986 110218 505222 110454
rect 504986 109898 505222 110134
rect 504986 74218 505222 74454
rect 504986 73898 505222 74134
rect 504986 38218 505222 38454
rect 504986 37898 505222 38134
rect 504986 2218 505222 2454
rect 504986 1898 505222 2134
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 508586 689818 508822 690054
rect 508586 689498 508822 689734
rect 508586 653818 508822 654054
rect 508586 653498 508822 653734
rect 508586 617818 508822 618054
rect 508586 617498 508822 617734
rect 508586 581818 508822 582054
rect 508586 581498 508822 581734
rect 508586 545818 508822 546054
rect 508586 545498 508822 545734
rect 508586 509818 508822 510054
rect 508586 509498 508822 509734
rect 508586 473818 508822 474054
rect 508586 473498 508822 473734
rect 508586 437818 508822 438054
rect 508586 437498 508822 437734
rect 508586 401818 508822 402054
rect 508586 401498 508822 401734
rect 508586 365818 508822 366054
rect 508586 365498 508822 365734
rect 508586 329818 508822 330054
rect 508586 329498 508822 329734
rect 508586 293818 508822 294054
rect 508586 293498 508822 293734
rect 508586 257818 508822 258054
rect 508586 257498 508822 257734
rect 508586 221818 508822 222054
rect 508586 221498 508822 221734
rect 508586 185818 508822 186054
rect 508586 185498 508822 185734
rect 508586 149818 508822 150054
rect 508586 149498 508822 149734
rect 508586 113818 508822 114054
rect 508586 113498 508822 113734
rect 508586 77818 508822 78054
rect 508586 77498 508822 77734
rect 508586 41818 508822 42054
rect 508586 41498 508822 41734
rect 508586 5818 508822 6054
rect 508586 5498 508822 5734
rect 508586 -2422 508822 -2186
rect 508586 -2742 508822 -2506
rect 512186 693418 512422 693654
rect 512186 693098 512422 693334
rect 512186 657418 512422 657654
rect 512186 657098 512422 657334
rect 512186 621418 512422 621654
rect 512186 621098 512422 621334
rect 512186 585418 512422 585654
rect 512186 585098 512422 585334
rect 512186 549418 512422 549654
rect 512186 549098 512422 549334
rect 512186 513418 512422 513654
rect 512186 513098 512422 513334
rect 512186 477418 512422 477654
rect 512186 477098 512422 477334
rect 512186 441418 512422 441654
rect 512186 441098 512422 441334
rect 512186 405418 512422 405654
rect 512186 405098 512422 405334
rect 512186 369418 512422 369654
rect 512186 369098 512422 369334
rect 512186 333418 512422 333654
rect 512186 333098 512422 333334
rect 512186 297418 512422 297654
rect 512186 297098 512422 297334
rect 512186 261418 512422 261654
rect 512186 261098 512422 261334
rect 512186 225418 512422 225654
rect 512186 225098 512422 225334
rect 512186 189418 512422 189654
rect 512186 189098 512422 189334
rect 512186 153418 512422 153654
rect 512186 153098 512422 153334
rect 512186 117418 512422 117654
rect 512186 117098 512422 117334
rect 512186 81418 512422 81654
rect 512186 81098 512422 81334
rect 512186 45418 512422 45654
rect 512186 45098 512422 45334
rect 512186 9418 512422 9654
rect 512186 9098 512422 9334
rect 512186 -4262 512422 -4026
rect 512186 -4582 512422 -4346
rect 533786 711042 534022 711278
rect 533786 710722 534022 710958
rect 530186 709202 530422 709438
rect 530186 708882 530422 709118
rect 526586 707362 526822 707598
rect 526586 707042 526822 707278
rect 515786 697018 516022 697254
rect 515786 696698 516022 696934
rect 515786 661018 516022 661254
rect 515786 660698 516022 660934
rect 515786 625018 516022 625254
rect 515786 624698 516022 624934
rect 515786 589018 516022 589254
rect 515786 588698 516022 588934
rect 515786 553018 516022 553254
rect 515786 552698 516022 552934
rect 515786 517018 516022 517254
rect 515786 516698 516022 516934
rect 515786 481018 516022 481254
rect 515786 480698 516022 480934
rect 515786 445018 516022 445254
rect 515786 444698 516022 444934
rect 515786 409018 516022 409254
rect 515786 408698 516022 408934
rect 515786 373018 516022 373254
rect 515786 372698 516022 372934
rect 515786 337018 516022 337254
rect 515786 336698 516022 336934
rect 515786 301018 516022 301254
rect 515786 300698 516022 300934
rect 515786 265018 516022 265254
rect 515786 264698 516022 264934
rect 515786 229018 516022 229254
rect 515786 228698 516022 228934
rect 515786 193018 516022 193254
rect 515786 192698 516022 192934
rect 515786 157018 516022 157254
rect 515786 156698 516022 156934
rect 515786 121018 516022 121254
rect 515786 120698 516022 120934
rect 515786 85018 516022 85254
rect 515786 84698 516022 84934
rect 515786 49018 516022 49254
rect 515786 48698 516022 48934
rect 515786 13018 516022 13254
rect 515786 12698 516022 12934
rect 497786 -7022 498022 -6786
rect 497786 -7342 498022 -7106
rect 522986 705522 523222 705758
rect 522986 705202 523222 705438
rect 522986 668218 523222 668454
rect 522986 667898 523222 668134
rect 522986 632218 523222 632454
rect 522986 631898 523222 632134
rect 522986 596218 523222 596454
rect 522986 595898 523222 596134
rect 522986 560218 523222 560454
rect 522986 559898 523222 560134
rect 522986 524218 523222 524454
rect 522986 523898 523222 524134
rect 522986 488218 523222 488454
rect 522986 487898 523222 488134
rect 522986 452218 523222 452454
rect 522986 451898 523222 452134
rect 522986 416218 523222 416454
rect 522986 415898 523222 416134
rect 522986 380218 523222 380454
rect 522986 379898 523222 380134
rect 522986 344218 523222 344454
rect 522986 343898 523222 344134
rect 522986 308218 523222 308454
rect 522986 307898 523222 308134
rect 522986 272218 523222 272454
rect 522986 271898 523222 272134
rect 522986 236218 523222 236454
rect 522986 235898 523222 236134
rect 522986 200218 523222 200454
rect 522986 199898 523222 200134
rect 522986 164218 523222 164454
rect 522986 163898 523222 164134
rect 522986 128218 523222 128454
rect 522986 127898 523222 128134
rect 522986 92218 523222 92454
rect 522986 91898 523222 92134
rect 522986 56218 523222 56454
rect 522986 55898 523222 56134
rect 522986 20218 523222 20454
rect 522986 19898 523222 20134
rect 522986 -1502 523222 -1266
rect 522986 -1822 523222 -1586
rect 526586 671818 526822 672054
rect 526586 671498 526822 671734
rect 526586 635818 526822 636054
rect 526586 635498 526822 635734
rect 526586 599818 526822 600054
rect 526586 599498 526822 599734
rect 526586 563818 526822 564054
rect 526586 563498 526822 563734
rect 526586 527818 526822 528054
rect 526586 527498 526822 527734
rect 526586 491818 526822 492054
rect 526586 491498 526822 491734
rect 526586 455818 526822 456054
rect 526586 455498 526822 455734
rect 526586 419818 526822 420054
rect 526586 419498 526822 419734
rect 526586 383818 526822 384054
rect 526586 383498 526822 383734
rect 526586 347818 526822 348054
rect 526586 347498 526822 347734
rect 526586 311818 526822 312054
rect 526586 311498 526822 311734
rect 526586 275818 526822 276054
rect 526586 275498 526822 275734
rect 526586 239818 526822 240054
rect 526586 239498 526822 239734
rect 526586 203818 526822 204054
rect 526586 203498 526822 203734
rect 526586 167818 526822 168054
rect 526586 167498 526822 167734
rect 526586 131818 526822 132054
rect 526586 131498 526822 131734
rect 526586 95818 526822 96054
rect 526586 95498 526822 95734
rect 526586 59818 526822 60054
rect 526586 59498 526822 59734
rect 526586 23818 526822 24054
rect 526586 23498 526822 23734
rect 526586 -3342 526822 -3106
rect 526586 -3662 526822 -3426
rect 530186 675418 530422 675654
rect 530186 675098 530422 675334
rect 530186 639418 530422 639654
rect 530186 639098 530422 639334
rect 530186 603418 530422 603654
rect 530186 603098 530422 603334
rect 530186 567418 530422 567654
rect 530186 567098 530422 567334
rect 530186 531418 530422 531654
rect 530186 531098 530422 531334
rect 530186 495418 530422 495654
rect 530186 495098 530422 495334
rect 530186 459418 530422 459654
rect 530186 459098 530422 459334
rect 530186 423418 530422 423654
rect 530186 423098 530422 423334
rect 530186 387418 530422 387654
rect 530186 387098 530422 387334
rect 530186 351418 530422 351654
rect 530186 351098 530422 351334
rect 530186 315418 530422 315654
rect 530186 315098 530422 315334
rect 530186 279418 530422 279654
rect 530186 279098 530422 279334
rect 530186 243418 530422 243654
rect 530186 243098 530422 243334
rect 530186 207418 530422 207654
rect 530186 207098 530422 207334
rect 530186 171418 530422 171654
rect 530186 171098 530422 171334
rect 530186 135418 530422 135654
rect 530186 135098 530422 135334
rect 530186 99418 530422 99654
rect 530186 99098 530422 99334
rect 530186 63418 530422 63654
rect 530186 63098 530422 63334
rect 530186 27418 530422 27654
rect 530186 27098 530422 27334
rect 530186 -5182 530422 -4946
rect 530186 -5502 530422 -5266
rect 551786 710122 552022 710358
rect 551786 709802 552022 710038
rect 548186 708282 548422 708518
rect 548186 707962 548422 708198
rect 544586 706442 544822 706678
rect 544586 706122 544822 706358
rect 533786 679018 534022 679254
rect 533786 678698 534022 678934
rect 533786 643018 534022 643254
rect 533786 642698 534022 642934
rect 533786 607018 534022 607254
rect 533786 606698 534022 606934
rect 533786 571018 534022 571254
rect 533786 570698 534022 570934
rect 533786 535018 534022 535254
rect 533786 534698 534022 534934
rect 533786 499018 534022 499254
rect 533786 498698 534022 498934
rect 533786 463018 534022 463254
rect 533786 462698 534022 462934
rect 533786 427018 534022 427254
rect 533786 426698 534022 426934
rect 533786 391018 534022 391254
rect 533786 390698 534022 390934
rect 533786 355018 534022 355254
rect 533786 354698 534022 354934
rect 533786 319018 534022 319254
rect 533786 318698 534022 318934
rect 533786 283018 534022 283254
rect 533786 282698 534022 282934
rect 533786 247018 534022 247254
rect 533786 246698 534022 246934
rect 533786 211018 534022 211254
rect 533786 210698 534022 210934
rect 533786 175018 534022 175254
rect 533786 174698 534022 174934
rect 533786 139018 534022 139254
rect 533786 138698 534022 138934
rect 533786 103018 534022 103254
rect 533786 102698 534022 102934
rect 533786 67018 534022 67254
rect 533786 66698 534022 66934
rect 533786 31018 534022 31254
rect 533786 30698 534022 30934
rect 515786 -6102 516022 -5866
rect 515786 -6422 516022 -6186
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 540986 686218 541222 686454
rect 540986 685898 541222 686134
rect 540986 650218 541222 650454
rect 540986 649898 541222 650134
rect 540986 614218 541222 614454
rect 540986 613898 541222 614134
rect 540986 578218 541222 578454
rect 540986 577898 541222 578134
rect 540986 542218 541222 542454
rect 540986 541898 541222 542134
rect 540986 506218 541222 506454
rect 540986 505898 541222 506134
rect 540986 470218 541222 470454
rect 540986 469898 541222 470134
rect 540986 434218 541222 434454
rect 540986 433898 541222 434134
rect 540986 398218 541222 398454
rect 540986 397898 541222 398134
rect 540986 362218 541222 362454
rect 540986 361898 541222 362134
rect 540986 326218 541222 326454
rect 540986 325898 541222 326134
rect 540986 290218 541222 290454
rect 540986 289898 541222 290134
rect 540986 254218 541222 254454
rect 540986 253898 541222 254134
rect 540986 218218 541222 218454
rect 540986 217898 541222 218134
rect 540986 182218 541222 182454
rect 540986 181898 541222 182134
rect 540986 146218 541222 146454
rect 540986 145898 541222 146134
rect 540986 110218 541222 110454
rect 540986 109898 541222 110134
rect 540986 74218 541222 74454
rect 540986 73898 541222 74134
rect 540986 38218 541222 38454
rect 540986 37898 541222 38134
rect 540986 2218 541222 2454
rect 540986 1898 541222 2134
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 544586 689818 544822 690054
rect 544586 689498 544822 689734
rect 544586 653818 544822 654054
rect 544586 653498 544822 653734
rect 544586 617818 544822 618054
rect 544586 617498 544822 617734
rect 544586 581818 544822 582054
rect 544586 581498 544822 581734
rect 544586 545818 544822 546054
rect 544586 545498 544822 545734
rect 544586 509818 544822 510054
rect 544586 509498 544822 509734
rect 544586 473818 544822 474054
rect 544586 473498 544822 473734
rect 544586 437818 544822 438054
rect 544586 437498 544822 437734
rect 544586 401818 544822 402054
rect 544586 401498 544822 401734
rect 544586 365818 544822 366054
rect 544586 365498 544822 365734
rect 544586 329818 544822 330054
rect 544586 329498 544822 329734
rect 544586 293818 544822 294054
rect 544586 293498 544822 293734
rect 544586 257818 544822 258054
rect 544586 257498 544822 257734
rect 544586 221818 544822 222054
rect 544586 221498 544822 221734
rect 544586 185818 544822 186054
rect 544586 185498 544822 185734
rect 544586 149818 544822 150054
rect 544586 149498 544822 149734
rect 544586 113818 544822 114054
rect 544586 113498 544822 113734
rect 544586 77818 544822 78054
rect 544586 77498 544822 77734
rect 544586 41818 544822 42054
rect 544586 41498 544822 41734
rect 544586 5818 544822 6054
rect 544586 5498 544822 5734
rect 544586 -2422 544822 -2186
rect 544586 -2742 544822 -2506
rect 548186 693418 548422 693654
rect 548186 693098 548422 693334
rect 548186 657418 548422 657654
rect 548186 657098 548422 657334
rect 548186 621418 548422 621654
rect 548186 621098 548422 621334
rect 548186 585418 548422 585654
rect 548186 585098 548422 585334
rect 548186 549418 548422 549654
rect 548186 549098 548422 549334
rect 548186 513418 548422 513654
rect 548186 513098 548422 513334
rect 548186 477418 548422 477654
rect 548186 477098 548422 477334
rect 548186 441418 548422 441654
rect 548186 441098 548422 441334
rect 548186 405418 548422 405654
rect 548186 405098 548422 405334
rect 548186 369418 548422 369654
rect 548186 369098 548422 369334
rect 548186 333418 548422 333654
rect 548186 333098 548422 333334
rect 548186 297418 548422 297654
rect 548186 297098 548422 297334
rect 548186 261418 548422 261654
rect 548186 261098 548422 261334
rect 548186 225418 548422 225654
rect 548186 225098 548422 225334
rect 548186 189418 548422 189654
rect 548186 189098 548422 189334
rect 548186 153418 548422 153654
rect 548186 153098 548422 153334
rect 548186 117418 548422 117654
rect 548186 117098 548422 117334
rect 548186 81418 548422 81654
rect 548186 81098 548422 81334
rect 548186 45418 548422 45654
rect 548186 45098 548422 45334
rect 548186 9418 548422 9654
rect 548186 9098 548422 9334
rect 548186 -4262 548422 -4026
rect 548186 -4582 548422 -4346
rect 569786 711042 570022 711278
rect 569786 710722 570022 710958
rect 566186 709202 566422 709438
rect 566186 708882 566422 709118
rect 562586 707362 562822 707598
rect 562586 707042 562822 707278
rect 551786 697018 552022 697254
rect 551786 696698 552022 696934
rect 551786 661018 552022 661254
rect 551786 660698 552022 660934
rect 551786 625018 552022 625254
rect 551786 624698 552022 624934
rect 551786 589018 552022 589254
rect 551786 588698 552022 588934
rect 551786 553018 552022 553254
rect 551786 552698 552022 552934
rect 551786 517018 552022 517254
rect 551786 516698 552022 516934
rect 551786 481018 552022 481254
rect 551786 480698 552022 480934
rect 551786 445018 552022 445254
rect 551786 444698 552022 444934
rect 551786 409018 552022 409254
rect 551786 408698 552022 408934
rect 551786 373018 552022 373254
rect 551786 372698 552022 372934
rect 551786 337018 552022 337254
rect 551786 336698 552022 336934
rect 551786 301018 552022 301254
rect 551786 300698 552022 300934
rect 551786 265018 552022 265254
rect 551786 264698 552022 264934
rect 551786 229018 552022 229254
rect 551786 228698 552022 228934
rect 551786 193018 552022 193254
rect 551786 192698 552022 192934
rect 551786 157018 552022 157254
rect 551786 156698 552022 156934
rect 551786 121018 552022 121254
rect 551786 120698 552022 120934
rect 551786 85018 552022 85254
rect 551786 84698 552022 84934
rect 551786 49018 552022 49254
rect 551786 48698 552022 48934
rect 551786 13018 552022 13254
rect 551786 12698 552022 12934
rect 533786 -7022 534022 -6786
rect 533786 -7342 534022 -7106
rect 558986 705522 559222 705758
rect 558986 705202 559222 705438
rect 558986 668218 559222 668454
rect 558986 667898 559222 668134
rect 558986 632218 559222 632454
rect 558986 631898 559222 632134
rect 558986 596218 559222 596454
rect 558986 595898 559222 596134
rect 558986 560218 559222 560454
rect 558986 559898 559222 560134
rect 558986 524218 559222 524454
rect 558986 523898 559222 524134
rect 558986 488218 559222 488454
rect 558986 487898 559222 488134
rect 558986 452218 559222 452454
rect 558986 451898 559222 452134
rect 558986 416218 559222 416454
rect 558986 415898 559222 416134
rect 558986 380218 559222 380454
rect 558986 379898 559222 380134
rect 558986 344218 559222 344454
rect 558986 343898 559222 344134
rect 558986 308218 559222 308454
rect 558986 307898 559222 308134
rect 558986 272218 559222 272454
rect 558986 271898 559222 272134
rect 558986 236218 559222 236454
rect 558986 235898 559222 236134
rect 558986 200218 559222 200454
rect 558986 199898 559222 200134
rect 558986 164218 559222 164454
rect 558986 163898 559222 164134
rect 558986 128218 559222 128454
rect 558986 127898 559222 128134
rect 558986 92218 559222 92454
rect 558986 91898 559222 92134
rect 558986 56218 559222 56454
rect 558986 55898 559222 56134
rect 558986 20218 559222 20454
rect 558986 19898 559222 20134
rect 558986 -1502 559222 -1266
rect 558986 -1822 559222 -1586
rect 562586 671818 562822 672054
rect 562586 671498 562822 671734
rect 562586 635818 562822 636054
rect 562586 635498 562822 635734
rect 562586 599818 562822 600054
rect 562586 599498 562822 599734
rect 562586 563818 562822 564054
rect 562586 563498 562822 563734
rect 562586 527818 562822 528054
rect 562586 527498 562822 527734
rect 562586 491818 562822 492054
rect 562586 491498 562822 491734
rect 562586 455818 562822 456054
rect 562586 455498 562822 455734
rect 562586 419818 562822 420054
rect 562586 419498 562822 419734
rect 562586 383818 562822 384054
rect 562586 383498 562822 383734
rect 562586 347818 562822 348054
rect 562586 347498 562822 347734
rect 562586 311818 562822 312054
rect 562586 311498 562822 311734
rect 562586 275818 562822 276054
rect 562586 275498 562822 275734
rect 562586 239818 562822 240054
rect 562586 239498 562822 239734
rect 562586 203818 562822 204054
rect 562586 203498 562822 203734
rect 562586 167818 562822 168054
rect 562586 167498 562822 167734
rect 562586 131818 562822 132054
rect 562586 131498 562822 131734
rect 562586 95818 562822 96054
rect 562586 95498 562822 95734
rect 562586 59818 562822 60054
rect 562586 59498 562822 59734
rect 562586 23818 562822 24054
rect 562586 23498 562822 23734
rect 562586 -3342 562822 -3106
rect 562586 -3662 562822 -3426
rect 566186 675418 566422 675654
rect 566186 675098 566422 675334
rect 566186 639418 566422 639654
rect 566186 639098 566422 639334
rect 566186 603418 566422 603654
rect 566186 603098 566422 603334
rect 566186 567418 566422 567654
rect 566186 567098 566422 567334
rect 566186 531418 566422 531654
rect 566186 531098 566422 531334
rect 566186 495418 566422 495654
rect 566186 495098 566422 495334
rect 566186 459418 566422 459654
rect 566186 459098 566422 459334
rect 566186 423418 566422 423654
rect 566186 423098 566422 423334
rect 566186 387418 566422 387654
rect 566186 387098 566422 387334
rect 566186 351418 566422 351654
rect 566186 351098 566422 351334
rect 566186 315418 566422 315654
rect 566186 315098 566422 315334
rect 566186 279418 566422 279654
rect 566186 279098 566422 279334
rect 566186 243418 566422 243654
rect 566186 243098 566422 243334
rect 566186 207418 566422 207654
rect 566186 207098 566422 207334
rect 566186 171418 566422 171654
rect 566186 171098 566422 171334
rect 566186 135418 566422 135654
rect 566186 135098 566422 135334
rect 566186 99418 566422 99654
rect 566186 99098 566422 99334
rect 566186 63418 566422 63654
rect 566186 63098 566422 63334
rect 566186 27418 566422 27654
rect 566186 27098 566422 27334
rect 566186 -5182 566422 -4946
rect 566186 -5502 566422 -5266
rect 591942 711042 592178 711278
rect 591942 710722 592178 710958
rect 591022 710122 591258 710358
rect 591022 709802 591258 710038
rect 590102 709202 590338 709438
rect 590102 708882 590338 709118
rect 589182 708282 589418 708518
rect 589182 707962 589418 708198
rect 588262 707362 588498 707598
rect 588262 707042 588498 707278
rect 580586 706442 580822 706678
rect 580586 706122 580822 706358
rect 569786 679018 570022 679254
rect 569786 678698 570022 678934
rect 569786 643018 570022 643254
rect 569786 642698 570022 642934
rect 569786 607018 570022 607254
rect 569786 606698 570022 606934
rect 569786 571018 570022 571254
rect 569786 570698 570022 570934
rect 569786 535018 570022 535254
rect 569786 534698 570022 534934
rect 569786 499018 570022 499254
rect 569786 498698 570022 498934
rect 569786 463018 570022 463254
rect 569786 462698 570022 462934
rect 569786 427018 570022 427254
rect 569786 426698 570022 426934
rect 569786 391018 570022 391254
rect 569786 390698 570022 390934
rect 569786 355018 570022 355254
rect 569786 354698 570022 354934
rect 569786 319018 570022 319254
rect 569786 318698 570022 318934
rect 569786 283018 570022 283254
rect 569786 282698 570022 282934
rect 569786 247018 570022 247254
rect 569786 246698 570022 246934
rect 569786 211018 570022 211254
rect 569786 210698 570022 210934
rect 569786 175018 570022 175254
rect 569786 174698 570022 174934
rect 569786 139018 570022 139254
rect 569786 138698 570022 138934
rect 569786 103018 570022 103254
rect 569786 102698 570022 102934
rect 569786 67018 570022 67254
rect 569786 66698 570022 66934
rect 569786 31018 570022 31254
rect 569786 30698 570022 30934
rect 551786 -6102 552022 -5866
rect 551786 -6422 552022 -6186
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 576986 686218 577222 686454
rect 576986 685898 577222 686134
rect 576986 650218 577222 650454
rect 576986 649898 577222 650134
rect 576986 614218 577222 614454
rect 576986 613898 577222 614134
rect 576986 578218 577222 578454
rect 576986 577898 577222 578134
rect 576986 542218 577222 542454
rect 576986 541898 577222 542134
rect 576986 506218 577222 506454
rect 576986 505898 577222 506134
rect 576986 470218 577222 470454
rect 576986 469898 577222 470134
rect 576986 434218 577222 434454
rect 576986 433898 577222 434134
rect 576986 398218 577222 398454
rect 576986 397898 577222 398134
rect 576986 362218 577222 362454
rect 576986 361898 577222 362134
rect 576986 326218 577222 326454
rect 576986 325898 577222 326134
rect 576986 290218 577222 290454
rect 576986 289898 577222 290134
rect 576986 254218 577222 254454
rect 576986 253898 577222 254134
rect 576986 218218 577222 218454
rect 576986 217898 577222 218134
rect 576986 182218 577222 182454
rect 576986 181898 577222 182134
rect 576986 146218 577222 146454
rect 576986 145898 577222 146134
rect 576986 110218 577222 110454
rect 576986 109898 577222 110134
rect 576986 74218 577222 74454
rect 576986 73898 577222 74134
rect 576986 38218 577222 38454
rect 576986 37898 577222 38134
rect 576986 2218 577222 2454
rect 576986 1898 577222 2134
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 587342 706442 587578 706678
rect 587342 706122 587578 706358
rect 586422 705522 586658 705758
rect 586422 705202 586658 705438
rect 580586 689818 580822 690054
rect 580586 689498 580822 689734
rect 580586 653818 580822 654054
rect 580586 653498 580822 653734
rect 580586 617818 580822 618054
rect 580586 617498 580822 617734
rect 580586 581818 580822 582054
rect 580586 581498 580822 581734
rect 580586 545818 580822 546054
rect 580586 545498 580822 545734
rect 580586 509818 580822 510054
rect 580586 509498 580822 509734
rect 580586 473818 580822 474054
rect 580586 473498 580822 473734
rect 580586 437818 580822 438054
rect 580586 437498 580822 437734
rect 580586 401818 580822 402054
rect 580586 401498 580822 401734
rect 580586 365818 580822 366054
rect 580586 365498 580822 365734
rect 580586 329818 580822 330054
rect 580586 329498 580822 329734
rect 580586 293818 580822 294054
rect 580586 293498 580822 293734
rect 580586 257818 580822 258054
rect 580586 257498 580822 257734
rect 580586 221818 580822 222054
rect 580586 221498 580822 221734
rect 580586 185818 580822 186054
rect 580586 185498 580822 185734
rect 580586 149818 580822 150054
rect 580586 149498 580822 149734
rect 580586 113818 580822 114054
rect 580586 113498 580822 113734
rect 580586 77818 580822 78054
rect 580586 77498 580822 77734
rect 580586 41818 580822 42054
rect 580586 41498 580822 41734
rect 580586 5818 580822 6054
rect 580586 5498 580822 5734
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 686218 585738 686454
rect 585502 685898 585738 686134
rect 585502 650218 585738 650454
rect 585502 649898 585738 650134
rect 585502 614218 585738 614454
rect 585502 613898 585738 614134
rect 585502 578218 585738 578454
rect 585502 577898 585738 578134
rect 585502 542218 585738 542454
rect 585502 541898 585738 542134
rect 585502 506218 585738 506454
rect 585502 505898 585738 506134
rect 585502 470218 585738 470454
rect 585502 469898 585738 470134
rect 585502 434218 585738 434454
rect 585502 433898 585738 434134
rect 585502 398218 585738 398454
rect 585502 397898 585738 398134
rect 585502 362218 585738 362454
rect 585502 361898 585738 362134
rect 585502 326218 585738 326454
rect 585502 325898 585738 326134
rect 585502 290218 585738 290454
rect 585502 289898 585738 290134
rect 585502 254218 585738 254454
rect 585502 253898 585738 254134
rect 585502 218218 585738 218454
rect 585502 217898 585738 218134
rect 585502 182218 585738 182454
rect 585502 181898 585738 182134
rect 585502 146218 585738 146454
rect 585502 145898 585738 146134
rect 585502 110218 585738 110454
rect 585502 109898 585738 110134
rect 585502 74218 585738 74454
rect 585502 73898 585738 74134
rect 585502 38218 585738 38454
rect 585502 37898 585738 38134
rect 585502 2218 585738 2454
rect 585502 1898 585738 2134
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586422 668218 586658 668454
rect 586422 667898 586658 668134
rect 586422 632218 586658 632454
rect 586422 631898 586658 632134
rect 586422 596218 586658 596454
rect 586422 595898 586658 596134
rect 586422 560218 586658 560454
rect 586422 559898 586658 560134
rect 586422 524218 586658 524454
rect 586422 523898 586658 524134
rect 586422 488218 586658 488454
rect 586422 487898 586658 488134
rect 586422 452218 586658 452454
rect 586422 451898 586658 452134
rect 586422 416218 586658 416454
rect 586422 415898 586658 416134
rect 586422 380218 586658 380454
rect 586422 379898 586658 380134
rect 586422 344218 586658 344454
rect 586422 343898 586658 344134
rect 586422 308218 586658 308454
rect 586422 307898 586658 308134
rect 586422 272218 586658 272454
rect 586422 271898 586658 272134
rect 586422 236218 586658 236454
rect 586422 235898 586658 236134
rect 586422 200218 586658 200454
rect 586422 199898 586658 200134
rect 586422 164218 586658 164454
rect 586422 163898 586658 164134
rect 586422 128218 586658 128454
rect 586422 127898 586658 128134
rect 586422 92218 586658 92454
rect 586422 91898 586658 92134
rect 586422 56218 586658 56454
rect 586422 55898 586658 56134
rect 586422 20218 586658 20454
rect 586422 19898 586658 20134
rect 586422 -1502 586658 -1266
rect 586422 -1822 586658 -1586
rect 587342 689818 587578 690054
rect 587342 689498 587578 689734
rect 587342 653818 587578 654054
rect 587342 653498 587578 653734
rect 587342 617818 587578 618054
rect 587342 617498 587578 617734
rect 587342 581818 587578 582054
rect 587342 581498 587578 581734
rect 587342 545818 587578 546054
rect 587342 545498 587578 545734
rect 587342 509818 587578 510054
rect 587342 509498 587578 509734
rect 587342 473818 587578 474054
rect 587342 473498 587578 473734
rect 587342 437818 587578 438054
rect 587342 437498 587578 437734
rect 587342 401818 587578 402054
rect 587342 401498 587578 401734
rect 587342 365818 587578 366054
rect 587342 365498 587578 365734
rect 587342 329818 587578 330054
rect 587342 329498 587578 329734
rect 587342 293818 587578 294054
rect 587342 293498 587578 293734
rect 587342 257818 587578 258054
rect 587342 257498 587578 257734
rect 587342 221818 587578 222054
rect 587342 221498 587578 221734
rect 587342 185818 587578 186054
rect 587342 185498 587578 185734
rect 587342 149818 587578 150054
rect 587342 149498 587578 149734
rect 587342 113818 587578 114054
rect 587342 113498 587578 113734
rect 587342 77818 587578 78054
rect 587342 77498 587578 77734
rect 587342 41818 587578 42054
rect 587342 41498 587578 41734
rect 587342 5818 587578 6054
rect 587342 5498 587578 5734
rect 580586 -2422 580822 -2186
rect 580586 -2742 580822 -2506
rect 587342 -2422 587578 -2186
rect 587342 -2742 587578 -2506
rect 588262 671818 588498 672054
rect 588262 671498 588498 671734
rect 588262 635818 588498 636054
rect 588262 635498 588498 635734
rect 588262 599818 588498 600054
rect 588262 599498 588498 599734
rect 588262 563818 588498 564054
rect 588262 563498 588498 563734
rect 588262 527818 588498 528054
rect 588262 527498 588498 527734
rect 588262 491818 588498 492054
rect 588262 491498 588498 491734
rect 588262 455818 588498 456054
rect 588262 455498 588498 455734
rect 588262 419818 588498 420054
rect 588262 419498 588498 419734
rect 588262 383818 588498 384054
rect 588262 383498 588498 383734
rect 588262 347818 588498 348054
rect 588262 347498 588498 347734
rect 588262 311818 588498 312054
rect 588262 311498 588498 311734
rect 588262 275818 588498 276054
rect 588262 275498 588498 275734
rect 588262 239818 588498 240054
rect 588262 239498 588498 239734
rect 588262 203818 588498 204054
rect 588262 203498 588498 203734
rect 588262 167818 588498 168054
rect 588262 167498 588498 167734
rect 588262 131818 588498 132054
rect 588262 131498 588498 131734
rect 588262 95818 588498 96054
rect 588262 95498 588498 95734
rect 588262 59818 588498 60054
rect 588262 59498 588498 59734
rect 588262 23818 588498 24054
rect 588262 23498 588498 23734
rect 588262 -3342 588498 -3106
rect 588262 -3662 588498 -3426
rect 589182 693418 589418 693654
rect 589182 693098 589418 693334
rect 589182 657418 589418 657654
rect 589182 657098 589418 657334
rect 589182 621418 589418 621654
rect 589182 621098 589418 621334
rect 589182 585418 589418 585654
rect 589182 585098 589418 585334
rect 589182 549418 589418 549654
rect 589182 549098 589418 549334
rect 589182 513418 589418 513654
rect 589182 513098 589418 513334
rect 589182 477418 589418 477654
rect 589182 477098 589418 477334
rect 589182 441418 589418 441654
rect 589182 441098 589418 441334
rect 589182 405418 589418 405654
rect 589182 405098 589418 405334
rect 589182 369418 589418 369654
rect 589182 369098 589418 369334
rect 589182 333418 589418 333654
rect 589182 333098 589418 333334
rect 589182 297418 589418 297654
rect 589182 297098 589418 297334
rect 589182 261418 589418 261654
rect 589182 261098 589418 261334
rect 589182 225418 589418 225654
rect 589182 225098 589418 225334
rect 589182 189418 589418 189654
rect 589182 189098 589418 189334
rect 589182 153418 589418 153654
rect 589182 153098 589418 153334
rect 589182 117418 589418 117654
rect 589182 117098 589418 117334
rect 589182 81418 589418 81654
rect 589182 81098 589418 81334
rect 589182 45418 589418 45654
rect 589182 45098 589418 45334
rect 589182 9418 589418 9654
rect 589182 9098 589418 9334
rect 589182 -4262 589418 -4026
rect 589182 -4582 589418 -4346
rect 590102 675418 590338 675654
rect 590102 675098 590338 675334
rect 590102 639418 590338 639654
rect 590102 639098 590338 639334
rect 590102 603418 590338 603654
rect 590102 603098 590338 603334
rect 590102 567418 590338 567654
rect 590102 567098 590338 567334
rect 590102 531418 590338 531654
rect 590102 531098 590338 531334
rect 590102 495418 590338 495654
rect 590102 495098 590338 495334
rect 590102 459418 590338 459654
rect 590102 459098 590338 459334
rect 590102 423418 590338 423654
rect 590102 423098 590338 423334
rect 590102 387418 590338 387654
rect 590102 387098 590338 387334
rect 590102 351418 590338 351654
rect 590102 351098 590338 351334
rect 590102 315418 590338 315654
rect 590102 315098 590338 315334
rect 590102 279418 590338 279654
rect 590102 279098 590338 279334
rect 590102 243418 590338 243654
rect 590102 243098 590338 243334
rect 590102 207418 590338 207654
rect 590102 207098 590338 207334
rect 590102 171418 590338 171654
rect 590102 171098 590338 171334
rect 590102 135418 590338 135654
rect 590102 135098 590338 135334
rect 590102 99418 590338 99654
rect 590102 99098 590338 99334
rect 590102 63418 590338 63654
rect 590102 63098 590338 63334
rect 590102 27418 590338 27654
rect 590102 27098 590338 27334
rect 590102 -5182 590338 -4946
rect 590102 -5502 590338 -5266
rect 591022 697018 591258 697254
rect 591022 696698 591258 696934
rect 591022 661018 591258 661254
rect 591022 660698 591258 660934
rect 591022 625018 591258 625254
rect 591022 624698 591258 624934
rect 591022 589018 591258 589254
rect 591022 588698 591258 588934
rect 591022 553018 591258 553254
rect 591022 552698 591258 552934
rect 591022 517018 591258 517254
rect 591022 516698 591258 516934
rect 591022 481018 591258 481254
rect 591022 480698 591258 480934
rect 591022 445018 591258 445254
rect 591022 444698 591258 444934
rect 591022 409018 591258 409254
rect 591022 408698 591258 408934
rect 591022 373018 591258 373254
rect 591022 372698 591258 372934
rect 591022 337018 591258 337254
rect 591022 336698 591258 336934
rect 591022 301018 591258 301254
rect 591022 300698 591258 300934
rect 591022 265018 591258 265254
rect 591022 264698 591258 264934
rect 591022 229018 591258 229254
rect 591022 228698 591258 228934
rect 591022 193018 591258 193254
rect 591022 192698 591258 192934
rect 591022 157018 591258 157254
rect 591022 156698 591258 156934
rect 591022 121018 591258 121254
rect 591022 120698 591258 120934
rect 591022 85018 591258 85254
rect 591022 84698 591258 84934
rect 591022 49018 591258 49254
rect 591022 48698 591258 48934
rect 591022 13018 591258 13254
rect 591022 12698 591258 12934
rect 591022 -6102 591258 -5866
rect 591022 -6422 591258 -6186
rect 591942 679018 592178 679254
rect 591942 678698 592178 678934
rect 591942 643018 592178 643254
rect 591942 642698 592178 642934
rect 591942 607018 592178 607254
rect 591942 606698 592178 606934
rect 591942 571018 592178 571254
rect 591942 570698 592178 570934
rect 591942 535018 592178 535254
rect 591942 534698 592178 534934
rect 591942 499018 592178 499254
rect 591942 498698 592178 498934
rect 591942 463018 592178 463254
rect 591942 462698 592178 462934
rect 591942 427018 592178 427254
rect 591942 426698 592178 426934
rect 591942 391018 592178 391254
rect 591942 390698 592178 390934
rect 591942 355018 592178 355254
rect 591942 354698 592178 354934
rect 591942 319018 592178 319254
rect 591942 318698 592178 318934
rect 591942 283018 592178 283254
rect 591942 282698 592178 282934
rect 591942 247018 592178 247254
rect 591942 246698 592178 246934
rect 591942 211018 592178 211254
rect 591942 210698 592178 210934
rect 591942 175018 592178 175254
rect 591942 174698 592178 174934
rect 591942 139018 592178 139254
rect 591942 138698 592178 138934
rect 591942 103018 592178 103254
rect 591942 102698 592178 102934
rect 591942 67018 592178 67254
rect 591942 66698 592178 66934
rect 591942 31018 592178 31254
rect 591942 30698 592178 30934
rect 569786 -7022 570022 -6786
rect 569786 -7342 570022 -7106
rect 591942 -7022 592178 -6786
rect 591942 -7342 592178 -7106
<< metal5 >>
rect -8436 711300 -7836 711302
rect 29604 711300 30204 711302
rect 65604 711300 66204 711302
rect 101604 711300 102204 711302
rect 137604 711300 138204 711302
rect 173604 711300 174204 711302
rect 209604 711300 210204 711302
rect 245604 711300 246204 711302
rect 281604 711300 282204 711302
rect 317604 711300 318204 711302
rect 353604 711300 354204 711302
rect 389604 711300 390204 711302
rect 425604 711300 426204 711302
rect 461604 711300 462204 711302
rect 497604 711300 498204 711302
rect 533604 711300 534204 711302
rect 569604 711300 570204 711302
rect 591760 711300 592360 711302
rect -8436 711278 592360 711300
rect -8436 711042 -8254 711278
rect -8018 711042 29786 711278
rect 30022 711042 65786 711278
rect 66022 711042 101786 711278
rect 102022 711042 137786 711278
rect 138022 711042 173786 711278
rect 174022 711042 209786 711278
rect 210022 711042 245786 711278
rect 246022 711042 281786 711278
rect 282022 711042 317786 711278
rect 318022 711042 353786 711278
rect 354022 711042 389786 711278
rect 390022 711042 425786 711278
rect 426022 711042 461786 711278
rect 462022 711042 497786 711278
rect 498022 711042 533786 711278
rect 534022 711042 569786 711278
rect 570022 711042 591942 711278
rect 592178 711042 592360 711278
rect -8436 710958 592360 711042
rect -8436 710722 -8254 710958
rect -8018 710722 29786 710958
rect 30022 710722 65786 710958
rect 66022 710722 101786 710958
rect 102022 710722 137786 710958
rect 138022 710722 173786 710958
rect 174022 710722 209786 710958
rect 210022 710722 245786 710958
rect 246022 710722 281786 710958
rect 282022 710722 317786 710958
rect 318022 710722 353786 710958
rect 354022 710722 389786 710958
rect 390022 710722 425786 710958
rect 426022 710722 461786 710958
rect 462022 710722 497786 710958
rect 498022 710722 533786 710958
rect 534022 710722 569786 710958
rect 570022 710722 591942 710958
rect 592178 710722 592360 710958
rect -8436 710700 592360 710722
rect -8436 710698 -7836 710700
rect 29604 710698 30204 710700
rect 65604 710698 66204 710700
rect 101604 710698 102204 710700
rect 137604 710698 138204 710700
rect 173604 710698 174204 710700
rect 209604 710698 210204 710700
rect 245604 710698 246204 710700
rect 281604 710698 282204 710700
rect 317604 710698 318204 710700
rect 353604 710698 354204 710700
rect 389604 710698 390204 710700
rect 425604 710698 426204 710700
rect 461604 710698 462204 710700
rect 497604 710698 498204 710700
rect 533604 710698 534204 710700
rect 569604 710698 570204 710700
rect 591760 710698 592360 710700
rect -7516 710380 -6916 710382
rect 11604 710380 12204 710382
rect 47604 710380 48204 710382
rect 83604 710380 84204 710382
rect 119604 710380 120204 710382
rect 155604 710380 156204 710382
rect 191604 710380 192204 710382
rect 227604 710380 228204 710382
rect 263604 710380 264204 710382
rect 299604 710380 300204 710382
rect 335604 710380 336204 710382
rect 371604 710380 372204 710382
rect 407604 710380 408204 710382
rect 443604 710380 444204 710382
rect 479604 710380 480204 710382
rect 515604 710380 516204 710382
rect 551604 710380 552204 710382
rect 590840 710380 591440 710382
rect -7516 710358 591440 710380
rect -7516 710122 -7334 710358
rect -7098 710122 11786 710358
rect 12022 710122 47786 710358
rect 48022 710122 83786 710358
rect 84022 710122 119786 710358
rect 120022 710122 155786 710358
rect 156022 710122 191786 710358
rect 192022 710122 227786 710358
rect 228022 710122 263786 710358
rect 264022 710122 299786 710358
rect 300022 710122 335786 710358
rect 336022 710122 371786 710358
rect 372022 710122 407786 710358
rect 408022 710122 443786 710358
rect 444022 710122 479786 710358
rect 480022 710122 515786 710358
rect 516022 710122 551786 710358
rect 552022 710122 591022 710358
rect 591258 710122 591440 710358
rect -7516 710038 591440 710122
rect -7516 709802 -7334 710038
rect -7098 709802 11786 710038
rect 12022 709802 47786 710038
rect 48022 709802 83786 710038
rect 84022 709802 119786 710038
rect 120022 709802 155786 710038
rect 156022 709802 191786 710038
rect 192022 709802 227786 710038
rect 228022 709802 263786 710038
rect 264022 709802 299786 710038
rect 300022 709802 335786 710038
rect 336022 709802 371786 710038
rect 372022 709802 407786 710038
rect 408022 709802 443786 710038
rect 444022 709802 479786 710038
rect 480022 709802 515786 710038
rect 516022 709802 551786 710038
rect 552022 709802 591022 710038
rect 591258 709802 591440 710038
rect -7516 709780 591440 709802
rect -7516 709778 -6916 709780
rect 11604 709778 12204 709780
rect 47604 709778 48204 709780
rect 83604 709778 84204 709780
rect 119604 709778 120204 709780
rect 155604 709778 156204 709780
rect 191604 709778 192204 709780
rect 227604 709778 228204 709780
rect 263604 709778 264204 709780
rect 299604 709778 300204 709780
rect 335604 709778 336204 709780
rect 371604 709778 372204 709780
rect 407604 709778 408204 709780
rect 443604 709778 444204 709780
rect 479604 709778 480204 709780
rect 515604 709778 516204 709780
rect 551604 709778 552204 709780
rect 590840 709778 591440 709780
rect -6596 709460 -5996 709462
rect 26004 709460 26604 709462
rect 62004 709460 62604 709462
rect 98004 709460 98604 709462
rect 134004 709460 134604 709462
rect 170004 709460 170604 709462
rect 206004 709460 206604 709462
rect 242004 709460 242604 709462
rect 278004 709460 278604 709462
rect 314004 709460 314604 709462
rect 350004 709460 350604 709462
rect 386004 709460 386604 709462
rect 422004 709460 422604 709462
rect 458004 709460 458604 709462
rect 494004 709460 494604 709462
rect 530004 709460 530604 709462
rect 566004 709460 566604 709462
rect 589920 709460 590520 709462
rect -6596 709438 590520 709460
rect -6596 709202 -6414 709438
rect -6178 709202 26186 709438
rect 26422 709202 62186 709438
rect 62422 709202 98186 709438
rect 98422 709202 134186 709438
rect 134422 709202 170186 709438
rect 170422 709202 206186 709438
rect 206422 709202 242186 709438
rect 242422 709202 278186 709438
rect 278422 709202 314186 709438
rect 314422 709202 350186 709438
rect 350422 709202 386186 709438
rect 386422 709202 422186 709438
rect 422422 709202 458186 709438
rect 458422 709202 494186 709438
rect 494422 709202 530186 709438
rect 530422 709202 566186 709438
rect 566422 709202 590102 709438
rect 590338 709202 590520 709438
rect -6596 709118 590520 709202
rect -6596 708882 -6414 709118
rect -6178 708882 26186 709118
rect 26422 708882 62186 709118
rect 62422 708882 98186 709118
rect 98422 708882 134186 709118
rect 134422 708882 170186 709118
rect 170422 708882 206186 709118
rect 206422 708882 242186 709118
rect 242422 708882 278186 709118
rect 278422 708882 314186 709118
rect 314422 708882 350186 709118
rect 350422 708882 386186 709118
rect 386422 708882 422186 709118
rect 422422 708882 458186 709118
rect 458422 708882 494186 709118
rect 494422 708882 530186 709118
rect 530422 708882 566186 709118
rect 566422 708882 590102 709118
rect 590338 708882 590520 709118
rect -6596 708860 590520 708882
rect -6596 708858 -5996 708860
rect 26004 708858 26604 708860
rect 62004 708858 62604 708860
rect 98004 708858 98604 708860
rect 134004 708858 134604 708860
rect 170004 708858 170604 708860
rect 206004 708858 206604 708860
rect 242004 708858 242604 708860
rect 278004 708858 278604 708860
rect 314004 708858 314604 708860
rect 350004 708858 350604 708860
rect 386004 708858 386604 708860
rect 422004 708858 422604 708860
rect 458004 708858 458604 708860
rect 494004 708858 494604 708860
rect 530004 708858 530604 708860
rect 566004 708858 566604 708860
rect 589920 708858 590520 708860
rect -5676 708540 -5076 708542
rect 8004 708540 8604 708542
rect 44004 708540 44604 708542
rect 80004 708540 80604 708542
rect 116004 708540 116604 708542
rect 152004 708540 152604 708542
rect 188004 708540 188604 708542
rect 224004 708540 224604 708542
rect 260004 708540 260604 708542
rect 296004 708540 296604 708542
rect 332004 708540 332604 708542
rect 368004 708540 368604 708542
rect 404004 708540 404604 708542
rect 440004 708540 440604 708542
rect 476004 708540 476604 708542
rect 512004 708540 512604 708542
rect 548004 708540 548604 708542
rect 589000 708540 589600 708542
rect -5676 708518 589600 708540
rect -5676 708282 -5494 708518
rect -5258 708282 8186 708518
rect 8422 708282 44186 708518
rect 44422 708282 80186 708518
rect 80422 708282 116186 708518
rect 116422 708282 152186 708518
rect 152422 708282 188186 708518
rect 188422 708282 224186 708518
rect 224422 708282 260186 708518
rect 260422 708282 296186 708518
rect 296422 708282 332186 708518
rect 332422 708282 368186 708518
rect 368422 708282 404186 708518
rect 404422 708282 440186 708518
rect 440422 708282 476186 708518
rect 476422 708282 512186 708518
rect 512422 708282 548186 708518
rect 548422 708282 589182 708518
rect 589418 708282 589600 708518
rect -5676 708198 589600 708282
rect -5676 707962 -5494 708198
rect -5258 707962 8186 708198
rect 8422 707962 44186 708198
rect 44422 707962 80186 708198
rect 80422 707962 116186 708198
rect 116422 707962 152186 708198
rect 152422 707962 188186 708198
rect 188422 707962 224186 708198
rect 224422 707962 260186 708198
rect 260422 707962 296186 708198
rect 296422 707962 332186 708198
rect 332422 707962 368186 708198
rect 368422 707962 404186 708198
rect 404422 707962 440186 708198
rect 440422 707962 476186 708198
rect 476422 707962 512186 708198
rect 512422 707962 548186 708198
rect 548422 707962 589182 708198
rect 589418 707962 589600 708198
rect -5676 707940 589600 707962
rect -5676 707938 -5076 707940
rect 8004 707938 8604 707940
rect 44004 707938 44604 707940
rect 80004 707938 80604 707940
rect 116004 707938 116604 707940
rect 152004 707938 152604 707940
rect 188004 707938 188604 707940
rect 224004 707938 224604 707940
rect 260004 707938 260604 707940
rect 296004 707938 296604 707940
rect 332004 707938 332604 707940
rect 368004 707938 368604 707940
rect 404004 707938 404604 707940
rect 440004 707938 440604 707940
rect 476004 707938 476604 707940
rect 512004 707938 512604 707940
rect 548004 707938 548604 707940
rect 589000 707938 589600 707940
rect -4756 707620 -4156 707622
rect 22404 707620 23004 707622
rect 58404 707620 59004 707622
rect 94404 707620 95004 707622
rect 130404 707620 131004 707622
rect 166404 707620 167004 707622
rect 202404 707620 203004 707622
rect 238404 707620 239004 707622
rect 274404 707620 275004 707622
rect 310404 707620 311004 707622
rect 346404 707620 347004 707622
rect 382404 707620 383004 707622
rect 418404 707620 419004 707622
rect 454404 707620 455004 707622
rect 490404 707620 491004 707622
rect 526404 707620 527004 707622
rect 562404 707620 563004 707622
rect 588080 707620 588680 707622
rect -4756 707598 588680 707620
rect -4756 707362 -4574 707598
rect -4338 707362 22586 707598
rect 22822 707362 58586 707598
rect 58822 707362 94586 707598
rect 94822 707362 130586 707598
rect 130822 707362 166586 707598
rect 166822 707362 202586 707598
rect 202822 707362 238586 707598
rect 238822 707362 274586 707598
rect 274822 707362 310586 707598
rect 310822 707362 346586 707598
rect 346822 707362 382586 707598
rect 382822 707362 418586 707598
rect 418822 707362 454586 707598
rect 454822 707362 490586 707598
rect 490822 707362 526586 707598
rect 526822 707362 562586 707598
rect 562822 707362 588262 707598
rect 588498 707362 588680 707598
rect -4756 707278 588680 707362
rect -4756 707042 -4574 707278
rect -4338 707042 22586 707278
rect 22822 707042 58586 707278
rect 58822 707042 94586 707278
rect 94822 707042 130586 707278
rect 130822 707042 166586 707278
rect 166822 707042 202586 707278
rect 202822 707042 238586 707278
rect 238822 707042 274586 707278
rect 274822 707042 310586 707278
rect 310822 707042 346586 707278
rect 346822 707042 382586 707278
rect 382822 707042 418586 707278
rect 418822 707042 454586 707278
rect 454822 707042 490586 707278
rect 490822 707042 526586 707278
rect 526822 707042 562586 707278
rect 562822 707042 588262 707278
rect 588498 707042 588680 707278
rect -4756 707020 588680 707042
rect -4756 707018 -4156 707020
rect 22404 707018 23004 707020
rect 58404 707018 59004 707020
rect 94404 707018 95004 707020
rect 130404 707018 131004 707020
rect 166404 707018 167004 707020
rect 202404 707018 203004 707020
rect 238404 707018 239004 707020
rect 274404 707018 275004 707020
rect 310404 707018 311004 707020
rect 346404 707018 347004 707020
rect 382404 707018 383004 707020
rect 418404 707018 419004 707020
rect 454404 707018 455004 707020
rect 490404 707018 491004 707020
rect 526404 707018 527004 707020
rect 562404 707018 563004 707020
rect 588080 707018 588680 707020
rect -3836 706700 -3236 706702
rect 4404 706700 5004 706702
rect 40404 706700 41004 706702
rect 76404 706700 77004 706702
rect 112404 706700 113004 706702
rect 148404 706700 149004 706702
rect 184404 706700 185004 706702
rect 220404 706700 221004 706702
rect 256404 706700 257004 706702
rect 292404 706700 293004 706702
rect 328404 706700 329004 706702
rect 364404 706700 365004 706702
rect 400404 706700 401004 706702
rect 436404 706700 437004 706702
rect 472404 706700 473004 706702
rect 508404 706700 509004 706702
rect 544404 706700 545004 706702
rect 580404 706700 581004 706702
rect 587160 706700 587760 706702
rect -3836 706678 587760 706700
rect -3836 706442 -3654 706678
rect -3418 706442 4586 706678
rect 4822 706442 40586 706678
rect 40822 706442 76586 706678
rect 76822 706442 112586 706678
rect 112822 706442 148586 706678
rect 148822 706442 184586 706678
rect 184822 706442 220586 706678
rect 220822 706442 256586 706678
rect 256822 706442 292586 706678
rect 292822 706442 328586 706678
rect 328822 706442 364586 706678
rect 364822 706442 400586 706678
rect 400822 706442 436586 706678
rect 436822 706442 472586 706678
rect 472822 706442 508586 706678
rect 508822 706442 544586 706678
rect 544822 706442 580586 706678
rect 580822 706442 587342 706678
rect 587578 706442 587760 706678
rect -3836 706358 587760 706442
rect -3836 706122 -3654 706358
rect -3418 706122 4586 706358
rect 4822 706122 40586 706358
rect 40822 706122 76586 706358
rect 76822 706122 112586 706358
rect 112822 706122 148586 706358
rect 148822 706122 184586 706358
rect 184822 706122 220586 706358
rect 220822 706122 256586 706358
rect 256822 706122 292586 706358
rect 292822 706122 328586 706358
rect 328822 706122 364586 706358
rect 364822 706122 400586 706358
rect 400822 706122 436586 706358
rect 436822 706122 472586 706358
rect 472822 706122 508586 706358
rect 508822 706122 544586 706358
rect 544822 706122 580586 706358
rect 580822 706122 587342 706358
rect 587578 706122 587760 706358
rect -3836 706100 587760 706122
rect -3836 706098 -3236 706100
rect 4404 706098 5004 706100
rect 40404 706098 41004 706100
rect 76404 706098 77004 706100
rect 112404 706098 113004 706100
rect 148404 706098 149004 706100
rect 184404 706098 185004 706100
rect 220404 706098 221004 706100
rect 256404 706098 257004 706100
rect 292404 706098 293004 706100
rect 328404 706098 329004 706100
rect 364404 706098 365004 706100
rect 400404 706098 401004 706100
rect 436404 706098 437004 706100
rect 472404 706098 473004 706100
rect 508404 706098 509004 706100
rect 544404 706098 545004 706100
rect 580404 706098 581004 706100
rect 587160 706098 587760 706100
rect -2916 705780 -2316 705782
rect 18804 705780 19404 705782
rect 54804 705780 55404 705782
rect 90804 705780 91404 705782
rect 126804 705780 127404 705782
rect 162804 705780 163404 705782
rect 198804 705780 199404 705782
rect 234804 705780 235404 705782
rect 270804 705780 271404 705782
rect 306804 705780 307404 705782
rect 342804 705780 343404 705782
rect 378804 705780 379404 705782
rect 414804 705780 415404 705782
rect 450804 705780 451404 705782
rect 486804 705780 487404 705782
rect 522804 705780 523404 705782
rect 558804 705780 559404 705782
rect 586240 705780 586840 705782
rect -2916 705758 586840 705780
rect -2916 705522 -2734 705758
rect -2498 705522 18986 705758
rect 19222 705522 54986 705758
rect 55222 705522 90986 705758
rect 91222 705522 126986 705758
rect 127222 705522 162986 705758
rect 163222 705522 198986 705758
rect 199222 705522 234986 705758
rect 235222 705522 270986 705758
rect 271222 705522 306986 705758
rect 307222 705522 342986 705758
rect 343222 705522 378986 705758
rect 379222 705522 414986 705758
rect 415222 705522 450986 705758
rect 451222 705522 486986 705758
rect 487222 705522 522986 705758
rect 523222 705522 558986 705758
rect 559222 705522 586422 705758
rect 586658 705522 586840 705758
rect -2916 705438 586840 705522
rect -2916 705202 -2734 705438
rect -2498 705202 18986 705438
rect 19222 705202 54986 705438
rect 55222 705202 90986 705438
rect 91222 705202 126986 705438
rect 127222 705202 162986 705438
rect 163222 705202 198986 705438
rect 199222 705202 234986 705438
rect 235222 705202 270986 705438
rect 271222 705202 306986 705438
rect 307222 705202 342986 705438
rect 343222 705202 378986 705438
rect 379222 705202 414986 705438
rect 415222 705202 450986 705438
rect 451222 705202 486986 705438
rect 487222 705202 522986 705438
rect 523222 705202 558986 705438
rect 559222 705202 586422 705438
rect 586658 705202 586840 705438
rect -2916 705180 586840 705202
rect -2916 705178 -2316 705180
rect 18804 705178 19404 705180
rect 54804 705178 55404 705180
rect 90804 705178 91404 705180
rect 126804 705178 127404 705180
rect 162804 705178 163404 705180
rect 198804 705178 199404 705180
rect 234804 705178 235404 705180
rect 270804 705178 271404 705180
rect 306804 705178 307404 705180
rect 342804 705178 343404 705180
rect 378804 705178 379404 705180
rect 414804 705178 415404 705180
rect 450804 705178 451404 705180
rect 486804 705178 487404 705180
rect 522804 705178 523404 705180
rect 558804 705178 559404 705180
rect 586240 705178 586840 705180
rect -1996 704860 -1396 704862
rect 804 704860 1404 704862
rect 36804 704860 37404 704862
rect 72804 704860 73404 704862
rect 108804 704860 109404 704862
rect 144804 704860 145404 704862
rect 180804 704860 181404 704862
rect 216804 704860 217404 704862
rect 252804 704860 253404 704862
rect 288804 704860 289404 704862
rect 324804 704860 325404 704862
rect 360804 704860 361404 704862
rect 396804 704860 397404 704862
rect 432804 704860 433404 704862
rect 468804 704860 469404 704862
rect 504804 704860 505404 704862
rect 540804 704860 541404 704862
rect 576804 704860 577404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 804 704258 1404 704260
rect 36804 704258 37404 704260
rect 72804 704258 73404 704260
rect 108804 704258 109404 704260
rect 144804 704258 145404 704260
rect 180804 704258 181404 704260
rect 216804 704258 217404 704260
rect 252804 704258 253404 704260
rect 288804 704258 289404 704260
rect 324804 704258 325404 704260
rect 360804 704258 361404 704260
rect 396804 704258 397404 704260
rect 432804 704258 433404 704260
rect 468804 704258 469404 704260
rect 504804 704258 505404 704260
rect 540804 704258 541404 704260
rect 576804 704258 577404 704260
rect 585320 704258 585920 704260
rect -7516 697276 -6916 697278
rect 11604 697276 12204 697278
rect 47604 697276 48204 697278
rect 83604 697276 84204 697278
rect 119604 697276 120204 697278
rect 155604 697276 156204 697278
rect 191604 697276 192204 697278
rect 227604 697276 228204 697278
rect 263604 697276 264204 697278
rect 299604 697276 300204 697278
rect 335604 697276 336204 697278
rect 371604 697276 372204 697278
rect 407604 697276 408204 697278
rect 443604 697276 444204 697278
rect 479604 697276 480204 697278
rect 515604 697276 516204 697278
rect 551604 697276 552204 697278
rect 590840 697276 591440 697278
rect -8436 697254 592360 697276
rect -8436 697018 -7334 697254
rect -7098 697018 11786 697254
rect 12022 697018 47786 697254
rect 48022 697018 83786 697254
rect 84022 697018 119786 697254
rect 120022 697018 155786 697254
rect 156022 697018 191786 697254
rect 192022 697018 227786 697254
rect 228022 697018 263786 697254
rect 264022 697018 299786 697254
rect 300022 697018 335786 697254
rect 336022 697018 371786 697254
rect 372022 697018 407786 697254
rect 408022 697018 443786 697254
rect 444022 697018 479786 697254
rect 480022 697018 515786 697254
rect 516022 697018 551786 697254
rect 552022 697018 591022 697254
rect 591258 697018 592360 697254
rect -8436 696934 592360 697018
rect -8436 696698 -7334 696934
rect -7098 696698 11786 696934
rect 12022 696698 47786 696934
rect 48022 696698 83786 696934
rect 84022 696698 119786 696934
rect 120022 696698 155786 696934
rect 156022 696698 191786 696934
rect 192022 696698 227786 696934
rect 228022 696698 263786 696934
rect 264022 696698 299786 696934
rect 300022 696698 335786 696934
rect 336022 696698 371786 696934
rect 372022 696698 407786 696934
rect 408022 696698 443786 696934
rect 444022 696698 479786 696934
rect 480022 696698 515786 696934
rect 516022 696698 551786 696934
rect 552022 696698 591022 696934
rect 591258 696698 592360 696934
rect -8436 696676 592360 696698
rect -7516 696674 -6916 696676
rect 11604 696674 12204 696676
rect 47604 696674 48204 696676
rect 83604 696674 84204 696676
rect 119604 696674 120204 696676
rect 155604 696674 156204 696676
rect 191604 696674 192204 696676
rect 227604 696674 228204 696676
rect 263604 696674 264204 696676
rect 299604 696674 300204 696676
rect 335604 696674 336204 696676
rect 371604 696674 372204 696676
rect 407604 696674 408204 696676
rect 443604 696674 444204 696676
rect 479604 696674 480204 696676
rect 515604 696674 516204 696676
rect 551604 696674 552204 696676
rect 590840 696674 591440 696676
rect -5676 693676 -5076 693678
rect 8004 693676 8604 693678
rect 44004 693676 44604 693678
rect 80004 693676 80604 693678
rect 116004 693676 116604 693678
rect 152004 693676 152604 693678
rect 188004 693676 188604 693678
rect 224004 693676 224604 693678
rect 260004 693676 260604 693678
rect 296004 693676 296604 693678
rect 332004 693676 332604 693678
rect 368004 693676 368604 693678
rect 404004 693676 404604 693678
rect 440004 693676 440604 693678
rect 476004 693676 476604 693678
rect 512004 693676 512604 693678
rect 548004 693676 548604 693678
rect 589000 693676 589600 693678
rect -6596 693654 590520 693676
rect -6596 693418 -5494 693654
rect -5258 693418 8186 693654
rect 8422 693418 44186 693654
rect 44422 693418 80186 693654
rect 80422 693418 116186 693654
rect 116422 693418 152186 693654
rect 152422 693418 188186 693654
rect 188422 693418 224186 693654
rect 224422 693418 260186 693654
rect 260422 693418 296186 693654
rect 296422 693418 332186 693654
rect 332422 693418 368186 693654
rect 368422 693418 404186 693654
rect 404422 693418 440186 693654
rect 440422 693418 476186 693654
rect 476422 693418 512186 693654
rect 512422 693418 548186 693654
rect 548422 693418 589182 693654
rect 589418 693418 590520 693654
rect -6596 693334 590520 693418
rect -6596 693098 -5494 693334
rect -5258 693098 8186 693334
rect 8422 693098 44186 693334
rect 44422 693098 80186 693334
rect 80422 693098 116186 693334
rect 116422 693098 152186 693334
rect 152422 693098 188186 693334
rect 188422 693098 224186 693334
rect 224422 693098 260186 693334
rect 260422 693098 296186 693334
rect 296422 693098 332186 693334
rect 332422 693098 368186 693334
rect 368422 693098 404186 693334
rect 404422 693098 440186 693334
rect 440422 693098 476186 693334
rect 476422 693098 512186 693334
rect 512422 693098 548186 693334
rect 548422 693098 589182 693334
rect 589418 693098 590520 693334
rect -6596 693076 590520 693098
rect -5676 693074 -5076 693076
rect 8004 693074 8604 693076
rect 44004 693074 44604 693076
rect 80004 693074 80604 693076
rect 116004 693074 116604 693076
rect 152004 693074 152604 693076
rect 188004 693074 188604 693076
rect 224004 693074 224604 693076
rect 260004 693074 260604 693076
rect 296004 693074 296604 693076
rect 332004 693074 332604 693076
rect 368004 693074 368604 693076
rect 404004 693074 404604 693076
rect 440004 693074 440604 693076
rect 476004 693074 476604 693076
rect 512004 693074 512604 693076
rect 548004 693074 548604 693076
rect 589000 693074 589600 693076
rect -3836 690076 -3236 690078
rect 4404 690076 5004 690078
rect 40404 690076 41004 690078
rect 76404 690076 77004 690078
rect 112404 690076 113004 690078
rect 148404 690076 149004 690078
rect 184404 690076 185004 690078
rect 220404 690076 221004 690078
rect 256404 690076 257004 690078
rect 292404 690076 293004 690078
rect 328404 690076 329004 690078
rect 364404 690076 365004 690078
rect 400404 690076 401004 690078
rect 436404 690076 437004 690078
rect 472404 690076 473004 690078
rect 508404 690076 509004 690078
rect 544404 690076 545004 690078
rect 580404 690076 581004 690078
rect 587160 690076 587760 690078
rect -4756 690054 588680 690076
rect -4756 689818 -3654 690054
rect -3418 689818 4586 690054
rect 4822 689818 40586 690054
rect 40822 689818 76586 690054
rect 76822 689818 112586 690054
rect 112822 689818 148586 690054
rect 148822 689818 184586 690054
rect 184822 689818 220586 690054
rect 220822 689818 256586 690054
rect 256822 689818 292586 690054
rect 292822 689818 328586 690054
rect 328822 689818 364586 690054
rect 364822 689818 400586 690054
rect 400822 689818 436586 690054
rect 436822 689818 472586 690054
rect 472822 689818 508586 690054
rect 508822 689818 544586 690054
rect 544822 689818 580586 690054
rect 580822 689818 587342 690054
rect 587578 689818 588680 690054
rect -4756 689734 588680 689818
rect -4756 689498 -3654 689734
rect -3418 689498 4586 689734
rect 4822 689498 40586 689734
rect 40822 689498 76586 689734
rect 76822 689498 112586 689734
rect 112822 689498 148586 689734
rect 148822 689498 184586 689734
rect 184822 689498 220586 689734
rect 220822 689498 256586 689734
rect 256822 689498 292586 689734
rect 292822 689498 328586 689734
rect 328822 689498 364586 689734
rect 364822 689498 400586 689734
rect 400822 689498 436586 689734
rect 436822 689498 472586 689734
rect 472822 689498 508586 689734
rect 508822 689498 544586 689734
rect 544822 689498 580586 689734
rect 580822 689498 587342 689734
rect 587578 689498 588680 689734
rect -4756 689476 588680 689498
rect -3836 689474 -3236 689476
rect 4404 689474 5004 689476
rect 40404 689474 41004 689476
rect 76404 689474 77004 689476
rect 112404 689474 113004 689476
rect 148404 689474 149004 689476
rect 184404 689474 185004 689476
rect 220404 689474 221004 689476
rect 256404 689474 257004 689476
rect 292404 689474 293004 689476
rect 328404 689474 329004 689476
rect 364404 689474 365004 689476
rect 400404 689474 401004 689476
rect 436404 689474 437004 689476
rect 472404 689474 473004 689476
rect 508404 689474 509004 689476
rect 544404 689474 545004 689476
rect 580404 689474 581004 689476
rect 587160 689474 587760 689476
rect -1996 686476 -1396 686478
rect 804 686476 1404 686478
rect 36804 686476 37404 686478
rect 72804 686476 73404 686478
rect 108804 686476 109404 686478
rect 144804 686476 145404 686478
rect 180804 686476 181404 686478
rect 216804 686476 217404 686478
rect 252804 686476 253404 686478
rect 288804 686476 289404 686478
rect 324804 686476 325404 686478
rect 360804 686476 361404 686478
rect 396804 686476 397404 686478
rect 432804 686476 433404 686478
rect 468804 686476 469404 686478
rect 504804 686476 505404 686478
rect 540804 686476 541404 686478
rect 576804 686476 577404 686478
rect 585320 686476 585920 686478
rect -2916 686454 586840 686476
rect -2916 686218 -1814 686454
rect -1578 686218 986 686454
rect 1222 686218 36986 686454
rect 37222 686218 72986 686454
rect 73222 686218 108986 686454
rect 109222 686218 144986 686454
rect 145222 686218 180986 686454
rect 181222 686218 216986 686454
rect 217222 686218 252986 686454
rect 253222 686218 288986 686454
rect 289222 686218 324986 686454
rect 325222 686218 360986 686454
rect 361222 686218 396986 686454
rect 397222 686218 432986 686454
rect 433222 686218 468986 686454
rect 469222 686218 504986 686454
rect 505222 686218 540986 686454
rect 541222 686218 576986 686454
rect 577222 686218 585502 686454
rect 585738 686218 586840 686454
rect -2916 686134 586840 686218
rect -2916 685898 -1814 686134
rect -1578 685898 986 686134
rect 1222 685898 36986 686134
rect 37222 685898 72986 686134
rect 73222 685898 108986 686134
rect 109222 685898 144986 686134
rect 145222 685898 180986 686134
rect 181222 685898 216986 686134
rect 217222 685898 252986 686134
rect 253222 685898 288986 686134
rect 289222 685898 324986 686134
rect 325222 685898 360986 686134
rect 361222 685898 396986 686134
rect 397222 685898 432986 686134
rect 433222 685898 468986 686134
rect 469222 685898 504986 686134
rect 505222 685898 540986 686134
rect 541222 685898 576986 686134
rect 577222 685898 585502 686134
rect 585738 685898 586840 686134
rect -2916 685876 586840 685898
rect -1996 685874 -1396 685876
rect 804 685874 1404 685876
rect 36804 685874 37404 685876
rect 72804 685874 73404 685876
rect 108804 685874 109404 685876
rect 144804 685874 145404 685876
rect 180804 685874 181404 685876
rect 216804 685874 217404 685876
rect 252804 685874 253404 685876
rect 288804 685874 289404 685876
rect 324804 685874 325404 685876
rect 360804 685874 361404 685876
rect 396804 685874 397404 685876
rect 432804 685874 433404 685876
rect 468804 685874 469404 685876
rect 504804 685874 505404 685876
rect 540804 685874 541404 685876
rect 576804 685874 577404 685876
rect 585320 685874 585920 685876
rect -8436 679276 -7836 679278
rect 29604 679276 30204 679278
rect 65604 679276 66204 679278
rect 101604 679276 102204 679278
rect 137604 679276 138204 679278
rect 173604 679276 174204 679278
rect 209604 679276 210204 679278
rect 245604 679276 246204 679278
rect 281604 679276 282204 679278
rect 317604 679276 318204 679278
rect 353604 679276 354204 679278
rect 389604 679276 390204 679278
rect 425604 679276 426204 679278
rect 461604 679276 462204 679278
rect 497604 679276 498204 679278
rect 533604 679276 534204 679278
rect 569604 679276 570204 679278
rect 591760 679276 592360 679278
rect -8436 679254 592360 679276
rect -8436 679018 -8254 679254
rect -8018 679018 29786 679254
rect 30022 679018 65786 679254
rect 66022 679018 101786 679254
rect 102022 679018 137786 679254
rect 138022 679018 173786 679254
rect 174022 679018 209786 679254
rect 210022 679018 245786 679254
rect 246022 679018 281786 679254
rect 282022 679018 317786 679254
rect 318022 679018 353786 679254
rect 354022 679018 389786 679254
rect 390022 679018 425786 679254
rect 426022 679018 461786 679254
rect 462022 679018 497786 679254
rect 498022 679018 533786 679254
rect 534022 679018 569786 679254
rect 570022 679018 591942 679254
rect 592178 679018 592360 679254
rect -8436 678934 592360 679018
rect -8436 678698 -8254 678934
rect -8018 678698 29786 678934
rect 30022 678698 65786 678934
rect 66022 678698 101786 678934
rect 102022 678698 137786 678934
rect 138022 678698 173786 678934
rect 174022 678698 209786 678934
rect 210022 678698 245786 678934
rect 246022 678698 281786 678934
rect 282022 678698 317786 678934
rect 318022 678698 353786 678934
rect 354022 678698 389786 678934
rect 390022 678698 425786 678934
rect 426022 678698 461786 678934
rect 462022 678698 497786 678934
rect 498022 678698 533786 678934
rect 534022 678698 569786 678934
rect 570022 678698 591942 678934
rect 592178 678698 592360 678934
rect -8436 678676 592360 678698
rect -8436 678674 -7836 678676
rect 29604 678674 30204 678676
rect 65604 678674 66204 678676
rect 101604 678674 102204 678676
rect 137604 678674 138204 678676
rect 173604 678674 174204 678676
rect 209604 678674 210204 678676
rect 245604 678674 246204 678676
rect 281604 678674 282204 678676
rect 317604 678674 318204 678676
rect 353604 678674 354204 678676
rect 389604 678674 390204 678676
rect 425604 678674 426204 678676
rect 461604 678674 462204 678676
rect 497604 678674 498204 678676
rect 533604 678674 534204 678676
rect 569604 678674 570204 678676
rect 591760 678674 592360 678676
rect -6596 675676 -5996 675678
rect 26004 675676 26604 675678
rect 62004 675676 62604 675678
rect 98004 675676 98604 675678
rect 134004 675676 134604 675678
rect 170004 675676 170604 675678
rect 206004 675676 206604 675678
rect 242004 675676 242604 675678
rect 278004 675676 278604 675678
rect 314004 675676 314604 675678
rect 350004 675676 350604 675678
rect 386004 675676 386604 675678
rect 422004 675676 422604 675678
rect 458004 675676 458604 675678
rect 494004 675676 494604 675678
rect 530004 675676 530604 675678
rect 566004 675676 566604 675678
rect 589920 675676 590520 675678
rect -6596 675654 590520 675676
rect -6596 675418 -6414 675654
rect -6178 675418 26186 675654
rect 26422 675418 62186 675654
rect 62422 675418 98186 675654
rect 98422 675418 134186 675654
rect 134422 675418 170186 675654
rect 170422 675418 206186 675654
rect 206422 675418 242186 675654
rect 242422 675418 278186 675654
rect 278422 675418 314186 675654
rect 314422 675418 350186 675654
rect 350422 675418 386186 675654
rect 386422 675418 422186 675654
rect 422422 675418 458186 675654
rect 458422 675418 494186 675654
rect 494422 675418 530186 675654
rect 530422 675418 566186 675654
rect 566422 675418 590102 675654
rect 590338 675418 590520 675654
rect -6596 675334 590520 675418
rect -6596 675098 -6414 675334
rect -6178 675098 26186 675334
rect 26422 675098 62186 675334
rect 62422 675098 98186 675334
rect 98422 675098 134186 675334
rect 134422 675098 170186 675334
rect 170422 675098 206186 675334
rect 206422 675098 242186 675334
rect 242422 675098 278186 675334
rect 278422 675098 314186 675334
rect 314422 675098 350186 675334
rect 350422 675098 386186 675334
rect 386422 675098 422186 675334
rect 422422 675098 458186 675334
rect 458422 675098 494186 675334
rect 494422 675098 530186 675334
rect 530422 675098 566186 675334
rect 566422 675098 590102 675334
rect 590338 675098 590520 675334
rect -6596 675076 590520 675098
rect -6596 675074 -5996 675076
rect 26004 675074 26604 675076
rect 62004 675074 62604 675076
rect 98004 675074 98604 675076
rect 134004 675074 134604 675076
rect 170004 675074 170604 675076
rect 206004 675074 206604 675076
rect 242004 675074 242604 675076
rect 278004 675074 278604 675076
rect 314004 675074 314604 675076
rect 350004 675074 350604 675076
rect 386004 675074 386604 675076
rect 422004 675074 422604 675076
rect 458004 675074 458604 675076
rect 494004 675074 494604 675076
rect 530004 675074 530604 675076
rect 566004 675074 566604 675076
rect 589920 675074 590520 675076
rect -4756 672076 -4156 672078
rect 22404 672076 23004 672078
rect 58404 672076 59004 672078
rect 94404 672076 95004 672078
rect 130404 672076 131004 672078
rect 166404 672076 167004 672078
rect 202404 672076 203004 672078
rect 238404 672076 239004 672078
rect 274404 672076 275004 672078
rect 310404 672076 311004 672078
rect 346404 672076 347004 672078
rect 382404 672076 383004 672078
rect 418404 672076 419004 672078
rect 454404 672076 455004 672078
rect 490404 672076 491004 672078
rect 526404 672076 527004 672078
rect 562404 672076 563004 672078
rect 588080 672076 588680 672078
rect -4756 672054 588680 672076
rect -4756 671818 -4574 672054
rect -4338 671818 22586 672054
rect 22822 671818 58586 672054
rect 58822 671818 94586 672054
rect 94822 671818 130586 672054
rect 130822 671818 166586 672054
rect 166822 671818 202586 672054
rect 202822 671818 238586 672054
rect 238822 671818 274586 672054
rect 274822 671818 310586 672054
rect 310822 671818 346586 672054
rect 346822 671818 382586 672054
rect 382822 671818 418586 672054
rect 418822 671818 454586 672054
rect 454822 671818 490586 672054
rect 490822 671818 526586 672054
rect 526822 671818 562586 672054
rect 562822 671818 588262 672054
rect 588498 671818 588680 672054
rect -4756 671734 588680 671818
rect -4756 671498 -4574 671734
rect -4338 671498 22586 671734
rect 22822 671498 58586 671734
rect 58822 671498 94586 671734
rect 94822 671498 130586 671734
rect 130822 671498 166586 671734
rect 166822 671498 202586 671734
rect 202822 671498 238586 671734
rect 238822 671498 274586 671734
rect 274822 671498 310586 671734
rect 310822 671498 346586 671734
rect 346822 671498 382586 671734
rect 382822 671498 418586 671734
rect 418822 671498 454586 671734
rect 454822 671498 490586 671734
rect 490822 671498 526586 671734
rect 526822 671498 562586 671734
rect 562822 671498 588262 671734
rect 588498 671498 588680 671734
rect -4756 671476 588680 671498
rect -4756 671474 -4156 671476
rect 22404 671474 23004 671476
rect 58404 671474 59004 671476
rect 94404 671474 95004 671476
rect 130404 671474 131004 671476
rect 166404 671474 167004 671476
rect 202404 671474 203004 671476
rect 238404 671474 239004 671476
rect 274404 671474 275004 671476
rect 310404 671474 311004 671476
rect 346404 671474 347004 671476
rect 382404 671474 383004 671476
rect 418404 671474 419004 671476
rect 454404 671474 455004 671476
rect 490404 671474 491004 671476
rect 526404 671474 527004 671476
rect 562404 671474 563004 671476
rect 588080 671474 588680 671476
rect -2916 668476 -2316 668478
rect 18804 668476 19404 668478
rect 54804 668476 55404 668478
rect 90804 668476 91404 668478
rect 126804 668476 127404 668478
rect 162804 668476 163404 668478
rect 198804 668476 199404 668478
rect 234804 668476 235404 668478
rect 270804 668476 271404 668478
rect 306804 668476 307404 668478
rect 342804 668476 343404 668478
rect 378804 668476 379404 668478
rect 414804 668476 415404 668478
rect 450804 668476 451404 668478
rect 486804 668476 487404 668478
rect 522804 668476 523404 668478
rect 558804 668476 559404 668478
rect 586240 668476 586840 668478
rect -2916 668454 586840 668476
rect -2916 668218 -2734 668454
rect -2498 668218 18986 668454
rect 19222 668218 54986 668454
rect 55222 668218 90986 668454
rect 91222 668218 126986 668454
rect 127222 668218 162986 668454
rect 163222 668218 198986 668454
rect 199222 668218 234986 668454
rect 235222 668218 270986 668454
rect 271222 668218 306986 668454
rect 307222 668218 342986 668454
rect 343222 668218 378986 668454
rect 379222 668218 414986 668454
rect 415222 668218 450986 668454
rect 451222 668218 486986 668454
rect 487222 668218 522986 668454
rect 523222 668218 558986 668454
rect 559222 668218 586422 668454
rect 586658 668218 586840 668454
rect -2916 668134 586840 668218
rect -2916 667898 -2734 668134
rect -2498 667898 18986 668134
rect 19222 667898 54986 668134
rect 55222 667898 90986 668134
rect 91222 667898 126986 668134
rect 127222 667898 162986 668134
rect 163222 667898 198986 668134
rect 199222 667898 234986 668134
rect 235222 667898 270986 668134
rect 271222 667898 306986 668134
rect 307222 667898 342986 668134
rect 343222 667898 378986 668134
rect 379222 667898 414986 668134
rect 415222 667898 450986 668134
rect 451222 667898 486986 668134
rect 487222 667898 522986 668134
rect 523222 667898 558986 668134
rect 559222 667898 586422 668134
rect 586658 667898 586840 668134
rect -2916 667876 586840 667898
rect -2916 667874 -2316 667876
rect 18804 667874 19404 667876
rect 54804 667874 55404 667876
rect 90804 667874 91404 667876
rect 126804 667874 127404 667876
rect 162804 667874 163404 667876
rect 198804 667874 199404 667876
rect 234804 667874 235404 667876
rect 270804 667874 271404 667876
rect 306804 667874 307404 667876
rect 342804 667874 343404 667876
rect 378804 667874 379404 667876
rect 414804 667874 415404 667876
rect 450804 667874 451404 667876
rect 486804 667874 487404 667876
rect 522804 667874 523404 667876
rect 558804 667874 559404 667876
rect 586240 667874 586840 667876
rect -7516 661276 -6916 661278
rect 11604 661276 12204 661278
rect 47604 661276 48204 661278
rect 83604 661276 84204 661278
rect 119604 661276 120204 661278
rect 155604 661276 156204 661278
rect 191604 661276 192204 661278
rect 227604 661276 228204 661278
rect 263604 661276 264204 661278
rect 299604 661276 300204 661278
rect 335604 661276 336204 661278
rect 371604 661276 372204 661278
rect 407604 661276 408204 661278
rect 443604 661276 444204 661278
rect 479604 661276 480204 661278
rect 515604 661276 516204 661278
rect 551604 661276 552204 661278
rect 590840 661276 591440 661278
rect -8436 661254 592360 661276
rect -8436 661018 -7334 661254
rect -7098 661018 11786 661254
rect 12022 661018 47786 661254
rect 48022 661018 83786 661254
rect 84022 661018 119786 661254
rect 120022 661018 155786 661254
rect 156022 661018 191786 661254
rect 192022 661018 227786 661254
rect 228022 661018 263786 661254
rect 264022 661018 299786 661254
rect 300022 661018 335786 661254
rect 336022 661018 371786 661254
rect 372022 661018 407786 661254
rect 408022 661018 443786 661254
rect 444022 661018 479786 661254
rect 480022 661018 515786 661254
rect 516022 661018 551786 661254
rect 552022 661018 591022 661254
rect 591258 661018 592360 661254
rect -8436 660934 592360 661018
rect -8436 660698 -7334 660934
rect -7098 660698 11786 660934
rect 12022 660698 47786 660934
rect 48022 660698 83786 660934
rect 84022 660698 119786 660934
rect 120022 660698 155786 660934
rect 156022 660698 191786 660934
rect 192022 660698 227786 660934
rect 228022 660698 263786 660934
rect 264022 660698 299786 660934
rect 300022 660698 335786 660934
rect 336022 660698 371786 660934
rect 372022 660698 407786 660934
rect 408022 660698 443786 660934
rect 444022 660698 479786 660934
rect 480022 660698 515786 660934
rect 516022 660698 551786 660934
rect 552022 660698 591022 660934
rect 591258 660698 592360 660934
rect -8436 660676 592360 660698
rect -7516 660674 -6916 660676
rect 11604 660674 12204 660676
rect 47604 660674 48204 660676
rect 83604 660674 84204 660676
rect 119604 660674 120204 660676
rect 155604 660674 156204 660676
rect 191604 660674 192204 660676
rect 227604 660674 228204 660676
rect 263604 660674 264204 660676
rect 299604 660674 300204 660676
rect 335604 660674 336204 660676
rect 371604 660674 372204 660676
rect 407604 660674 408204 660676
rect 443604 660674 444204 660676
rect 479604 660674 480204 660676
rect 515604 660674 516204 660676
rect 551604 660674 552204 660676
rect 590840 660674 591440 660676
rect -5676 657676 -5076 657678
rect 8004 657676 8604 657678
rect 44004 657676 44604 657678
rect 80004 657676 80604 657678
rect 116004 657676 116604 657678
rect 152004 657676 152604 657678
rect 188004 657676 188604 657678
rect 224004 657676 224604 657678
rect 260004 657676 260604 657678
rect 296004 657676 296604 657678
rect 332004 657676 332604 657678
rect 368004 657676 368604 657678
rect 404004 657676 404604 657678
rect 440004 657676 440604 657678
rect 476004 657676 476604 657678
rect 512004 657676 512604 657678
rect 548004 657676 548604 657678
rect 589000 657676 589600 657678
rect -6596 657654 590520 657676
rect -6596 657418 -5494 657654
rect -5258 657418 8186 657654
rect 8422 657418 44186 657654
rect 44422 657418 80186 657654
rect 80422 657418 116186 657654
rect 116422 657418 152186 657654
rect 152422 657418 188186 657654
rect 188422 657418 224186 657654
rect 224422 657418 260186 657654
rect 260422 657418 296186 657654
rect 296422 657418 332186 657654
rect 332422 657418 368186 657654
rect 368422 657418 404186 657654
rect 404422 657418 440186 657654
rect 440422 657418 476186 657654
rect 476422 657418 512186 657654
rect 512422 657418 548186 657654
rect 548422 657418 589182 657654
rect 589418 657418 590520 657654
rect -6596 657334 590520 657418
rect -6596 657098 -5494 657334
rect -5258 657098 8186 657334
rect 8422 657098 44186 657334
rect 44422 657098 80186 657334
rect 80422 657098 116186 657334
rect 116422 657098 152186 657334
rect 152422 657098 188186 657334
rect 188422 657098 224186 657334
rect 224422 657098 260186 657334
rect 260422 657098 296186 657334
rect 296422 657098 332186 657334
rect 332422 657098 368186 657334
rect 368422 657098 404186 657334
rect 404422 657098 440186 657334
rect 440422 657098 476186 657334
rect 476422 657098 512186 657334
rect 512422 657098 548186 657334
rect 548422 657098 589182 657334
rect 589418 657098 590520 657334
rect -6596 657076 590520 657098
rect -5676 657074 -5076 657076
rect 8004 657074 8604 657076
rect 44004 657074 44604 657076
rect 80004 657074 80604 657076
rect 116004 657074 116604 657076
rect 152004 657074 152604 657076
rect 188004 657074 188604 657076
rect 224004 657074 224604 657076
rect 260004 657074 260604 657076
rect 296004 657074 296604 657076
rect 332004 657074 332604 657076
rect 368004 657074 368604 657076
rect 404004 657074 404604 657076
rect 440004 657074 440604 657076
rect 476004 657074 476604 657076
rect 512004 657074 512604 657076
rect 548004 657074 548604 657076
rect 589000 657074 589600 657076
rect -3836 654076 -3236 654078
rect 4404 654076 5004 654078
rect 40404 654076 41004 654078
rect 76404 654076 77004 654078
rect 112404 654076 113004 654078
rect 148404 654076 149004 654078
rect 184404 654076 185004 654078
rect 220404 654076 221004 654078
rect 256404 654076 257004 654078
rect 292404 654076 293004 654078
rect 328404 654076 329004 654078
rect 364404 654076 365004 654078
rect 400404 654076 401004 654078
rect 436404 654076 437004 654078
rect 472404 654076 473004 654078
rect 508404 654076 509004 654078
rect 544404 654076 545004 654078
rect 580404 654076 581004 654078
rect 587160 654076 587760 654078
rect -4756 654054 588680 654076
rect -4756 653818 -3654 654054
rect -3418 653818 4586 654054
rect 4822 653818 40586 654054
rect 40822 653818 76586 654054
rect 76822 653818 112586 654054
rect 112822 653818 148586 654054
rect 148822 653818 184586 654054
rect 184822 653818 220586 654054
rect 220822 653818 256586 654054
rect 256822 653818 292586 654054
rect 292822 653818 328586 654054
rect 328822 653818 364586 654054
rect 364822 653818 400586 654054
rect 400822 653818 436586 654054
rect 436822 653818 472586 654054
rect 472822 653818 508586 654054
rect 508822 653818 544586 654054
rect 544822 653818 580586 654054
rect 580822 653818 587342 654054
rect 587578 653818 588680 654054
rect -4756 653734 588680 653818
rect -4756 653498 -3654 653734
rect -3418 653498 4586 653734
rect 4822 653498 40586 653734
rect 40822 653498 76586 653734
rect 76822 653498 112586 653734
rect 112822 653498 148586 653734
rect 148822 653498 184586 653734
rect 184822 653498 220586 653734
rect 220822 653498 256586 653734
rect 256822 653498 292586 653734
rect 292822 653498 328586 653734
rect 328822 653498 364586 653734
rect 364822 653498 400586 653734
rect 400822 653498 436586 653734
rect 436822 653498 472586 653734
rect 472822 653498 508586 653734
rect 508822 653498 544586 653734
rect 544822 653498 580586 653734
rect 580822 653498 587342 653734
rect 587578 653498 588680 653734
rect -4756 653476 588680 653498
rect -3836 653474 -3236 653476
rect 4404 653474 5004 653476
rect 40404 653474 41004 653476
rect 76404 653474 77004 653476
rect 112404 653474 113004 653476
rect 148404 653474 149004 653476
rect 184404 653474 185004 653476
rect 220404 653474 221004 653476
rect 256404 653474 257004 653476
rect 292404 653474 293004 653476
rect 328404 653474 329004 653476
rect 364404 653474 365004 653476
rect 400404 653474 401004 653476
rect 436404 653474 437004 653476
rect 472404 653474 473004 653476
rect 508404 653474 509004 653476
rect 544404 653474 545004 653476
rect 580404 653474 581004 653476
rect 587160 653474 587760 653476
rect -1996 650476 -1396 650478
rect 804 650476 1404 650478
rect 36804 650476 37404 650478
rect 72804 650476 73404 650478
rect 108804 650476 109404 650478
rect 144804 650476 145404 650478
rect 180804 650476 181404 650478
rect 216804 650476 217404 650478
rect 252804 650476 253404 650478
rect 288804 650476 289404 650478
rect 324804 650476 325404 650478
rect 360804 650476 361404 650478
rect 396804 650476 397404 650478
rect 432804 650476 433404 650478
rect 468804 650476 469404 650478
rect 504804 650476 505404 650478
rect 540804 650476 541404 650478
rect 576804 650476 577404 650478
rect 585320 650476 585920 650478
rect -2916 650454 586840 650476
rect -2916 650218 -1814 650454
rect -1578 650218 986 650454
rect 1222 650218 36986 650454
rect 37222 650218 72986 650454
rect 73222 650218 108986 650454
rect 109222 650218 144986 650454
rect 145222 650218 180986 650454
rect 181222 650218 216986 650454
rect 217222 650218 252986 650454
rect 253222 650218 288986 650454
rect 289222 650218 324986 650454
rect 325222 650218 360986 650454
rect 361222 650218 396986 650454
rect 397222 650218 432986 650454
rect 433222 650218 468986 650454
rect 469222 650218 504986 650454
rect 505222 650218 540986 650454
rect 541222 650218 576986 650454
rect 577222 650218 585502 650454
rect 585738 650218 586840 650454
rect -2916 650134 586840 650218
rect -2916 649898 -1814 650134
rect -1578 649898 986 650134
rect 1222 649898 36986 650134
rect 37222 649898 72986 650134
rect 73222 649898 108986 650134
rect 109222 649898 144986 650134
rect 145222 649898 180986 650134
rect 181222 649898 216986 650134
rect 217222 649898 252986 650134
rect 253222 649898 288986 650134
rect 289222 649898 324986 650134
rect 325222 649898 360986 650134
rect 361222 649898 396986 650134
rect 397222 649898 432986 650134
rect 433222 649898 468986 650134
rect 469222 649898 504986 650134
rect 505222 649898 540986 650134
rect 541222 649898 576986 650134
rect 577222 649898 585502 650134
rect 585738 649898 586840 650134
rect -2916 649876 586840 649898
rect -1996 649874 -1396 649876
rect 804 649874 1404 649876
rect 36804 649874 37404 649876
rect 72804 649874 73404 649876
rect 108804 649874 109404 649876
rect 144804 649874 145404 649876
rect 180804 649874 181404 649876
rect 216804 649874 217404 649876
rect 252804 649874 253404 649876
rect 288804 649874 289404 649876
rect 324804 649874 325404 649876
rect 360804 649874 361404 649876
rect 396804 649874 397404 649876
rect 432804 649874 433404 649876
rect 468804 649874 469404 649876
rect 504804 649874 505404 649876
rect 540804 649874 541404 649876
rect 576804 649874 577404 649876
rect 585320 649874 585920 649876
rect -8436 643276 -7836 643278
rect 29604 643276 30204 643278
rect 65604 643276 66204 643278
rect 101604 643276 102204 643278
rect 137604 643276 138204 643278
rect 173604 643276 174204 643278
rect 209604 643276 210204 643278
rect 245604 643276 246204 643278
rect 281604 643276 282204 643278
rect 317604 643276 318204 643278
rect 353604 643276 354204 643278
rect 389604 643276 390204 643278
rect 425604 643276 426204 643278
rect 461604 643276 462204 643278
rect 497604 643276 498204 643278
rect 533604 643276 534204 643278
rect 569604 643276 570204 643278
rect 591760 643276 592360 643278
rect -8436 643254 592360 643276
rect -8436 643018 -8254 643254
rect -8018 643018 29786 643254
rect 30022 643018 65786 643254
rect 66022 643018 101786 643254
rect 102022 643018 137786 643254
rect 138022 643018 173786 643254
rect 174022 643018 209786 643254
rect 210022 643018 245786 643254
rect 246022 643018 281786 643254
rect 282022 643018 317786 643254
rect 318022 643018 353786 643254
rect 354022 643018 389786 643254
rect 390022 643018 425786 643254
rect 426022 643018 461786 643254
rect 462022 643018 497786 643254
rect 498022 643018 533786 643254
rect 534022 643018 569786 643254
rect 570022 643018 591942 643254
rect 592178 643018 592360 643254
rect -8436 642934 592360 643018
rect -8436 642698 -8254 642934
rect -8018 642698 29786 642934
rect 30022 642698 65786 642934
rect 66022 642698 101786 642934
rect 102022 642698 137786 642934
rect 138022 642698 173786 642934
rect 174022 642698 209786 642934
rect 210022 642698 245786 642934
rect 246022 642698 281786 642934
rect 282022 642698 317786 642934
rect 318022 642698 353786 642934
rect 354022 642698 389786 642934
rect 390022 642698 425786 642934
rect 426022 642698 461786 642934
rect 462022 642698 497786 642934
rect 498022 642698 533786 642934
rect 534022 642698 569786 642934
rect 570022 642698 591942 642934
rect 592178 642698 592360 642934
rect -8436 642676 592360 642698
rect -8436 642674 -7836 642676
rect 29604 642674 30204 642676
rect 65604 642674 66204 642676
rect 101604 642674 102204 642676
rect 137604 642674 138204 642676
rect 173604 642674 174204 642676
rect 209604 642674 210204 642676
rect 245604 642674 246204 642676
rect 281604 642674 282204 642676
rect 317604 642674 318204 642676
rect 353604 642674 354204 642676
rect 389604 642674 390204 642676
rect 425604 642674 426204 642676
rect 461604 642674 462204 642676
rect 497604 642674 498204 642676
rect 533604 642674 534204 642676
rect 569604 642674 570204 642676
rect 591760 642674 592360 642676
rect -6596 639676 -5996 639678
rect 26004 639676 26604 639678
rect 62004 639676 62604 639678
rect 98004 639676 98604 639678
rect 134004 639676 134604 639678
rect 170004 639676 170604 639678
rect 206004 639676 206604 639678
rect 242004 639676 242604 639678
rect 278004 639676 278604 639678
rect 314004 639676 314604 639678
rect 350004 639676 350604 639678
rect 386004 639676 386604 639678
rect 422004 639676 422604 639678
rect 458004 639676 458604 639678
rect 494004 639676 494604 639678
rect 530004 639676 530604 639678
rect 566004 639676 566604 639678
rect 589920 639676 590520 639678
rect -6596 639654 590520 639676
rect -6596 639418 -6414 639654
rect -6178 639418 26186 639654
rect 26422 639418 62186 639654
rect 62422 639418 98186 639654
rect 98422 639418 134186 639654
rect 134422 639418 170186 639654
rect 170422 639418 206186 639654
rect 206422 639418 242186 639654
rect 242422 639418 278186 639654
rect 278422 639418 314186 639654
rect 314422 639418 350186 639654
rect 350422 639418 386186 639654
rect 386422 639418 422186 639654
rect 422422 639418 458186 639654
rect 458422 639418 494186 639654
rect 494422 639418 530186 639654
rect 530422 639418 566186 639654
rect 566422 639418 590102 639654
rect 590338 639418 590520 639654
rect -6596 639334 590520 639418
rect -6596 639098 -6414 639334
rect -6178 639098 26186 639334
rect 26422 639098 62186 639334
rect 62422 639098 98186 639334
rect 98422 639098 134186 639334
rect 134422 639098 170186 639334
rect 170422 639098 206186 639334
rect 206422 639098 242186 639334
rect 242422 639098 278186 639334
rect 278422 639098 314186 639334
rect 314422 639098 350186 639334
rect 350422 639098 386186 639334
rect 386422 639098 422186 639334
rect 422422 639098 458186 639334
rect 458422 639098 494186 639334
rect 494422 639098 530186 639334
rect 530422 639098 566186 639334
rect 566422 639098 590102 639334
rect 590338 639098 590520 639334
rect -6596 639076 590520 639098
rect -6596 639074 -5996 639076
rect 26004 639074 26604 639076
rect 62004 639074 62604 639076
rect 98004 639074 98604 639076
rect 134004 639074 134604 639076
rect 170004 639074 170604 639076
rect 206004 639074 206604 639076
rect 242004 639074 242604 639076
rect 278004 639074 278604 639076
rect 314004 639074 314604 639076
rect 350004 639074 350604 639076
rect 386004 639074 386604 639076
rect 422004 639074 422604 639076
rect 458004 639074 458604 639076
rect 494004 639074 494604 639076
rect 530004 639074 530604 639076
rect 566004 639074 566604 639076
rect 589920 639074 590520 639076
rect -4756 636076 -4156 636078
rect 22404 636076 23004 636078
rect 58404 636076 59004 636078
rect 94404 636076 95004 636078
rect 130404 636076 131004 636078
rect 166404 636076 167004 636078
rect 202404 636076 203004 636078
rect 238404 636076 239004 636078
rect 274404 636076 275004 636078
rect 310404 636076 311004 636078
rect 346404 636076 347004 636078
rect 382404 636076 383004 636078
rect 418404 636076 419004 636078
rect 454404 636076 455004 636078
rect 490404 636076 491004 636078
rect 526404 636076 527004 636078
rect 562404 636076 563004 636078
rect 588080 636076 588680 636078
rect -4756 636054 588680 636076
rect -4756 635818 -4574 636054
rect -4338 635818 22586 636054
rect 22822 635818 58586 636054
rect 58822 635818 94586 636054
rect 94822 635818 130586 636054
rect 130822 635818 166586 636054
rect 166822 635818 202586 636054
rect 202822 635818 238586 636054
rect 238822 635818 274586 636054
rect 274822 635818 310586 636054
rect 310822 635818 346586 636054
rect 346822 635818 382586 636054
rect 382822 635818 418586 636054
rect 418822 635818 454586 636054
rect 454822 635818 490586 636054
rect 490822 635818 526586 636054
rect 526822 635818 562586 636054
rect 562822 635818 588262 636054
rect 588498 635818 588680 636054
rect -4756 635734 588680 635818
rect -4756 635498 -4574 635734
rect -4338 635498 22586 635734
rect 22822 635498 58586 635734
rect 58822 635498 94586 635734
rect 94822 635498 130586 635734
rect 130822 635498 166586 635734
rect 166822 635498 202586 635734
rect 202822 635498 238586 635734
rect 238822 635498 274586 635734
rect 274822 635498 310586 635734
rect 310822 635498 346586 635734
rect 346822 635498 382586 635734
rect 382822 635498 418586 635734
rect 418822 635498 454586 635734
rect 454822 635498 490586 635734
rect 490822 635498 526586 635734
rect 526822 635498 562586 635734
rect 562822 635498 588262 635734
rect 588498 635498 588680 635734
rect -4756 635476 588680 635498
rect -4756 635474 -4156 635476
rect 22404 635474 23004 635476
rect 58404 635474 59004 635476
rect 94404 635474 95004 635476
rect 130404 635474 131004 635476
rect 166404 635474 167004 635476
rect 202404 635474 203004 635476
rect 238404 635474 239004 635476
rect 274404 635474 275004 635476
rect 310404 635474 311004 635476
rect 346404 635474 347004 635476
rect 382404 635474 383004 635476
rect 418404 635474 419004 635476
rect 454404 635474 455004 635476
rect 490404 635474 491004 635476
rect 526404 635474 527004 635476
rect 562404 635474 563004 635476
rect 588080 635474 588680 635476
rect -2916 632476 -2316 632478
rect 18804 632476 19404 632478
rect 54804 632476 55404 632478
rect 90804 632476 91404 632478
rect 126804 632476 127404 632478
rect 162804 632476 163404 632478
rect 198804 632476 199404 632478
rect 234804 632476 235404 632478
rect 270804 632476 271404 632478
rect 306804 632476 307404 632478
rect 342804 632476 343404 632478
rect 378804 632476 379404 632478
rect 414804 632476 415404 632478
rect 450804 632476 451404 632478
rect 486804 632476 487404 632478
rect 522804 632476 523404 632478
rect 558804 632476 559404 632478
rect 586240 632476 586840 632478
rect -2916 632454 586840 632476
rect -2916 632218 -2734 632454
rect -2498 632218 18986 632454
rect 19222 632218 54986 632454
rect 55222 632218 90986 632454
rect 91222 632218 126986 632454
rect 127222 632218 162986 632454
rect 163222 632218 198986 632454
rect 199222 632218 234986 632454
rect 235222 632218 270986 632454
rect 271222 632218 306986 632454
rect 307222 632218 342986 632454
rect 343222 632218 378986 632454
rect 379222 632218 414986 632454
rect 415222 632218 450986 632454
rect 451222 632218 486986 632454
rect 487222 632218 522986 632454
rect 523222 632218 558986 632454
rect 559222 632218 586422 632454
rect 586658 632218 586840 632454
rect -2916 632134 586840 632218
rect -2916 631898 -2734 632134
rect -2498 631898 18986 632134
rect 19222 631898 54986 632134
rect 55222 631898 90986 632134
rect 91222 631898 126986 632134
rect 127222 631898 162986 632134
rect 163222 631898 198986 632134
rect 199222 631898 234986 632134
rect 235222 631898 270986 632134
rect 271222 631898 306986 632134
rect 307222 631898 342986 632134
rect 343222 631898 378986 632134
rect 379222 631898 414986 632134
rect 415222 631898 450986 632134
rect 451222 631898 486986 632134
rect 487222 631898 522986 632134
rect 523222 631898 558986 632134
rect 559222 631898 586422 632134
rect 586658 631898 586840 632134
rect -2916 631876 586840 631898
rect -2916 631874 -2316 631876
rect 18804 631874 19404 631876
rect 54804 631874 55404 631876
rect 90804 631874 91404 631876
rect 126804 631874 127404 631876
rect 162804 631874 163404 631876
rect 198804 631874 199404 631876
rect 234804 631874 235404 631876
rect 270804 631874 271404 631876
rect 306804 631874 307404 631876
rect 342804 631874 343404 631876
rect 378804 631874 379404 631876
rect 414804 631874 415404 631876
rect 450804 631874 451404 631876
rect 486804 631874 487404 631876
rect 522804 631874 523404 631876
rect 558804 631874 559404 631876
rect 586240 631874 586840 631876
rect -7516 625276 -6916 625278
rect 11604 625276 12204 625278
rect 47604 625276 48204 625278
rect 83604 625276 84204 625278
rect 119604 625276 120204 625278
rect 155604 625276 156204 625278
rect 191604 625276 192204 625278
rect 227604 625276 228204 625278
rect 263604 625276 264204 625278
rect 299604 625276 300204 625278
rect 335604 625276 336204 625278
rect 371604 625276 372204 625278
rect 407604 625276 408204 625278
rect 443604 625276 444204 625278
rect 479604 625276 480204 625278
rect 515604 625276 516204 625278
rect 551604 625276 552204 625278
rect 590840 625276 591440 625278
rect -8436 625254 592360 625276
rect -8436 625018 -7334 625254
rect -7098 625018 11786 625254
rect 12022 625018 47786 625254
rect 48022 625018 83786 625254
rect 84022 625018 119786 625254
rect 120022 625018 155786 625254
rect 156022 625018 191786 625254
rect 192022 625018 227786 625254
rect 228022 625018 263786 625254
rect 264022 625018 299786 625254
rect 300022 625018 335786 625254
rect 336022 625018 371786 625254
rect 372022 625018 407786 625254
rect 408022 625018 443786 625254
rect 444022 625018 479786 625254
rect 480022 625018 515786 625254
rect 516022 625018 551786 625254
rect 552022 625018 591022 625254
rect 591258 625018 592360 625254
rect -8436 624934 592360 625018
rect -8436 624698 -7334 624934
rect -7098 624698 11786 624934
rect 12022 624698 47786 624934
rect 48022 624698 83786 624934
rect 84022 624698 119786 624934
rect 120022 624698 155786 624934
rect 156022 624698 191786 624934
rect 192022 624698 227786 624934
rect 228022 624698 263786 624934
rect 264022 624698 299786 624934
rect 300022 624698 335786 624934
rect 336022 624698 371786 624934
rect 372022 624698 407786 624934
rect 408022 624698 443786 624934
rect 444022 624698 479786 624934
rect 480022 624698 515786 624934
rect 516022 624698 551786 624934
rect 552022 624698 591022 624934
rect 591258 624698 592360 624934
rect -8436 624676 592360 624698
rect -7516 624674 -6916 624676
rect 11604 624674 12204 624676
rect 47604 624674 48204 624676
rect 83604 624674 84204 624676
rect 119604 624674 120204 624676
rect 155604 624674 156204 624676
rect 191604 624674 192204 624676
rect 227604 624674 228204 624676
rect 263604 624674 264204 624676
rect 299604 624674 300204 624676
rect 335604 624674 336204 624676
rect 371604 624674 372204 624676
rect 407604 624674 408204 624676
rect 443604 624674 444204 624676
rect 479604 624674 480204 624676
rect 515604 624674 516204 624676
rect 551604 624674 552204 624676
rect 590840 624674 591440 624676
rect -5676 621676 -5076 621678
rect 8004 621676 8604 621678
rect 44004 621676 44604 621678
rect 80004 621676 80604 621678
rect 116004 621676 116604 621678
rect 152004 621676 152604 621678
rect 188004 621676 188604 621678
rect 224004 621676 224604 621678
rect 260004 621676 260604 621678
rect 296004 621676 296604 621678
rect 332004 621676 332604 621678
rect 368004 621676 368604 621678
rect 404004 621676 404604 621678
rect 440004 621676 440604 621678
rect 476004 621676 476604 621678
rect 512004 621676 512604 621678
rect 548004 621676 548604 621678
rect 589000 621676 589600 621678
rect -6596 621654 590520 621676
rect -6596 621418 -5494 621654
rect -5258 621418 8186 621654
rect 8422 621418 44186 621654
rect 44422 621418 80186 621654
rect 80422 621418 116186 621654
rect 116422 621418 152186 621654
rect 152422 621418 188186 621654
rect 188422 621418 224186 621654
rect 224422 621418 260186 621654
rect 260422 621418 296186 621654
rect 296422 621418 332186 621654
rect 332422 621418 368186 621654
rect 368422 621418 404186 621654
rect 404422 621418 440186 621654
rect 440422 621418 476186 621654
rect 476422 621418 512186 621654
rect 512422 621418 548186 621654
rect 548422 621418 589182 621654
rect 589418 621418 590520 621654
rect -6596 621334 590520 621418
rect -6596 621098 -5494 621334
rect -5258 621098 8186 621334
rect 8422 621098 44186 621334
rect 44422 621098 80186 621334
rect 80422 621098 116186 621334
rect 116422 621098 152186 621334
rect 152422 621098 188186 621334
rect 188422 621098 224186 621334
rect 224422 621098 260186 621334
rect 260422 621098 296186 621334
rect 296422 621098 332186 621334
rect 332422 621098 368186 621334
rect 368422 621098 404186 621334
rect 404422 621098 440186 621334
rect 440422 621098 476186 621334
rect 476422 621098 512186 621334
rect 512422 621098 548186 621334
rect 548422 621098 589182 621334
rect 589418 621098 590520 621334
rect -6596 621076 590520 621098
rect -5676 621074 -5076 621076
rect 8004 621074 8604 621076
rect 44004 621074 44604 621076
rect 80004 621074 80604 621076
rect 116004 621074 116604 621076
rect 152004 621074 152604 621076
rect 188004 621074 188604 621076
rect 224004 621074 224604 621076
rect 260004 621074 260604 621076
rect 296004 621074 296604 621076
rect 332004 621074 332604 621076
rect 368004 621074 368604 621076
rect 404004 621074 404604 621076
rect 440004 621074 440604 621076
rect 476004 621074 476604 621076
rect 512004 621074 512604 621076
rect 548004 621074 548604 621076
rect 589000 621074 589600 621076
rect -3836 618076 -3236 618078
rect 4404 618076 5004 618078
rect 40404 618076 41004 618078
rect 76404 618076 77004 618078
rect 112404 618076 113004 618078
rect 148404 618076 149004 618078
rect 184404 618076 185004 618078
rect 220404 618076 221004 618078
rect 256404 618076 257004 618078
rect 292404 618076 293004 618078
rect 328404 618076 329004 618078
rect 364404 618076 365004 618078
rect 400404 618076 401004 618078
rect 436404 618076 437004 618078
rect 472404 618076 473004 618078
rect 508404 618076 509004 618078
rect 544404 618076 545004 618078
rect 580404 618076 581004 618078
rect 587160 618076 587760 618078
rect -4756 618054 588680 618076
rect -4756 617818 -3654 618054
rect -3418 617818 4586 618054
rect 4822 617818 40586 618054
rect 40822 617818 76586 618054
rect 76822 617818 112586 618054
rect 112822 617818 148586 618054
rect 148822 617818 184586 618054
rect 184822 617818 220586 618054
rect 220822 617818 256586 618054
rect 256822 617818 292586 618054
rect 292822 617818 328586 618054
rect 328822 617818 364586 618054
rect 364822 617818 400586 618054
rect 400822 617818 436586 618054
rect 436822 617818 472586 618054
rect 472822 617818 508586 618054
rect 508822 617818 544586 618054
rect 544822 617818 580586 618054
rect 580822 617818 587342 618054
rect 587578 617818 588680 618054
rect -4756 617734 588680 617818
rect -4756 617498 -3654 617734
rect -3418 617498 4586 617734
rect 4822 617498 40586 617734
rect 40822 617498 76586 617734
rect 76822 617498 112586 617734
rect 112822 617498 148586 617734
rect 148822 617498 184586 617734
rect 184822 617498 220586 617734
rect 220822 617498 256586 617734
rect 256822 617498 292586 617734
rect 292822 617498 328586 617734
rect 328822 617498 364586 617734
rect 364822 617498 400586 617734
rect 400822 617498 436586 617734
rect 436822 617498 472586 617734
rect 472822 617498 508586 617734
rect 508822 617498 544586 617734
rect 544822 617498 580586 617734
rect 580822 617498 587342 617734
rect 587578 617498 588680 617734
rect -4756 617476 588680 617498
rect -3836 617474 -3236 617476
rect 4404 617474 5004 617476
rect 40404 617474 41004 617476
rect 76404 617474 77004 617476
rect 112404 617474 113004 617476
rect 148404 617474 149004 617476
rect 184404 617474 185004 617476
rect 220404 617474 221004 617476
rect 256404 617474 257004 617476
rect 292404 617474 293004 617476
rect 328404 617474 329004 617476
rect 364404 617474 365004 617476
rect 400404 617474 401004 617476
rect 436404 617474 437004 617476
rect 472404 617474 473004 617476
rect 508404 617474 509004 617476
rect 544404 617474 545004 617476
rect 580404 617474 581004 617476
rect 587160 617474 587760 617476
rect -1996 614476 -1396 614478
rect 804 614476 1404 614478
rect 36804 614476 37404 614478
rect 72804 614476 73404 614478
rect 108804 614476 109404 614478
rect 144804 614476 145404 614478
rect 180804 614476 181404 614478
rect 216804 614476 217404 614478
rect 252804 614476 253404 614478
rect 288804 614476 289404 614478
rect 324804 614476 325404 614478
rect 360804 614476 361404 614478
rect 396804 614476 397404 614478
rect 432804 614476 433404 614478
rect 468804 614476 469404 614478
rect 504804 614476 505404 614478
rect 540804 614476 541404 614478
rect 576804 614476 577404 614478
rect 585320 614476 585920 614478
rect -2916 614454 586840 614476
rect -2916 614218 -1814 614454
rect -1578 614218 986 614454
rect 1222 614218 36986 614454
rect 37222 614218 72986 614454
rect 73222 614218 108986 614454
rect 109222 614218 144986 614454
rect 145222 614218 180986 614454
rect 181222 614218 216986 614454
rect 217222 614218 252986 614454
rect 253222 614218 288986 614454
rect 289222 614218 324986 614454
rect 325222 614218 360986 614454
rect 361222 614218 396986 614454
rect 397222 614218 432986 614454
rect 433222 614218 468986 614454
rect 469222 614218 504986 614454
rect 505222 614218 540986 614454
rect 541222 614218 576986 614454
rect 577222 614218 585502 614454
rect 585738 614218 586840 614454
rect -2916 614134 586840 614218
rect -2916 613898 -1814 614134
rect -1578 613898 986 614134
rect 1222 613898 36986 614134
rect 37222 613898 72986 614134
rect 73222 613898 108986 614134
rect 109222 613898 144986 614134
rect 145222 613898 180986 614134
rect 181222 613898 216986 614134
rect 217222 613898 252986 614134
rect 253222 613898 288986 614134
rect 289222 613898 324986 614134
rect 325222 613898 360986 614134
rect 361222 613898 396986 614134
rect 397222 613898 432986 614134
rect 433222 613898 468986 614134
rect 469222 613898 504986 614134
rect 505222 613898 540986 614134
rect 541222 613898 576986 614134
rect 577222 613898 585502 614134
rect 585738 613898 586840 614134
rect -2916 613876 586840 613898
rect -1996 613874 -1396 613876
rect 804 613874 1404 613876
rect 36804 613874 37404 613876
rect 72804 613874 73404 613876
rect 108804 613874 109404 613876
rect 144804 613874 145404 613876
rect 180804 613874 181404 613876
rect 216804 613874 217404 613876
rect 252804 613874 253404 613876
rect 288804 613874 289404 613876
rect 324804 613874 325404 613876
rect 360804 613874 361404 613876
rect 396804 613874 397404 613876
rect 432804 613874 433404 613876
rect 468804 613874 469404 613876
rect 504804 613874 505404 613876
rect 540804 613874 541404 613876
rect 576804 613874 577404 613876
rect 585320 613874 585920 613876
rect -8436 607276 -7836 607278
rect 29604 607276 30204 607278
rect 65604 607276 66204 607278
rect 101604 607276 102204 607278
rect 137604 607276 138204 607278
rect 173604 607276 174204 607278
rect 209604 607276 210204 607278
rect 245604 607276 246204 607278
rect 281604 607276 282204 607278
rect 317604 607276 318204 607278
rect 353604 607276 354204 607278
rect 389604 607276 390204 607278
rect 425604 607276 426204 607278
rect 461604 607276 462204 607278
rect 497604 607276 498204 607278
rect 533604 607276 534204 607278
rect 569604 607276 570204 607278
rect 591760 607276 592360 607278
rect -8436 607254 592360 607276
rect -8436 607018 -8254 607254
rect -8018 607018 29786 607254
rect 30022 607018 65786 607254
rect 66022 607018 101786 607254
rect 102022 607018 137786 607254
rect 138022 607018 173786 607254
rect 174022 607018 209786 607254
rect 210022 607018 245786 607254
rect 246022 607018 281786 607254
rect 282022 607018 317786 607254
rect 318022 607018 353786 607254
rect 354022 607018 389786 607254
rect 390022 607018 425786 607254
rect 426022 607018 461786 607254
rect 462022 607018 497786 607254
rect 498022 607018 533786 607254
rect 534022 607018 569786 607254
rect 570022 607018 591942 607254
rect 592178 607018 592360 607254
rect -8436 606934 592360 607018
rect -8436 606698 -8254 606934
rect -8018 606698 29786 606934
rect 30022 606698 65786 606934
rect 66022 606698 101786 606934
rect 102022 606698 137786 606934
rect 138022 606698 173786 606934
rect 174022 606698 209786 606934
rect 210022 606698 245786 606934
rect 246022 606698 281786 606934
rect 282022 606698 317786 606934
rect 318022 606698 353786 606934
rect 354022 606698 389786 606934
rect 390022 606698 425786 606934
rect 426022 606698 461786 606934
rect 462022 606698 497786 606934
rect 498022 606698 533786 606934
rect 534022 606698 569786 606934
rect 570022 606698 591942 606934
rect 592178 606698 592360 606934
rect -8436 606676 592360 606698
rect -8436 606674 -7836 606676
rect 29604 606674 30204 606676
rect 65604 606674 66204 606676
rect 101604 606674 102204 606676
rect 137604 606674 138204 606676
rect 173604 606674 174204 606676
rect 209604 606674 210204 606676
rect 245604 606674 246204 606676
rect 281604 606674 282204 606676
rect 317604 606674 318204 606676
rect 353604 606674 354204 606676
rect 389604 606674 390204 606676
rect 425604 606674 426204 606676
rect 461604 606674 462204 606676
rect 497604 606674 498204 606676
rect 533604 606674 534204 606676
rect 569604 606674 570204 606676
rect 591760 606674 592360 606676
rect -6596 603676 -5996 603678
rect 26004 603676 26604 603678
rect 62004 603676 62604 603678
rect 98004 603676 98604 603678
rect 134004 603676 134604 603678
rect 170004 603676 170604 603678
rect 206004 603676 206604 603678
rect 242004 603676 242604 603678
rect 278004 603676 278604 603678
rect 314004 603676 314604 603678
rect 350004 603676 350604 603678
rect 386004 603676 386604 603678
rect 422004 603676 422604 603678
rect 458004 603676 458604 603678
rect 494004 603676 494604 603678
rect 530004 603676 530604 603678
rect 566004 603676 566604 603678
rect 589920 603676 590520 603678
rect -6596 603654 590520 603676
rect -6596 603418 -6414 603654
rect -6178 603418 26186 603654
rect 26422 603418 62186 603654
rect 62422 603418 98186 603654
rect 98422 603418 134186 603654
rect 134422 603418 170186 603654
rect 170422 603418 206186 603654
rect 206422 603418 242186 603654
rect 242422 603418 278186 603654
rect 278422 603418 314186 603654
rect 314422 603418 350186 603654
rect 350422 603418 386186 603654
rect 386422 603418 422186 603654
rect 422422 603418 458186 603654
rect 458422 603418 494186 603654
rect 494422 603418 530186 603654
rect 530422 603418 566186 603654
rect 566422 603418 590102 603654
rect 590338 603418 590520 603654
rect -6596 603334 590520 603418
rect -6596 603098 -6414 603334
rect -6178 603098 26186 603334
rect 26422 603098 62186 603334
rect 62422 603098 98186 603334
rect 98422 603098 134186 603334
rect 134422 603098 170186 603334
rect 170422 603098 206186 603334
rect 206422 603098 242186 603334
rect 242422 603098 278186 603334
rect 278422 603098 314186 603334
rect 314422 603098 350186 603334
rect 350422 603098 386186 603334
rect 386422 603098 422186 603334
rect 422422 603098 458186 603334
rect 458422 603098 494186 603334
rect 494422 603098 530186 603334
rect 530422 603098 566186 603334
rect 566422 603098 590102 603334
rect 590338 603098 590520 603334
rect -6596 603076 590520 603098
rect -6596 603074 -5996 603076
rect 26004 603074 26604 603076
rect 62004 603074 62604 603076
rect 98004 603074 98604 603076
rect 134004 603074 134604 603076
rect 170004 603074 170604 603076
rect 206004 603074 206604 603076
rect 242004 603074 242604 603076
rect 278004 603074 278604 603076
rect 314004 603074 314604 603076
rect 350004 603074 350604 603076
rect 386004 603074 386604 603076
rect 422004 603074 422604 603076
rect 458004 603074 458604 603076
rect 494004 603074 494604 603076
rect 530004 603074 530604 603076
rect 566004 603074 566604 603076
rect 589920 603074 590520 603076
rect -4756 600076 -4156 600078
rect 22404 600076 23004 600078
rect 58404 600076 59004 600078
rect 94404 600076 95004 600078
rect 130404 600076 131004 600078
rect 166404 600076 167004 600078
rect 202404 600076 203004 600078
rect 238404 600076 239004 600078
rect 274404 600076 275004 600078
rect 310404 600076 311004 600078
rect 346404 600076 347004 600078
rect 382404 600076 383004 600078
rect 418404 600076 419004 600078
rect 454404 600076 455004 600078
rect 490404 600076 491004 600078
rect 526404 600076 527004 600078
rect 562404 600076 563004 600078
rect 588080 600076 588680 600078
rect -4756 600054 588680 600076
rect -4756 599818 -4574 600054
rect -4338 599818 22586 600054
rect 22822 599818 58586 600054
rect 58822 599818 94586 600054
rect 94822 599818 130586 600054
rect 130822 599818 166586 600054
rect 166822 599818 202586 600054
rect 202822 599818 238586 600054
rect 238822 599818 274586 600054
rect 274822 599818 310586 600054
rect 310822 599818 346586 600054
rect 346822 599818 382586 600054
rect 382822 599818 418586 600054
rect 418822 599818 454586 600054
rect 454822 599818 490586 600054
rect 490822 599818 526586 600054
rect 526822 599818 562586 600054
rect 562822 599818 588262 600054
rect 588498 599818 588680 600054
rect -4756 599734 588680 599818
rect -4756 599498 -4574 599734
rect -4338 599498 22586 599734
rect 22822 599498 58586 599734
rect 58822 599498 94586 599734
rect 94822 599498 130586 599734
rect 130822 599498 166586 599734
rect 166822 599498 202586 599734
rect 202822 599498 238586 599734
rect 238822 599498 274586 599734
rect 274822 599498 310586 599734
rect 310822 599498 346586 599734
rect 346822 599498 382586 599734
rect 382822 599498 418586 599734
rect 418822 599498 454586 599734
rect 454822 599498 490586 599734
rect 490822 599498 526586 599734
rect 526822 599498 562586 599734
rect 562822 599498 588262 599734
rect 588498 599498 588680 599734
rect -4756 599476 588680 599498
rect -4756 599474 -4156 599476
rect 22404 599474 23004 599476
rect 58404 599474 59004 599476
rect 94404 599474 95004 599476
rect 130404 599474 131004 599476
rect 166404 599474 167004 599476
rect 202404 599474 203004 599476
rect 238404 599474 239004 599476
rect 274404 599474 275004 599476
rect 310404 599474 311004 599476
rect 346404 599474 347004 599476
rect 382404 599474 383004 599476
rect 418404 599474 419004 599476
rect 454404 599474 455004 599476
rect 490404 599474 491004 599476
rect 526404 599474 527004 599476
rect 562404 599474 563004 599476
rect 588080 599474 588680 599476
rect -2916 596476 -2316 596478
rect 18804 596476 19404 596478
rect 54804 596476 55404 596478
rect 90804 596476 91404 596478
rect 126804 596476 127404 596478
rect 162804 596476 163404 596478
rect 198804 596476 199404 596478
rect 234804 596476 235404 596478
rect 270804 596476 271404 596478
rect 306804 596476 307404 596478
rect 342804 596476 343404 596478
rect 378804 596476 379404 596478
rect 414804 596476 415404 596478
rect 450804 596476 451404 596478
rect 486804 596476 487404 596478
rect 522804 596476 523404 596478
rect 558804 596476 559404 596478
rect 586240 596476 586840 596478
rect -2916 596454 586840 596476
rect -2916 596218 -2734 596454
rect -2498 596218 18986 596454
rect 19222 596218 54986 596454
rect 55222 596218 90986 596454
rect 91222 596218 126986 596454
rect 127222 596218 162986 596454
rect 163222 596218 198986 596454
rect 199222 596218 234986 596454
rect 235222 596218 270986 596454
rect 271222 596218 306986 596454
rect 307222 596218 342986 596454
rect 343222 596218 378986 596454
rect 379222 596218 414986 596454
rect 415222 596218 450986 596454
rect 451222 596218 486986 596454
rect 487222 596218 522986 596454
rect 523222 596218 558986 596454
rect 559222 596218 586422 596454
rect 586658 596218 586840 596454
rect -2916 596134 586840 596218
rect -2916 595898 -2734 596134
rect -2498 595898 18986 596134
rect 19222 595898 54986 596134
rect 55222 595898 90986 596134
rect 91222 595898 126986 596134
rect 127222 595898 162986 596134
rect 163222 595898 198986 596134
rect 199222 595898 234986 596134
rect 235222 595898 270986 596134
rect 271222 595898 306986 596134
rect 307222 595898 342986 596134
rect 343222 595898 378986 596134
rect 379222 595898 414986 596134
rect 415222 595898 450986 596134
rect 451222 595898 486986 596134
rect 487222 595898 522986 596134
rect 523222 595898 558986 596134
rect 559222 595898 586422 596134
rect 586658 595898 586840 596134
rect -2916 595876 586840 595898
rect -2916 595874 -2316 595876
rect 18804 595874 19404 595876
rect 54804 595874 55404 595876
rect 90804 595874 91404 595876
rect 126804 595874 127404 595876
rect 162804 595874 163404 595876
rect 198804 595874 199404 595876
rect 234804 595874 235404 595876
rect 270804 595874 271404 595876
rect 306804 595874 307404 595876
rect 342804 595874 343404 595876
rect 378804 595874 379404 595876
rect 414804 595874 415404 595876
rect 450804 595874 451404 595876
rect 486804 595874 487404 595876
rect 522804 595874 523404 595876
rect 558804 595874 559404 595876
rect 586240 595874 586840 595876
rect -7516 589276 -6916 589278
rect 11604 589276 12204 589278
rect 47604 589276 48204 589278
rect 83604 589276 84204 589278
rect 119604 589276 120204 589278
rect 155604 589276 156204 589278
rect 191604 589276 192204 589278
rect 227604 589276 228204 589278
rect 263604 589276 264204 589278
rect 299604 589276 300204 589278
rect 335604 589276 336204 589278
rect 371604 589276 372204 589278
rect 407604 589276 408204 589278
rect 443604 589276 444204 589278
rect 479604 589276 480204 589278
rect 515604 589276 516204 589278
rect 551604 589276 552204 589278
rect 590840 589276 591440 589278
rect -8436 589254 592360 589276
rect -8436 589018 -7334 589254
rect -7098 589018 11786 589254
rect 12022 589018 47786 589254
rect 48022 589018 83786 589254
rect 84022 589018 119786 589254
rect 120022 589018 155786 589254
rect 156022 589018 191786 589254
rect 192022 589018 227786 589254
rect 228022 589018 263786 589254
rect 264022 589018 299786 589254
rect 300022 589018 335786 589254
rect 336022 589018 371786 589254
rect 372022 589018 407786 589254
rect 408022 589018 443786 589254
rect 444022 589018 479786 589254
rect 480022 589018 515786 589254
rect 516022 589018 551786 589254
rect 552022 589018 591022 589254
rect 591258 589018 592360 589254
rect -8436 588934 592360 589018
rect -8436 588698 -7334 588934
rect -7098 588698 11786 588934
rect 12022 588698 47786 588934
rect 48022 588698 83786 588934
rect 84022 588698 119786 588934
rect 120022 588698 155786 588934
rect 156022 588698 191786 588934
rect 192022 588698 227786 588934
rect 228022 588698 263786 588934
rect 264022 588698 299786 588934
rect 300022 588698 335786 588934
rect 336022 588698 371786 588934
rect 372022 588698 407786 588934
rect 408022 588698 443786 588934
rect 444022 588698 479786 588934
rect 480022 588698 515786 588934
rect 516022 588698 551786 588934
rect 552022 588698 591022 588934
rect 591258 588698 592360 588934
rect -8436 588676 592360 588698
rect -7516 588674 -6916 588676
rect 11604 588674 12204 588676
rect 47604 588674 48204 588676
rect 83604 588674 84204 588676
rect 119604 588674 120204 588676
rect 155604 588674 156204 588676
rect 191604 588674 192204 588676
rect 227604 588674 228204 588676
rect 263604 588674 264204 588676
rect 299604 588674 300204 588676
rect 335604 588674 336204 588676
rect 371604 588674 372204 588676
rect 407604 588674 408204 588676
rect 443604 588674 444204 588676
rect 479604 588674 480204 588676
rect 515604 588674 516204 588676
rect 551604 588674 552204 588676
rect 590840 588674 591440 588676
rect -5676 585676 -5076 585678
rect 8004 585676 8604 585678
rect 44004 585676 44604 585678
rect 80004 585676 80604 585678
rect 116004 585676 116604 585678
rect 152004 585676 152604 585678
rect 188004 585676 188604 585678
rect 224004 585676 224604 585678
rect 260004 585676 260604 585678
rect 296004 585676 296604 585678
rect 332004 585676 332604 585678
rect 368004 585676 368604 585678
rect 404004 585676 404604 585678
rect 440004 585676 440604 585678
rect 476004 585676 476604 585678
rect 512004 585676 512604 585678
rect 548004 585676 548604 585678
rect 589000 585676 589600 585678
rect -6596 585654 590520 585676
rect -6596 585418 -5494 585654
rect -5258 585418 8186 585654
rect 8422 585418 44186 585654
rect 44422 585418 80186 585654
rect 80422 585418 116186 585654
rect 116422 585418 152186 585654
rect 152422 585418 188186 585654
rect 188422 585418 224186 585654
rect 224422 585418 260186 585654
rect 260422 585418 296186 585654
rect 296422 585418 332186 585654
rect 332422 585418 368186 585654
rect 368422 585418 404186 585654
rect 404422 585418 440186 585654
rect 440422 585418 476186 585654
rect 476422 585418 512186 585654
rect 512422 585418 548186 585654
rect 548422 585418 589182 585654
rect 589418 585418 590520 585654
rect -6596 585334 590520 585418
rect -6596 585098 -5494 585334
rect -5258 585098 8186 585334
rect 8422 585098 44186 585334
rect 44422 585098 80186 585334
rect 80422 585098 116186 585334
rect 116422 585098 152186 585334
rect 152422 585098 188186 585334
rect 188422 585098 224186 585334
rect 224422 585098 260186 585334
rect 260422 585098 296186 585334
rect 296422 585098 332186 585334
rect 332422 585098 368186 585334
rect 368422 585098 404186 585334
rect 404422 585098 440186 585334
rect 440422 585098 476186 585334
rect 476422 585098 512186 585334
rect 512422 585098 548186 585334
rect 548422 585098 589182 585334
rect 589418 585098 590520 585334
rect -6596 585076 590520 585098
rect -5676 585074 -5076 585076
rect 8004 585074 8604 585076
rect 44004 585074 44604 585076
rect 80004 585074 80604 585076
rect 116004 585074 116604 585076
rect 152004 585074 152604 585076
rect 188004 585074 188604 585076
rect 224004 585074 224604 585076
rect 260004 585074 260604 585076
rect 296004 585074 296604 585076
rect 332004 585074 332604 585076
rect 368004 585074 368604 585076
rect 404004 585074 404604 585076
rect 440004 585074 440604 585076
rect 476004 585074 476604 585076
rect 512004 585074 512604 585076
rect 548004 585074 548604 585076
rect 589000 585074 589600 585076
rect -3836 582076 -3236 582078
rect 4404 582076 5004 582078
rect 40404 582076 41004 582078
rect 76404 582076 77004 582078
rect 112404 582076 113004 582078
rect 148404 582076 149004 582078
rect 184404 582076 185004 582078
rect 220404 582076 221004 582078
rect 256404 582076 257004 582078
rect 292404 582076 293004 582078
rect 328404 582076 329004 582078
rect 364404 582076 365004 582078
rect 400404 582076 401004 582078
rect 436404 582076 437004 582078
rect 472404 582076 473004 582078
rect 508404 582076 509004 582078
rect 544404 582076 545004 582078
rect 580404 582076 581004 582078
rect 587160 582076 587760 582078
rect -4756 582054 588680 582076
rect -4756 581818 -3654 582054
rect -3418 581818 4586 582054
rect 4822 581818 40586 582054
rect 40822 581818 76586 582054
rect 76822 581818 112586 582054
rect 112822 581818 148586 582054
rect 148822 581818 184586 582054
rect 184822 581818 220586 582054
rect 220822 581818 256586 582054
rect 256822 581818 292586 582054
rect 292822 581818 328586 582054
rect 328822 581818 364586 582054
rect 364822 581818 400586 582054
rect 400822 581818 436586 582054
rect 436822 581818 472586 582054
rect 472822 581818 508586 582054
rect 508822 581818 544586 582054
rect 544822 581818 580586 582054
rect 580822 581818 587342 582054
rect 587578 581818 588680 582054
rect -4756 581734 588680 581818
rect -4756 581498 -3654 581734
rect -3418 581498 4586 581734
rect 4822 581498 40586 581734
rect 40822 581498 76586 581734
rect 76822 581498 112586 581734
rect 112822 581498 148586 581734
rect 148822 581498 184586 581734
rect 184822 581498 220586 581734
rect 220822 581498 256586 581734
rect 256822 581498 292586 581734
rect 292822 581498 328586 581734
rect 328822 581498 364586 581734
rect 364822 581498 400586 581734
rect 400822 581498 436586 581734
rect 436822 581498 472586 581734
rect 472822 581498 508586 581734
rect 508822 581498 544586 581734
rect 544822 581498 580586 581734
rect 580822 581498 587342 581734
rect 587578 581498 588680 581734
rect -4756 581476 588680 581498
rect -3836 581474 -3236 581476
rect 4404 581474 5004 581476
rect 40404 581474 41004 581476
rect 76404 581474 77004 581476
rect 112404 581474 113004 581476
rect 148404 581474 149004 581476
rect 184404 581474 185004 581476
rect 220404 581474 221004 581476
rect 256404 581474 257004 581476
rect 292404 581474 293004 581476
rect 328404 581474 329004 581476
rect 364404 581474 365004 581476
rect 400404 581474 401004 581476
rect 436404 581474 437004 581476
rect 472404 581474 473004 581476
rect 508404 581474 509004 581476
rect 544404 581474 545004 581476
rect 580404 581474 581004 581476
rect 587160 581474 587760 581476
rect -1996 578476 -1396 578478
rect 804 578476 1404 578478
rect 36804 578476 37404 578478
rect 72804 578476 73404 578478
rect 108804 578476 109404 578478
rect 144804 578476 145404 578478
rect 180804 578476 181404 578478
rect 216804 578476 217404 578478
rect 252804 578476 253404 578478
rect 288804 578476 289404 578478
rect 324804 578476 325404 578478
rect 360804 578476 361404 578478
rect 396804 578476 397404 578478
rect 432804 578476 433404 578478
rect 468804 578476 469404 578478
rect 504804 578476 505404 578478
rect 540804 578476 541404 578478
rect 576804 578476 577404 578478
rect 585320 578476 585920 578478
rect -2916 578454 586840 578476
rect -2916 578218 -1814 578454
rect -1578 578218 986 578454
rect 1222 578218 36986 578454
rect 37222 578218 72986 578454
rect 73222 578218 108986 578454
rect 109222 578218 144986 578454
rect 145222 578218 180986 578454
rect 181222 578218 216986 578454
rect 217222 578218 252986 578454
rect 253222 578218 288986 578454
rect 289222 578218 324986 578454
rect 325222 578218 360986 578454
rect 361222 578218 396986 578454
rect 397222 578218 432986 578454
rect 433222 578218 468986 578454
rect 469222 578218 504986 578454
rect 505222 578218 540986 578454
rect 541222 578218 576986 578454
rect 577222 578218 585502 578454
rect 585738 578218 586840 578454
rect -2916 578134 586840 578218
rect -2916 577898 -1814 578134
rect -1578 577898 986 578134
rect 1222 577898 36986 578134
rect 37222 577898 72986 578134
rect 73222 577898 108986 578134
rect 109222 577898 144986 578134
rect 145222 577898 180986 578134
rect 181222 577898 216986 578134
rect 217222 577898 252986 578134
rect 253222 577898 288986 578134
rect 289222 577898 324986 578134
rect 325222 577898 360986 578134
rect 361222 577898 396986 578134
rect 397222 577898 432986 578134
rect 433222 577898 468986 578134
rect 469222 577898 504986 578134
rect 505222 577898 540986 578134
rect 541222 577898 576986 578134
rect 577222 577898 585502 578134
rect 585738 577898 586840 578134
rect -2916 577876 586840 577898
rect -1996 577874 -1396 577876
rect 804 577874 1404 577876
rect 36804 577874 37404 577876
rect 72804 577874 73404 577876
rect 108804 577874 109404 577876
rect 144804 577874 145404 577876
rect 180804 577874 181404 577876
rect 216804 577874 217404 577876
rect 252804 577874 253404 577876
rect 288804 577874 289404 577876
rect 324804 577874 325404 577876
rect 360804 577874 361404 577876
rect 396804 577874 397404 577876
rect 432804 577874 433404 577876
rect 468804 577874 469404 577876
rect 504804 577874 505404 577876
rect 540804 577874 541404 577876
rect 576804 577874 577404 577876
rect 585320 577874 585920 577876
rect -8436 571276 -7836 571278
rect 29604 571276 30204 571278
rect 65604 571276 66204 571278
rect 101604 571276 102204 571278
rect 137604 571276 138204 571278
rect 173604 571276 174204 571278
rect 209604 571276 210204 571278
rect 245604 571276 246204 571278
rect 281604 571276 282204 571278
rect 317604 571276 318204 571278
rect 353604 571276 354204 571278
rect 389604 571276 390204 571278
rect 425604 571276 426204 571278
rect 461604 571276 462204 571278
rect 497604 571276 498204 571278
rect 533604 571276 534204 571278
rect 569604 571276 570204 571278
rect 591760 571276 592360 571278
rect -8436 571254 592360 571276
rect -8436 571018 -8254 571254
rect -8018 571018 29786 571254
rect 30022 571018 65786 571254
rect 66022 571018 101786 571254
rect 102022 571018 137786 571254
rect 138022 571018 173786 571254
rect 174022 571018 209786 571254
rect 210022 571018 245786 571254
rect 246022 571018 281786 571254
rect 282022 571018 317786 571254
rect 318022 571018 353786 571254
rect 354022 571018 389786 571254
rect 390022 571018 425786 571254
rect 426022 571018 461786 571254
rect 462022 571018 497786 571254
rect 498022 571018 533786 571254
rect 534022 571018 569786 571254
rect 570022 571018 591942 571254
rect 592178 571018 592360 571254
rect -8436 570934 592360 571018
rect -8436 570698 -8254 570934
rect -8018 570698 29786 570934
rect 30022 570698 65786 570934
rect 66022 570698 101786 570934
rect 102022 570698 137786 570934
rect 138022 570698 173786 570934
rect 174022 570698 209786 570934
rect 210022 570698 245786 570934
rect 246022 570698 281786 570934
rect 282022 570698 317786 570934
rect 318022 570698 353786 570934
rect 354022 570698 389786 570934
rect 390022 570698 425786 570934
rect 426022 570698 461786 570934
rect 462022 570698 497786 570934
rect 498022 570698 533786 570934
rect 534022 570698 569786 570934
rect 570022 570698 591942 570934
rect 592178 570698 592360 570934
rect -8436 570676 592360 570698
rect -8436 570674 -7836 570676
rect 29604 570674 30204 570676
rect 65604 570674 66204 570676
rect 101604 570674 102204 570676
rect 137604 570674 138204 570676
rect 173604 570674 174204 570676
rect 209604 570674 210204 570676
rect 245604 570674 246204 570676
rect 281604 570674 282204 570676
rect 317604 570674 318204 570676
rect 353604 570674 354204 570676
rect 389604 570674 390204 570676
rect 425604 570674 426204 570676
rect 461604 570674 462204 570676
rect 497604 570674 498204 570676
rect 533604 570674 534204 570676
rect 569604 570674 570204 570676
rect 591760 570674 592360 570676
rect -6596 567676 -5996 567678
rect 26004 567676 26604 567678
rect 62004 567676 62604 567678
rect 98004 567676 98604 567678
rect 134004 567676 134604 567678
rect 170004 567676 170604 567678
rect 206004 567676 206604 567678
rect 242004 567676 242604 567678
rect 278004 567676 278604 567678
rect 314004 567676 314604 567678
rect 350004 567676 350604 567678
rect 386004 567676 386604 567678
rect 422004 567676 422604 567678
rect 458004 567676 458604 567678
rect 494004 567676 494604 567678
rect 530004 567676 530604 567678
rect 566004 567676 566604 567678
rect 589920 567676 590520 567678
rect -6596 567654 590520 567676
rect -6596 567418 -6414 567654
rect -6178 567418 26186 567654
rect 26422 567418 62186 567654
rect 62422 567418 98186 567654
rect 98422 567418 134186 567654
rect 134422 567418 170186 567654
rect 170422 567418 206186 567654
rect 206422 567418 242186 567654
rect 242422 567418 278186 567654
rect 278422 567418 314186 567654
rect 314422 567418 350186 567654
rect 350422 567418 386186 567654
rect 386422 567418 422186 567654
rect 422422 567418 458186 567654
rect 458422 567418 494186 567654
rect 494422 567418 530186 567654
rect 530422 567418 566186 567654
rect 566422 567418 590102 567654
rect 590338 567418 590520 567654
rect -6596 567334 590520 567418
rect -6596 567098 -6414 567334
rect -6178 567098 26186 567334
rect 26422 567098 62186 567334
rect 62422 567098 98186 567334
rect 98422 567098 134186 567334
rect 134422 567098 170186 567334
rect 170422 567098 206186 567334
rect 206422 567098 242186 567334
rect 242422 567098 278186 567334
rect 278422 567098 314186 567334
rect 314422 567098 350186 567334
rect 350422 567098 386186 567334
rect 386422 567098 422186 567334
rect 422422 567098 458186 567334
rect 458422 567098 494186 567334
rect 494422 567098 530186 567334
rect 530422 567098 566186 567334
rect 566422 567098 590102 567334
rect 590338 567098 590520 567334
rect -6596 567076 590520 567098
rect -6596 567074 -5996 567076
rect 26004 567074 26604 567076
rect 62004 567074 62604 567076
rect 98004 567074 98604 567076
rect 134004 567074 134604 567076
rect 170004 567074 170604 567076
rect 206004 567074 206604 567076
rect 242004 567074 242604 567076
rect 278004 567074 278604 567076
rect 314004 567074 314604 567076
rect 350004 567074 350604 567076
rect 386004 567074 386604 567076
rect 422004 567074 422604 567076
rect 458004 567074 458604 567076
rect 494004 567074 494604 567076
rect 530004 567074 530604 567076
rect 566004 567074 566604 567076
rect 589920 567074 590520 567076
rect -4756 564076 -4156 564078
rect 22404 564076 23004 564078
rect 58404 564076 59004 564078
rect 94404 564076 95004 564078
rect 130404 564076 131004 564078
rect 166404 564076 167004 564078
rect 202404 564076 203004 564078
rect 238404 564076 239004 564078
rect 274404 564076 275004 564078
rect 310404 564076 311004 564078
rect 346404 564076 347004 564078
rect 382404 564076 383004 564078
rect 418404 564076 419004 564078
rect 454404 564076 455004 564078
rect 490404 564076 491004 564078
rect 526404 564076 527004 564078
rect 562404 564076 563004 564078
rect 588080 564076 588680 564078
rect -4756 564054 588680 564076
rect -4756 563818 -4574 564054
rect -4338 563818 22586 564054
rect 22822 563818 58586 564054
rect 58822 563818 94586 564054
rect 94822 563818 130586 564054
rect 130822 563818 166586 564054
rect 166822 563818 202586 564054
rect 202822 563818 238586 564054
rect 238822 563818 274586 564054
rect 274822 563818 310586 564054
rect 310822 563818 346586 564054
rect 346822 563818 382586 564054
rect 382822 563818 418586 564054
rect 418822 563818 454586 564054
rect 454822 563818 490586 564054
rect 490822 563818 526586 564054
rect 526822 563818 562586 564054
rect 562822 563818 588262 564054
rect 588498 563818 588680 564054
rect -4756 563734 588680 563818
rect -4756 563498 -4574 563734
rect -4338 563498 22586 563734
rect 22822 563498 58586 563734
rect 58822 563498 94586 563734
rect 94822 563498 130586 563734
rect 130822 563498 166586 563734
rect 166822 563498 202586 563734
rect 202822 563498 238586 563734
rect 238822 563498 274586 563734
rect 274822 563498 310586 563734
rect 310822 563498 346586 563734
rect 346822 563498 382586 563734
rect 382822 563498 418586 563734
rect 418822 563498 454586 563734
rect 454822 563498 490586 563734
rect 490822 563498 526586 563734
rect 526822 563498 562586 563734
rect 562822 563498 588262 563734
rect 588498 563498 588680 563734
rect -4756 563476 588680 563498
rect -4756 563474 -4156 563476
rect 22404 563474 23004 563476
rect 58404 563474 59004 563476
rect 94404 563474 95004 563476
rect 130404 563474 131004 563476
rect 166404 563474 167004 563476
rect 202404 563474 203004 563476
rect 238404 563474 239004 563476
rect 274404 563474 275004 563476
rect 310404 563474 311004 563476
rect 346404 563474 347004 563476
rect 382404 563474 383004 563476
rect 418404 563474 419004 563476
rect 454404 563474 455004 563476
rect 490404 563474 491004 563476
rect 526404 563474 527004 563476
rect 562404 563474 563004 563476
rect 588080 563474 588680 563476
rect -2916 560476 -2316 560478
rect 18804 560476 19404 560478
rect 54804 560476 55404 560478
rect 90804 560476 91404 560478
rect 126804 560476 127404 560478
rect 162804 560476 163404 560478
rect 198804 560476 199404 560478
rect 234804 560476 235404 560478
rect 270804 560476 271404 560478
rect 306804 560476 307404 560478
rect 342804 560476 343404 560478
rect 378804 560476 379404 560478
rect 414804 560476 415404 560478
rect 450804 560476 451404 560478
rect 486804 560476 487404 560478
rect 522804 560476 523404 560478
rect 558804 560476 559404 560478
rect 586240 560476 586840 560478
rect -2916 560454 586840 560476
rect -2916 560218 -2734 560454
rect -2498 560218 18986 560454
rect 19222 560218 54986 560454
rect 55222 560218 90986 560454
rect 91222 560218 126986 560454
rect 127222 560218 162986 560454
rect 163222 560218 198986 560454
rect 199222 560218 234986 560454
rect 235222 560218 270986 560454
rect 271222 560218 306986 560454
rect 307222 560218 342986 560454
rect 343222 560218 378986 560454
rect 379222 560218 414986 560454
rect 415222 560218 450986 560454
rect 451222 560218 486986 560454
rect 487222 560218 522986 560454
rect 523222 560218 558986 560454
rect 559222 560218 586422 560454
rect 586658 560218 586840 560454
rect -2916 560134 586840 560218
rect -2916 559898 -2734 560134
rect -2498 559898 18986 560134
rect 19222 559898 54986 560134
rect 55222 559898 90986 560134
rect 91222 559898 126986 560134
rect 127222 559898 162986 560134
rect 163222 559898 198986 560134
rect 199222 559898 234986 560134
rect 235222 559898 270986 560134
rect 271222 559898 306986 560134
rect 307222 559898 342986 560134
rect 343222 559898 378986 560134
rect 379222 559898 414986 560134
rect 415222 559898 450986 560134
rect 451222 559898 486986 560134
rect 487222 559898 522986 560134
rect 523222 559898 558986 560134
rect 559222 559898 586422 560134
rect 586658 559898 586840 560134
rect -2916 559876 586840 559898
rect -2916 559874 -2316 559876
rect 18804 559874 19404 559876
rect 54804 559874 55404 559876
rect 90804 559874 91404 559876
rect 126804 559874 127404 559876
rect 162804 559874 163404 559876
rect 198804 559874 199404 559876
rect 234804 559874 235404 559876
rect 270804 559874 271404 559876
rect 306804 559874 307404 559876
rect 342804 559874 343404 559876
rect 378804 559874 379404 559876
rect 414804 559874 415404 559876
rect 450804 559874 451404 559876
rect 486804 559874 487404 559876
rect 522804 559874 523404 559876
rect 558804 559874 559404 559876
rect 586240 559874 586840 559876
rect -7516 553276 -6916 553278
rect 11604 553276 12204 553278
rect 47604 553276 48204 553278
rect 83604 553276 84204 553278
rect 119604 553276 120204 553278
rect 155604 553276 156204 553278
rect 191604 553276 192204 553278
rect 227604 553276 228204 553278
rect 263604 553276 264204 553278
rect 299604 553276 300204 553278
rect 335604 553276 336204 553278
rect 371604 553276 372204 553278
rect 407604 553276 408204 553278
rect 443604 553276 444204 553278
rect 479604 553276 480204 553278
rect 515604 553276 516204 553278
rect 551604 553276 552204 553278
rect 590840 553276 591440 553278
rect -8436 553254 592360 553276
rect -8436 553018 -7334 553254
rect -7098 553018 11786 553254
rect 12022 553018 47786 553254
rect 48022 553018 83786 553254
rect 84022 553018 119786 553254
rect 120022 553018 155786 553254
rect 156022 553018 191786 553254
rect 192022 553018 227786 553254
rect 228022 553018 263786 553254
rect 264022 553018 299786 553254
rect 300022 553018 335786 553254
rect 336022 553018 371786 553254
rect 372022 553018 407786 553254
rect 408022 553018 443786 553254
rect 444022 553018 479786 553254
rect 480022 553018 515786 553254
rect 516022 553018 551786 553254
rect 552022 553018 591022 553254
rect 591258 553018 592360 553254
rect -8436 552934 592360 553018
rect -8436 552698 -7334 552934
rect -7098 552698 11786 552934
rect 12022 552698 47786 552934
rect 48022 552698 83786 552934
rect 84022 552698 119786 552934
rect 120022 552698 155786 552934
rect 156022 552698 191786 552934
rect 192022 552698 227786 552934
rect 228022 552698 263786 552934
rect 264022 552698 299786 552934
rect 300022 552698 335786 552934
rect 336022 552698 371786 552934
rect 372022 552698 407786 552934
rect 408022 552698 443786 552934
rect 444022 552698 479786 552934
rect 480022 552698 515786 552934
rect 516022 552698 551786 552934
rect 552022 552698 591022 552934
rect 591258 552698 592360 552934
rect -8436 552676 592360 552698
rect -7516 552674 -6916 552676
rect 11604 552674 12204 552676
rect 47604 552674 48204 552676
rect 83604 552674 84204 552676
rect 119604 552674 120204 552676
rect 155604 552674 156204 552676
rect 191604 552674 192204 552676
rect 227604 552674 228204 552676
rect 263604 552674 264204 552676
rect 299604 552674 300204 552676
rect 335604 552674 336204 552676
rect 371604 552674 372204 552676
rect 407604 552674 408204 552676
rect 443604 552674 444204 552676
rect 479604 552674 480204 552676
rect 515604 552674 516204 552676
rect 551604 552674 552204 552676
rect 590840 552674 591440 552676
rect -5676 549676 -5076 549678
rect 8004 549676 8604 549678
rect 44004 549676 44604 549678
rect 80004 549676 80604 549678
rect 116004 549676 116604 549678
rect 152004 549676 152604 549678
rect 188004 549676 188604 549678
rect 224004 549676 224604 549678
rect 260004 549676 260604 549678
rect 296004 549676 296604 549678
rect 332004 549676 332604 549678
rect 368004 549676 368604 549678
rect 404004 549676 404604 549678
rect 440004 549676 440604 549678
rect 476004 549676 476604 549678
rect 512004 549676 512604 549678
rect 548004 549676 548604 549678
rect 589000 549676 589600 549678
rect -6596 549654 590520 549676
rect -6596 549418 -5494 549654
rect -5258 549418 8186 549654
rect 8422 549418 44186 549654
rect 44422 549418 80186 549654
rect 80422 549418 116186 549654
rect 116422 549418 152186 549654
rect 152422 549418 188186 549654
rect 188422 549418 224186 549654
rect 224422 549418 260186 549654
rect 260422 549418 296186 549654
rect 296422 549418 332186 549654
rect 332422 549418 368186 549654
rect 368422 549418 404186 549654
rect 404422 549418 440186 549654
rect 440422 549418 476186 549654
rect 476422 549418 512186 549654
rect 512422 549418 548186 549654
rect 548422 549418 589182 549654
rect 589418 549418 590520 549654
rect -6596 549334 590520 549418
rect -6596 549098 -5494 549334
rect -5258 549098 8186 549334
rect 8422 549098 44186 549334
rect 44422 549098 80186 549334
rect 80422 549098 116186 549334
rect 116422 549098 152186 549334
rect 152422 549098 188186 549334
rect 188422 549098 224186 549334
rect 224422 549098 260186 549334
rect 260422 549098 296186 549334
rect 296422 549098 332186 549334
rect 332422 549098 368186 549334
rect 368422 549098 404186 549334
rect 404422 549098 440186 549334
rect 440422 549098 476186 549334
rect 476422 549098 512186 549334
rect 512422 549098 548186 549334
rect 548422 549098 589182 549334
rect 589418 549098 590520 549334
rect -6596 549076 590520 549098
rect -5676 549074 -5076 549076
rect 8004 549074 8604 549076
rect 44004 549074 44604 549076
rect 80004 549074 80604 549076
rect 116004 549074 116604 549076
rect 152004 549074 152604 549076
rect 188004 549074 188604 549076
rect 224004 549074 224604 549076
rect 260004 549074 260604 549076
rect 296004 549074 296604 549076
rect 332004 549074 332604 549076
rect 368004 549074 368604 549076
rect 404004 549074 404604 549076
rect 440004 549074 440604 549076
rect 476004 549074 476604 549076
rect 512004 549074 512604 549076
rect 548004 549074 548604 549076
rect 589000 549074 589600 549076
rect -3836 546076 -3236 546078
rect 4404 546076 5004 546078
rect 40404 546076 41004 546078
rect 76404 546076 77004 546078
rect 112404 546076 113004 546078
rect 148404 546076 149004 546078
rect 184404 546076 185004 546078
rect 220404 546076 221004 546078
rect 256404 546076 257004 546078
rect 292404 546076 293004 546078
rect 328404 546076 329004 546078
rect 364404 546076 365004 546078
rect 400404 546076 401004 546078
rect 436404 546076 437004 546078
rect 472404 546076 473004 546078
rect 508404 546076 509004 546078
rect 544404 546076 545004 546078
rect 580404 546076 581004 546078
rect 587160 546076 587760 546078
rect -4756 546054 588680 546076
rect -4756 545818 -3654 546054
rect -3418 545818 4586 546054
rect 4822 545818 40586 546054
rect 40822 545818 76586 546054
rect 76822 545818 112586 546054
rect 112822 545818 148586 546054
rect 148822 545818 184586 546054
rect 184822 545818 220586 546054
rect 220822 545818 256586 546054
rect 256822 545818 292586 546054
rect 292822 545818 328586 546054
rect 328822 545818 364586 546054
rect 364822 545818 400586 546054
rect 400822 545818 436586 546054
rect 436822 545818 472586 546054
rect 472822 545818 508586 546054
rect 508822 545818 544586 546054
rect 544822 545818 580586 546054
rect 580822 545818 587342 546054
rect 587578 545818 588680 546054
rect -4756 545734 588680 545818
rect -4756 545498 -3654 545734
rect -3418 545498 4586 545734
rect 4822 545498 40586 545734
rect 40822 545498 76586 545734
rect 76822 545498 112586 545734
rect 112822 545498 148586 545734
rect 148822 545498 184586 545734
rect 184822 545498 220586 545734
rect 220822 545498 256586 545734
rect 256822 545498 292586 545734
rect 292822 545498 328586 545734
rect 328822 545498 364586 545734
rect 364822 545498 400586 545734
rect 400822 545498 436586 545734
rect 436822 545498 472586 545734
rect 472822 545498 508586 545734
rect 508822 545498 544586 545734
rect 544822 545498 580586 545734
rect 580822 545498 587342 545734
rect 587578 545498 588680 545734
rect -4756 545476 588680 545498
rect -3836 545474 -3236 545476
rect 4404 545474 5004 545476
rect 40404 545474 41004 545476
rect 76404 545474 77004 545476
rect 112404 545474 113004 545476
rect 148404 545474 149004 545476
rect 184404 545474 185004 545476
rect 220404 545474 221004 545476
rect 256404 545474 257004 545476
rect 292404 545474 293004 545476
rect 328404 545474 329004 545476
rect 364404 545474 365004 545476
rect 400404 545474 401004 545476
rect 436404 545474 437004 545476
rect 472404 545474 473004 545476
rect 508404 545474 509004 545476
rect 544404 545474 545004 545476
rect 580404 545474 581004 545476
rect 587160 545474 587760 545476
rect -1996 542476 -1396 542478
rect 804 542476 1404 542478
rect 36804 542476 37404 542478
rect 72804 542476 73404 542478
rect 108804 542476 109404 542478
rect 144804 542476 145404 542478
rect 180804 542476 181404 542478
rect 216804 542476 217404 542478
rect 252804 542476 253404 542478
rect 288804 542476 289404 542478
rect 324804 542476 325404 542478
rect 360804 542476 361404 542478
rect 396804 542476 397404 542478
rect 432804 542476 433404 542478
rect 468804 542476 469404 542478
rect 504804 542476 505404 542478
rect 540804 542476 541404 542478
rect 576804 542476 577404 542478
rect 585320 542476 585920 542478
rect -2916 542454 586840 542476
rect -2916 542218 -1814 542454
rect -1578 542218 986 542454
rect 1222 542218 36986 542454
rect 37222 542218 72986 542454
rect 73222 542218 108986 542454
rect 109222 542218 144986 542454
rect 145222 542218 180986 542454
rect 181222 542218 216986 542454
rect 217222 542218 252986 542454
rect 253222 542218 288986 542454
rect 289222 542218 324986 542454
rect 325222 542218 360986 542454
rect 361222 542218 396986 542454
rect 397222 542218 432986 542454
rect 433222 542218 468986 542454
rect 469222 542218 504986 542454
rect 505222 542218 540986 542454
rect 541222 542218 576986 542454
rect 577222 542218 585502 542454
rect 585738 542218 586840 542454
rect -2916 542134 586840 542218
rect -2916 541898 -1814 542134
rect -1578 541898 986 542134
rect 1222 541898 36986 542134
rect 37222 541898 72986 542134
rect 73222 541898 108986 542134
rect 109222 541898 144986 542134
rect 145222 541898 180986 542134
rect 181222 541898 216986 542134
rect 217222 541898 252986 542134
rect 253222 541898 288986 542134
rect 289222 541898 324986 542134
rect 325222 541898 360986 542134
rect 361222 541898 396986 542134
rect 397222 541898 432986 542134
rect 433222 541898 468986 542134
rect 469222 541898 504986 542134
rect 505222 541898 540986 542134
rect 541222 541898 576986 542134
rect 577222 541898 585502 542134
rect 585738 541898 586840 542134
rect -2916 541876 586840 541898
rect -1996 541874 -1396 541876
rect 804 541874 1404 541876
rect 36804 541874 37404 541876
rect 72804 541874 73404 541876
rect 108804 541874 109404 541876
rect 144804 541874 145404 541876
rect 180804 541874 181404 541876
rect 216804 541874 217404 541876
rect 252804 541874 253404 541876
rect 288804 541874 289404 541876
rect 324804 541874 325404 541876
rect 360804 541874 361404 541876
rect 396804 541874 397404 541876
rect 432804 541874 433404 541876
rect 468804 541874 469404 541876
rect 504804 541874 505404 541876
rect 540804 541874 541404 541876
rect 576804 541874 577404 541876
rect 585320 541874 585920 541876
rect -8436 535276 -7836 535278
rect 29604 535276 30204 535278
rect 65604 535276 66204 535278
rect 101604 535276 102204 535278
rect 137604 535276 138204 535278
rect 173604 535276 174204 535278
rect 209604 535276 210204 535278
rect 245604 535276 246204 535278
rect 281604 535276 282204 535278
rect 317604 535276 318204 535278
rect 353604 535276 354204 535278
rect 389604 535276 390204 535278
rect 425604 535276 426204 535278
rect 461604 535276 462204 535278
rect 497604 535276 498204 535278
rect 533604 535276 534204 535278
rect 569604 535276 570204 535278
rect 591760 535276 592360 535278
rect -8436 535254 592360 535276
rect -8436 535018 -8254 535254
rect -8018 535018 29786 535254
rect 30022 535018 65786 535254
rect 66022 535018 101786 535254
rect 102022 535018 137786 535254
rect 138022 535018 173786 535254
rect 174022 535018 209786 535254
rect 210022 535018 245786 535254
rect 246022 535018 281786 535254
rect 282022 535018 317786 535254
rect 318022 535018 353786 535254
rect 354022 535018 389786 535254
rect 390022 535018 425786 535254
rect 426022 535018 461786 535254
rect 462022 535018 497786 535254
rect 498022 535018 533786 535254
rect 534022 535018 569786 535254
rect 570022 535018 591942 535254
rect 592178 535018 592360 535254
rect -8436 534934 592360 535018
rect -8436 534698 -8254 534934
rect -8018 534698 29786 534934
rect 30022 534698 65786 534934
rect 66022 534698 101786 534934
rect 102022 534698 137786 534934
rect 138022 534698 173786 534934
rect 174022 534698 209786 534934
rect 210022 534698 245786 534934
rect 246022 534698 281786 534934
rect 282022 534698 317786 534934
rect 318022 534698 353786 534934
rect 354022 534698 389786 534934
rect 390022 534698 425786 534934
rect 426022 534698 461786 534934
rect 462022 534698 497786 534934
rect 498022 534698 533786 534934
rect 534022 534698 569786 534934
rect 570022 534698 591942 534934
rect 592178 534698 592360 534934
rect -8436 534676 592360 534698
rect -8436 534674 -7836 534676
rect 29604 534674 30204 534676
rect 65604 534674 66204 534676
rect 101604 534674 102204 534676
rect 137604 534674 138204 534676
rect 173604 534674 174204 534676
rect 209604 534674 210204 534676
rect 245604 534674 246204 534676
rect 281604 534674 282204 534676
rect 317604 534674 318204 534676
rect 353604 534674 354204 534676
rect 389604 534674 390204 534676
rect 425604 534674 426204 534676
rect 461604 534674 462204 534676
rect 497604 534674 498204 534676
rect 533604 534674 534204 534676
rect 569604 534674 570204 534676
rect 591760 534674 592360 534676
rect -6596 531676 -5996 531678
rect 26004 531676 26604 531678
rect 62004 531676 62604 531678
rect 98004 531676 98604 531678
rect 134004 531676 134604 531678
rect 170004 531676 170604 531678
rect 206004 531676 206604 531678
rect 242004 531676 242604 531678
rect 278004 531676 278604 531678
rect 314004 531676 314604 531678
rect 350004 531676 350604 531678
rect 386004 531676 386604 531678
rect 422004 531676 422604 531678
rect 458004 531676 458604 531678
rect 494004 531676 494604 531678
rect 530004 531676 530604 531678
rect 566004 531676 566604 531678
rect 589920 531676 590520 531678
rect -6596 531654 590520 531676
rect -6596 531418 -6414 531654
rect -6178 531418 26186 531654
rect 26422 531418 62186 531654
rect 62422 531418 98186 531654
rect 98422 531418 134186 531654
rect 134422 531418 170186 531654
rect 170422 531418 206186 531654
rect 206422 531418 242186 531654
rect 242422 531418 278186 531654
rect 278422 531418 314186 531654
rect 314422 531418 350186 531654
rect 350422 531418 386186 531654
rect 386422 531418 422186 531654
rect 422422 531418 458186 531654
rect 458422 531418 494186 531654
rect 494422 531418 530186 531654
rect 530422 531418 566186 531654
rect 566422 531418 590102 531654
rect 590338 531418 590520 531654
rect -6596 531334 590520 531418
rect -6596 531098 -6414 531334
rect -6178 531098 26186 531334
rect 26422 531098 62186 531334
rect 62422 531098 98186 531334
rect 98422 531098 134186 531334
rect 134422 531098 170186 531334
rect 170422 531098 206186 531334
rect 206422 531098 242186 531334
rect 242422 531098 278186 531334
rect 278422 531098 314186 531334
rect 314422 531098 350186 531334
rect 350422 531098 386186 531334
rect 386422 531098 422186 531334
rect 422422 531098 458186 531334
rect 458422 531098 494186 531334
rect 494422 531098 530186 531334
rect 530422 531098 566186 531334
rect 566422 531098 590102 531334
rect 590338 531098 590520 531334
rect -6596 531076 590520 531098
rect -6596 531074 -5996 531076
rect 26004 531074 26604 531076
rect 62004 531074 62604 531076
rect 98004 531074 98604 531076
rect 134004 531074 134604 531076
rect 170004 531074 170604 531076
rect 206004 531074 206604 531076
rect 242004 531074 242604 531076
rect 278004 531074 278604 531076
rect 314004 531074 314604 531076
rect 350004 531074 350604 531076
rect 386004 531074 386604 531076
rect 422004 531074 422604 531076
rect 458004 531074 458604 531076
rect 494004 531074 494604 531076
rect 530004 531074 530604 531076
rect 566004 531074 566604 531076
rect 589920 531074 590520 531076
rect -4756 528076 -4156 528078
rect 22404 528076 23004 528078
rect 58404 528076 59004 528078
rect 94404 528076 95004 528078
rect 130404 528076 131004 528078
rect 166404 528076 167004 528078
rect 202404 528076 203004 528078
rect 238404 528076 239004 528078
rect 274404 528076 275004 528078
rect 310404 528076 311004 528078
rect 346404 528076 347004 528078
rect 382404 528076 383004 528078
rect 418404 528076 419004 528078
rect 454404 528076 455004 528078
rect 490404 528076 491004 528078
rect 526404 528076 527004 528078
rect 562404 528076 563004 528078
rect 588080 528076 588680 528078
rect -4756 528054 588680 528076
rect -4756 527818 -4574 528054
rect -4338 527818 22586 528054
rect 22822 527818 58586 528054
rect 58822 527818 94586 528054
rect 94822 527818 130586 528054
rect 130822 527818 166586 528054
rect 166822 527818 202586 528054
rect 202822 527818 238586 528054
rect 238822 527818 274586 528054
rect 274822 527818 310586 528054
rect 310822 527818 346586 528054
rect 346822 527818 382586 528054
rect 382822 527818 418586 528054
rect 418822 527818 454586 528054
rect 454822 527818 490586 528054
rect 490822 527818 526586 528054
rect 526822 527818 562586 528054
rect 562822 527818 588262 528054
rect 588498 527818 588680 528054
rect -4756 527734 588680 527818
rect -4756 527498 -4574 527734
rect -4338 527498 22586 527734
rect 22822 527498 58586 527734
rect 58822 527498 94586 527734
rect 94822 527498 130586 527734
rect 130822 527498 166586 527734
rect 166822 527498 202586 527734
rect 202822 527498 238586 527734
rect 238822 527498 274586 527734
rect 274822 527498 310586 527734
rect 310822 527498 346586 527734
rect 346822 527498 382586 527734
rect 382822 527498 418586 527734
rect 418822 527498 454586 527734
rect 454822 527498 490586 527734
rect 490822 527498 526586 527734
rect 526822 527498 562586 527734
rect 562822 527498 588262 527734
rect 588498 527498 588680 527734
rect -4756 527476 588680 527498
rect -4756 527474 -4156 527476
rect 22404 527474 23004 527476
rect 58404 527474 59004 527476
rect 94404 527474 95004 527476
rect 130404 527474 131004 527476
rect 166404 527474 167004 527476
rect 202404 527474 203004 527476
rect 238404 527474 239004 527476
rect 274404 527474 275004 527476
rect 310404 527474 311004 527476
rect 346404 527474 347004 527476
rect 382404 527474 383004 527476
rect 418404 527474 419004 527476
rect 454404 527474 455004 527476
rect 490404 527474 491004 527476
rect 526404 527474 527004 527476
rect 562404 527474 563004 527476
rect 588080 527474 588680 527476
rect -2916 524476 -2316 524478
rect 18804 524476 19404 524478
rect 54804 524476 55404 524478
rect 90804 524476 91404 524478
rect 126804 524476 127404 524478
rect 162804 524476 163404 524478
rect 198804 524476 199404 524478
rect 234804 524476 235404 524478
rect 270804 524476 271404 524478
rect 306804 524476 307404 524478
rect 342804 524476 343404 524478
rect 378804 524476 379404 524478
rect 414804 524476 415404 524478
rect 450804 524476 451404 524478
rect 486804 524476 487404 524478
rect 522804 524476 523404 524478
rect 558804 524476 559404 524478
rect 586240 524476 586840 524478
rect -2916 524454 586840 524476
rect -2916 524218 -2734 524454
rect -2498 524218 18986 524454
rect 19222 524218 54986 524454
rect 55222 524218 90986 524454
rect 91222 524218 126986 524454
rect 127222 524218 162986 524454
rect 163222 524218 198986 524454
rect 199222 524218 234986 524454
rect 235222 524218 270986 524454
rect 271222 524218 306986 524454
rect 307222 524218 342986 524454
rect 343222 524218 378986 524454
rect 379222 524218 414986 524454
rect 415222 524218 450986 524454
rect 451222 524218 486986 524454
rect 487222 524218 522986 524454
rect 523222 524218 558986 524454
rect 559222 524218 586422 524454
rect 586658 524218 586840 524454
rect -2916 524134 586840 524218
rect -2916 523898 -2734 524134
rect -2498 523898 18986 524134
rect 19222 523898 54986 524134
rect 55222 523898 90986 524134
rect 91222 523898 126986 524134
rect 127222 523898 162986 524134
rect 163222 523898 198986 524134
rect 199222 523898 234986 524134
rect 235222 523898 270986 524134
rect 271222 523898 306986 524134
rect 307222 523898 342986 524134
rect 343222 523898 378986 524134
rect 379222 523898 414986 524134
rect 415222 523898 450986 524134
rect 451222 523898 486986 524134
rect 487222 523898 522986 524134
rect 523222 523898 558986 524134
rect 559222 523898 586422 524134
rect 586658 523898 586840 524134
rect -2916 523876 586840 523898
rect -2916 523874 -2316 523876
rect 18804 523874 19404 523876
rect 54804 523874 55404 523876
rect 90804 523874 91404 523876
rect 126804 523874 127404 523876
rect 162804 523874 163404 523876
rect 198804 523874 199404 523876
rect 234804 523874 235404 523876
rect 270804 523874 271404 523876
rect 306804 523874 307404 523876
rect 342804 523874 343404 523876
rect 378804 523874 379404 523876
rect 414804 523874 415404 523876
rect 450804 523874 451404 523876
rect 486804 523874 487404 523876
rect 522804 523874 523404 523876
rect 558804 523874 559404 523876
rect 586240 523874 586840 523876
rect 210244 517938 219396 517980
rect 210244 517702 210286 517938
rect 210522 517702 219118 517938
rect 219354 517702 219396 517938
rect 210244 517660 219396 517702
rect 234348 517938 243868 517980
rect 234348 517702 234390 517938
rect 234626 517702 243590 517938
rect 243826 517702 243868 517938
rect 234348 517660 243868 517702
rect 244652 517938 254356 517980
rect 244652 517702 244694 517938
rect 244930 517702 254078 517938
rect 254314 517702 254356 517938
rect 244652 517660 254356 517702
rect 264340 517938 273676 517980
rect 264340 517702 264382 517938
rect 264618 517702 273398 517938
rect 273634 517702 273676 517938
rect 264340 517660 273676 517702
rect 283292 517938 302932 517980
rect 283292 517702 283334 517938
rect 283570 517702 302654 517938
rect 302890 517702 302932 517938
rect 283292 517660 302932 517702
rect 335180 517938 336604 517980
rect 335180 517702 335222 517938
rect 335458 517702 336326 517938
rect 336562 517702 336604 517938
rect 335180 517660 336604 517702
rect -7516 517276 -6916 517278
rect 11604 517276 12204 517278
rect 47604 517276 48204 517278
rect 83604 517276 84204 517278
rect 119604 517276 120204 517278
rect 155604 517276 156204 517278
rect 191604 517276 192204 517278
rect 227604 517276 228204 517278
rect 263604 517276 264204 517278
rect 299604 517276 300204 517278
rect 335604 517276 336204 517278
rect 371604 517276 372204 517278
rect 407604 517276 408204 517278
rect 443604 517276 444204 517278
rect 479604 517276 480204 517278
rect 515604 517276 516204 517278
rect 551604 517276 552204 517278
rect 590840 517276 591440 517278
rect -8436 517254 592360 517276
rect -8436 517018 -7334 517254
rect -7098 517018 11786 517254
rect 12022 517018 47786 517254
rect 48022 517018 83786 517254
rect 84022 517018 119786 517254
rect 120022 517018 155786 517254
rect 156022 517018 191786 517254
rect 192022 517018 227786 517254
rect 228022 517018 263786 517254
rect 264022 517018 299786 517254
rect 300022 517018 335786 517254
rect 336022 517018 371786 517254
rect 372022 517018 407786 517254
rect 408022 517018 443786 517254
rect 444022 517018 479786 517254
rect 480022 517018 515786 517254
rect 516022 517018 551786 517254
rect 552022 517018 591022 517254
rect 591258 517018 592360 517254
rect -8436 516934 592360 517018
rect -8436 516698 -7334 516934
rect -7098 516698 11786 516934
rect 12022 516698 47786 516934
rect 48022 516698 83786 516934
rect 84022 516698 119786 516934
rect 120022 516698 155786 516934
rect 156022 516698 191786 516934
rect 192022 516698 227786 516934
rect 228022 516698 263786 516934
rect 264022 516698 299786 516934
rect 300022 516698 335786 516934
rect 336022 516698 371786 516934
rect 372022 516698 407786 516934
rect 408022 516698 443786 516934
rect 444022 516698 479786 516934
rect 480022 516698 515786 516934
rect 516022 516698 551786 516934
rect 552022 516698 591022 516934
rect 591258 516698 592360 516934
rect -8436 516676 592360 516698
rect -7516 516674 -6916 516676
rect 11604 516674 12204 516676
rect 47604 516674 48204 516676
rect 83604 516674 84204 516676
rect 119604 516674 120204 516676
rect 155604 516674 156204 516676
rect 191604 516674 192204 516676
rect 227604 516674 228204 516676
rect 263604 516674 264204 516676
rect 299604 516674 300204 516676
rect 335604 516674 336204 516676
rect 371604 516674 372204 516676
rect 407604 516674 408204 516676
rect 443604 516674 444204 516676
rect 479604 516674 480204 516676
rect 515604 516674 516204 516676
rect 551604 516674 552204 516676
rect 590840 516674 591440 516676
rect -5676 513676 -5076 513678
rect 8004 513676 8604 513678
rect 44004 513676 44604 513678
rect 80004 513676 80604 513678
rect 116004 513676 116604 513678
rect 152004 513676 152604 513678
rect 188004 513676 188604 513678
rect 224004 513676 224604 513678
rect 260004 513676 260604 513678
rect 296004 513676 296604 513678
rect 332004 513676 332604 513678
rect 368004 513676 368604 513678
rect 404004 513676 404604 513678
rect 440004 513676 440604 513678
rect 476004 513676 476604 513678
rect 512004 513676 512604 513678
rect 548004 513676 548604 513678
rect 589000 513676 589600 513678
rect -6596 513654 590520 513676
rect -6596 513418 -5494 513654
rect -5258 513418 8186 513654
rect 8422 513418 44186 513654
rect 44422 513418 80186 513654
rect 80422 513418 116186 513654
rect 116422 513418 152186 513654
rect 152422 513418 188186 513654
rect 188422 513418 224186 513654
rect 224422 513418 260186 513654
rect 260422 513418 296186 513654
rect 296422 513418 332186 513654
rect 332422 513418 368186 513654
rect 368422 513418 404186 513654
rect 404422 513418 440186 513654
rect 440422 513418 476186 513654
rect 476422 513418 512186 513654
rect 512422 513418 548186 513654
rect 548422 513418 589182 513654
rect 589418 513418 590520 513654
rect -6596 513334 590520 513418
rect -6596 513098 -5494 513334
rect -5258 513098 8186 513334
rect 8422 513098 44186 513334
rect 44422 513098 80186 513334
rect 80422 513098 116186 513334
rect 116422 513098 152186 513334
rect 152422 513098 188186 513334
rect 188422 513098 224186 513334
rect 224422 513098 260186 513334
rect 260422 513098 296186 513334
rect 296422 513098 332186 513334
rect 332422 513098 368186 513334
rect 368422 513098 404186 513334
rect 404422 513098 440186 513334
rect 440422 513098 476186 513334
rect 476422 513098 512186 513334
rect 512422 513098 548186 513334
rect 548422 513098 589182 513334
rect 589418 513098 590520 513334
rect -6596 513076 590520 513098
rect -5676 513074 -5076 513076
rect 8004 513074 8604 513076
rect 44004 513074 44604 513076
rect 80004 513074 80604 513076
rect 116004 513074 116604 513076
rect 152004 513074 152604 513076
rect 188004 513074 188604 513076
rect 224004 513074 224604 513076
rect 260004 513074 260604 513076
rect 296004 513074 296604 513076
rect 332004 513074 332604 513076
rect 368004 513074 368604 513076
rect 404004 513074 404604 513076
rect 440004 513074 440604 513076
rect 476004 513074 476604 513076
rect 512004 513074 512604 513076
rect 548004 513074 548604 513076
rect 589000 513074 589600 513076
rect -3836 510076 -3236 510078
rect 4404 510076 5004 510078
rect 40404 510076 41004 510078
rect 76404 510076 77004 510078
rect 112404 510076 113004 510078
rect 148404 510076 149004 510078
rect 184404 510076 185004 510078
rect 220404 510076 221004 510078
rect 256404 510076 257004 510078
rect 292404 510076 293004 510078
rect 328404 510076 329004 510078
rect 364404 510076 365004 510078
rect 400404 510076 401004 510078
rect 436404 510076 437004 510078
rect 472404 510076 473004 510078
rect 508404 510076 509004 510078
rect 544404 510076 545004 510078
rect 580404 510076 581004 510078
rect 587160 510076 587760 510078
rect -4756 510054 588680 510076
rect -4756 509818 -3654 510054
rect -3418 509818 4586 510054
rect 4822 509818 40586 510054
rect 40822 509818 76586 510054
rect 76822 509818 112586 510054
rect 112822 509818 148586 510054
rect 148822 509818 184586 510054
rect 184822 509818 220586 510054
rect 220822 509818 256586 510054
rect 256822 509818 292586 510054
rect 292822 509818 328586 510054
rect 328822 509818 364586 510054
rect 364822 509818 400586 510054
rect 400822 509818 436586 510054
rect 436822 509818 472586 510054
rect 472822 509818 508586 510054
rect 508822 509818 544586 510054
rect 544822 509818 580586 510054
rect 580822 509818 587342 510054
rect 587578 509818 588680 510054
rect -4756 509734 588680 509818
rect -4756 509498 -3654 509734
rect -3418 509498 4586 509734
rect 4822 509498 40586 509734
rect 40822 509498 76586 509734
rect 76822 509498 112586 509734
rect 112822 509498 148586 509734
rect 148822 509498 184586 509734
rect 184822 509498 220586 509734
rect 220822 509498 256586 509734
rect 256822 509498 292586 509734
rect 292822 509498 328586 509734
rect 328822 509498 364586 509734
rect 364822 509498 400586 509734
rect 400822 509498 436586 509734
rect 436822 509498 472586 509734
rect 472822 509498 508586 509734
rect 508822 509498 544586 509734
rect 544822 509498 580586 509734
rect 580822 509498 587342 509734
rect 587578 509498 588680 509734
rect -4756 509476 588680 509498
rect -3836 509474 -3236 509476
rect 4404 509474 5004 509476
rect 40404 509474 41004 509476
rect 76404 509474 77004 509476
rect 112404 509474 113004 509476
rect 148404 509474 149004 509476
rect 184404 509474 185004 509476
rect 220404 509474 221004 509476
rect 256404 509474 257004 509476
rect 292404 509474 293004 509476
rect 328404 509474 329004 509476
rect 364404 509474 365004 509476
rect 400404 509474 401004 509476
rect 436404 509474 437004 509476
rect 472404 509474 473004 509476
rect 508404 509474 509004 509476
rect 544404 509474 545004 509476
rect 580404 509474 581004 509476
rect 587160 509474 587760 509476
rect -1996 506476 -1396 506478
rect 804 506476 1404 506478
rect 36804 506476 37404 506478
rect 72804 506476 73404 506478
rect 108804 506476 109404 506478
rect 144804 506476 145404 506478
rect 180804 506476 181404 506478
rect 216804 506476 217404 506478
rect 252804 506476 253404 506478
rect 288804 506476 289404 506478
rect 324804 506476 325404 506478
rect 360804 506476 361404 506478
rect 396804 506476 397404 506478
rect 432804 506476 433404 506478
rect 468804 506476 469404 506478
rect 504804 506476 505404 506478
rect 540804 506476 541404 506478
rect 576804 506476 577404 506478
rect 585320 506476 585920 506478
rect -2916 506454 586840 506476
rect -2916 506218 -1814 506454
rect -1578 506218 986 506454
rect 1222 506218 36986 506454
rect 37222 506218 72986 506454
rect 73222 506218 108986 506454
rect 109222 506218 144986 506454
rect 145222 506218 180986 506454
rect 181222 506218 216986 506454
rect 217222 506218 252986 506454
rect 253222 506218 288986 506454
rect 289222 506218 324986 506454
rect 325222 506218 360986 506454
rect 361222 506218 396986 506454
rect 397222 506218 432986 506454
rect 433222 506218 468986 506454
rect 469222 506218 504986 506454
rect 505222 506218 540986 506454
rect 541222 506218 576986 506454
rect 577222 506218 585502 506454
rect 585738 506218 586840 506454
rect -2916 506134 586840 506218
rect -2916 505898 -1814 506134
rect -1578 505898 986 506134
rect 1222 505898 36986 506134
rect 37222 505898 72986 506134
rect 73222 505898 108986 506134
rect 109222 505898 144986 506134
rect 145222 505898 180986 506134
rect 181222 505898 216986 506134
rect 217222 505898 252986 506134
rect 253222 505898 288986 506134
rect 289222 505898 324986 506134
rect 325222 505898 360986 506134
rect 361222 505898 396986 506134
rect 397222 505898 432986 506134
rect 433222 505898 468986 506134
rect 469222 505898 504986 506134
rect 505222 505898 540986 506134
rect 541222 505898 576986 506134
rect 577222 505898 585502 506134
rect 585738 505898 586840 506134
rect -2916 505876 586840 505898
rect -1996 505874 -1396 505876
rect 804 505874 1404 505876
rect 36804 505874 37404 505876
rect 72804 505874 73404 505876
rect 108804 505874 109404 505876
rect 144804 505874 145404 505876
rect 180804 505874 181404 505876
rect 216804 505874 217404 505876
rect 252804 505874 253404 505876
rect 288804 505874 289404 505876
rect 324804 505874 325404 505876
rect 360804 505874 361404 505876
rect 396804 505874 397404 505876
rect 432804 505874 433404 505876
rect 468804 505874 469404 505876
rect 504804 505874 505404 505876
rect 540804 505874 541404 505876
rect 576804 505874 577404 505876
rect 585320 505874 585920 505876
rect -8436 499276 -7836 499278
rect 29604 499276 30204 499278
rect 65604 499276 66204 499278
rect 101604 499276 102204 499278
rect 137604 499276 138204 499278
rect 173604 499276 174204 499278
rect 209604 499276 210204 499278
rect 245604 499276 246204 499278
rect 281604 499276 282204 499278
rect 317604 499276 318204 499278
rect 353604 499276 354204 499278
rect 389604 499276 390204 499278
rect 425604 499276 426204 499278
rect 461604 499276 462204 499278
rect 497604 499276 498204 499278
rect 533604 499276 534204 499278
rect 569604 499276 570204 499278
rect 591760 499276 592360 499278
rect -8436 499254 592360 499276
rect -8436 499018 -8254 499254
rect -8018 499018 29786 499254
rect 30022 499018 65786 499254
rect 66022 499018 101786 499254
rect 102022 499018 137786 499254
rect 138022 499018 173786 499254
rect 174022 499018 209786 499254
rect 210022 499018 245786 499254
rect 246022 499018 281786 499254
rect 282022 499018 317786 499254
rect 318022 499018 353786 499254
rect 354022 499018 389786 499254
rect 390022 499018 425786 499254
rect 426022 499018 461786 499254
rect 462022 499018 497786 499254
rect 498022 499018 533786 499254
rect 534022 499018 569786 499254
rect 570022 499018 591942 499254
rect 592178 499018 592360 499254
rect -8436 498934 592360 499018
rect -8436 498698 -8254 498934
rect -8018 498698 29786 498934
rect 30022 498698 65786 498934
rect 66022 498698 101786 498934
rect 102022 498698 137786 498934
rect 138022 498698 173786 498934
rect 174022 498698 209786 498934
rect 210022 498698 245786 498934
rect 246022 498698 281786 498934
rect 282022 498698 317786 498934
rect 318022 498698 353786 498934
rect 354022 498698 389786 498934
rect 390022 498698 425786 498934
rect 426022 498698 461786 498934
rect 462022 498698 497786 498934
rect 498022 498698 533786 498934
rect 534022 498698 569786 498934
rect 570022 498698 591942 498934
rect 592178 498698 592360 498934
rect -8436 498676 592360 498698
rect -8436 498674 -7836 498676
rect 29604 498674 30204 498676
rect 65604 498674 66204 498676
rect 101604 498674 102204 498676
rect 137604 498674 138204 498676
rect 173604 498674 174204 498676
rect 209604 498674 210204 498676
rect 245604 498674 246204 498676
rect 281604 498674 282204 498676
rect 317604 498674 318204 498676
rect 353604 498674 354204 498676
rect 389604 498674 390204 498676
rect 425604 498674 426204 498676
rect 461604 498674 462204 498676
rect 497604 498674 498204 498676
rect 533604 498674 534204 498676
rect 569604 498674 570204 498676
rect 591760 498674 592360 498676
rect -6596 495676 -5996 495678
rect 26004 495676 26604 495678
rect 62004 495676 62604 495678
rect 98004 495676 98604 495678
rect 134004 495676 134604 495678
rect 170004 495676 170604 495678
rect 206004 495676 206604 495678
rect 242004 495676 242604 495678
rect 278004 495676 278604 495678
rect 314004 495676 314604 495678
rect 350004 495676 350604 495678
rect 386004 495676 386604 495678
rect 422004 495676 422604 495678
rect 458004 495676 458604 495678
rect 494004 495676 494604 495678
rect 530004 495676 530604 495678
rect 566004 495676 566604 495678
rect 589920 495676 590520 495678
rect -6596 495654 590520 495676
rect -6596 495418 -6414 495654
rect -6178 495418 26186 495654
rect 26422 495418 62186 495654
rect 62422 495418 98186 495654
rect 98422 495418 134186 495654
rect 134422 495418 170186 495654
rect 170422 495418 206186 495654
rect 206422 495418 242186 495654
rect 242422 495418 278186 495654
rect 278422 495418 314186 495654
rect 314422 495418 350186 495654
rect 350422 495418 386186 495654
rect 386422 495418 422186 495654
rect 422422 495418 458186 495654
rect 458422 495418 494186 495654
rect 494422 495418 530186 495654
rect 530422 495418 566186 495654
rect 566422 495418 590102 495654
rect 590338 495418 590520 495654
rect -6596 495334 590520 495418
rect -6596 495098 -6414 495334
rect -6178 495098 26186 495334
rect 26422 495098 62186 495334
rect 62422 495098 98186 495334
rect 98422 495098 134186 495334
rect 134422 495098 170186 495334
rect 170422 495098 206186 495334
rect 206422 495098 242186 495334
rect 242422 495098 278186 495334
rect 278422 495098 314186 495334
rect 314422 495098 350186 495334
rect 350422 495098 386186 495334
rect 386422 495098 422186 495334
rect 422422 495098 458186 495334
rect 458422 495098 494186 495334
rect 494422 495098 530186 495334
rect 530422 495098 566186 495334
rect 566422 495098 590102 495334
rect 590338 495098 590520 495334
rect -6596 495076 590520 495098
rect -6596 495074 -5996 495076
rect 26004 495074 26604 495076
rect 62004 495074 62604 495076
rect 98004 495074 98604 495076
rect 134004 495074 134604 495076
rect 170004 495074 170604 495076
rect 206004 495074 206604 495076
rect 242004 495074 242604 495076
rect 278004 495074 278604 495076
rect 314004 495074 314604 495076
rect 350004 495074 350604 495076
rect 386004 495074 386604 495076
rect 422004 495074 422604 495076
rect 458004 495074 458604 495076
rect 494004 495074 494604 495076
rect 530004 495074 530604 495076
rect 566004 495074 566604 495076
rect 589920 495074 590520 495076
rect -4756 492076 -4156 492078
rect 22404 492076 23004 492078
rect 58404 492076 59004 492078
rect 94404 492076 95004 492078
rect 130404 492076 131004 492078
rect 166404 492076 167004 492078
rect 202404 492076 203004 492078
rect 238404 492076 239004 492078
rect 274404 492076 275004 492078
rect 310404 492076 311004 492078
rect 346404 492076 347004 492078
rect 382404 492076 383004 492078
rect 418404 492076 419004 492078
rect 454404 492076 455004 492078
rect 490404 492076 491004 492078
rect 526404 492076 527004 492078
rect 562404 492076 563004 492078
rect 588080 492076 588680 492078
rect -4756 492054 588680 492076
rect -4756 491818 -4574 492054
rect -4338 491818 22586 492054
rect 22822 491818 58586 492054
rect 58822 491818 94586 492054
rect 94822 491818 130586 492054
rect 130822 491818 166586 492054
rect 166822 491818 202586 492054
rect 202822 491818 238586 492054
rect 238822 491818 274586 492054
rect 274822 491818 310586 492054
rect 310822 491818 346586 492054
rect 346822 491818 382586 492054
rect 382822 491818 418586 492054
rect 418822 491818 454586 492054
rect 454822 491818 490586 492054
rect 490822 491818 526586 492054
rect 526822 491818 562586 492054
rect 562822 491818 588262 492054
rect 588498 491818 588680 492054
rect -4756 491734 588680 491818
rect -4756 491498 -4574 491734
rect -4338 491498 22586 491734
rect 22822 491498 58586 491734
rect 58822 491498 94586 491734
rect 94822 491498 130586 491734
rect 130822 491498 166586 491734
rect 166822 491498 202586 491734
rect 202822 491498 238586 491734
rect 238822 491498 274586 491734
rect 274822 491498 310586 491734
rect 310822 491498 346586 491734
rect 346822 491498 382586 491734
rect 382822 491498 418586 491734
rect 418822 491498 454586 491734
rect 454822 491498 490586 491734
rect 490822 491498 526586 491734
rect 526822 491498 562586 491734
rect 562822 491498 588262 491734
rect 588498 491498 588680 491734
rect -4756 491476 588680 491498
rect -4756 491474 -4156 491476
rect 22404 491474 23004 491476
rect 58404 491474 59004 491476
rect 94404 491474 95004 491476
rect 130404 491474 131004 491476
rect 166404 491474 167004 491476
rect 202404 491474 203004 491476
rect 238404 491474 239004 491476
rect 274404 491474 275004 491476
rect 310404 491474 311004 491476
rect 346404 491474 347004 491476
rect 382404 491474 383004 491476
rect 418404 491474 419004 491476
rect 454404 491474 455004 491476
rect 490404 491474 491004 491476
rect 526404 491474 527004 491476
rect 562404 491474 563004 491476
rect 588080 491474 588680 491476
rect -2916 488476 -2316 488478
rect 18804 488476 19404 488478
rect 54804 488476 55404 488478
rect 90804 488476 91404 488478
rect 126804 488476 127404 488478
rect 162804 488476 163404 488478
rect 198804 488476 199404 488478
rect 234804 488476 235404 488478
rect 270804 488476 271404 488478
rect 306804 488476 307404 488478
rect 342804 488476 343404 488478
rect 378804 488476 379404 488478
rect 414804 488476 415404 488478
rect 450804 488476 451404 488478
rect 486804 488476 487404 488478
rect 522804 488476 523404 488478
rect 558804 488476 559404 488478
rect 586240 488476 586840 488478
rect -2916 488454 586840 488476
rect -2916 488218 -2734 488454
rect -2498 488218 18986 488454
rect 19222 488218 54986 488454
rect 55222 488218 90986 488454
rect 91222 488218 126986 488454
rect 127222 488218 162986 488454
rect 163222 488218 198986 488454
rect 199222 488218 234986 488454
rect 235222 488218 270986 488454
rect 271222 488218 306986 488454
rect 307222 488218 342986 488454
rect 343222 488218 378986 488454
rect 379222 488218 414986 488454
rect 415222 488218 450986 488454
rect 451222 488218 486986 488454
rect 487222 488218 522986 488454
rect 523222 488218 558986 488454
rect 559222 488218 586422 488454
rect 586658 488218 586840 488454
rect -2916 488134 586840 488218
rect -2916 487898 -2734 488134
rect -2498 487898 18986 488134
rect 19222 487898 54986 488134
rect 55222 487898 90986 488134
rect 91222 487898 126986 488134
rect 127222 487898 162986 488134
rect 163222 487898 198986 488134
rect 199222 487898 234986 488134
rect 235222 487898 270986 488134
rect 271222 487898 306986 488134
rect 307222 487898 342986 488134
rect 343222 487898 378986 488134
rect 379222 487898 414986 488134
rect 415222 487898 450986 488134
rect 451222 487898 486986 488134
rect 487222 487898 522986 488134
rect 523222 487898 558986 488134
rect 559222 487898 586422 488134
rect 586658 487898 586840 488134
rect -2916 487876 586840 487898
rect -2916 487874 -2316 487876
rect 18804 487874 19404 487876
rect 54804 487874 55404 487876
rect 90804 487874 91404 487876
rect 126804 487874 127404 487876
rect 162804 487874 163404 487876
rect 198804 487874 199404 487876
rect 234804 487874 235404 487876
rect 270804 487874 271404 487876
rect 306804 487874 307404 487876
rect 342804 487874 343404 487876
rect 378804 487874 379404 487876
rect 414804 487874 415404 487876
rect 450804 487874 451404 487876
rect 486804 487874 487404 487876
rect 522804 487874 523404 487876
rect 558804 487874 559404 487876
rect 586240 487874 586840 487876
rect -7516 481276 -6916 481278
rect 11604 481276 12204 481278
rect 47604 481276 48204 481278
rect 83604 481276 84204 481278
rect 119604 481276 120204 481278
rect 155604 481276 156204 481278
rect 191604 481276 192204 481278
rect 227604 481276 228204 481278
rect 263604 481276 264204 481278
rect 299604 481276 300204 481278
rect 335604 481276 336204 481278
rect 371604 481276 372204 481278
rect 407604 481276 408204 481278
rect 443604 481276 444204 481278
rect 479604 481276 480204 481278
rect 515604 481276 516204 481278
rect 551604 481276 552204 481278
rect 590840 481276 591440 481278
rect -8436 481254 592360 481276
rect -8436 481018 -7334 481254
rect -7098 481018 11786 481254
rect 12022 481018 47786 481254
rect 48022 481018 83786 481254
rect 84022 481018 119786 481254
rect 120022 481018 155786 481254
rect 156022 481018 191786 481254
rect 192022 481018 227786 481254
rect 228022 481018 263786 481254
rect 264022 481018 299786 481254
rect 300022 481018 335786 481254
rect 336022 481018 371786 481254
rect 372022 481018 407786 481254
rect 408022 481018 443786 481254
rect 444022 481018 479786 481254
rect 480022 481018 515786 481254
rect 516022 481018 551786 481254
rect 552022 481018 591022 481254
rect 591258 481018 592360 481254
rect -8436 480934 592360 481018
rect -8436 480698 -7334 480934
rect -7098 480698 11786 480934
rect 12022 480698 47786 480934
rect 48022 480698 83786 480934
rect 84022 480698 119786 480934
rect 120022 480698 155786 480934
rect 156022 480698 191786 480934
rect 192022 480698 227786 480934
rect 228022 480698 263786 480934
rect 264022 480698 299786 480934
rect 300022 480698 335786 480934
rect 336022 480698 371786 480934
rect 372022 480698 407786 480934
rect 408022 480698 443786 480934
rect 444022 480698 479786 480934
rect 480022 480698 515786 480934
rect 516022 480698 551786 480934
rect 552022 480698 591022 480934
rect 591258 480698 592360 480934
rect -8436 480676 592360 480698
rect -7516 480674 -6916 480676
rect 11604 480674 12204 480676
rect 47604 480674 48204 480676
rect 83604 480674 84204 480676
rect 119604 480674 120204 480676
rect 155604 480674 156204 480676
rect 191604 480674 192204 480676
rect 227604 480674 228204 480676
rect 263604 480674 264204 480676
rect 299604 480674 300204 480676
rect 335604 480674 336204 480676
rect 371604 480674 372204 480676
rect 407604 480674 408204 480676
rect 443604 480674 444204 480676
rect 479604 480674 480204 480676
rect 515604 480674 516204 480676
rect 551604 480674 552204 480676
rect 590840 480674 591440 480676
rect -5676 477676 -5076 477678
rect 8004 477676 8604 477678
rect 44004 477676 44604 477678
rect 80004 477676 80604 477678
rect 116004 477676 116604 477678
rect 152004 477676 152604 477678
rect 188004 477676 188604 477678
rect 224004 477676 224604 477678
rect 260004 477676 260604 477678
rect 296004 477676 296604 477678
rect 332004 477676 332604 477678
rect 368004 477676 368604 477678
rect 404004 477676 404604 477678
rect 440004 477676 440604 477678
rect 476004 477676 476604 477678
rect 512004 477676 512604 477678
rect 548004 477676 548604 477678
rect 589000 477676 589600 477678
rect -6596 477654 590520 477676
rect -6596 477418 -5494 477654
rect -5258 477418 8186 477654
rect 8422 477418 44186 477654
rect 44422 477418 80186 477654
rect 80422 477418 116186 477654
rect 116422 477418 152186 477654
rect 152422 477418 188186 477654
rect 188422 477418 224186 477654
rect 224422 477418 260186 477654
rect 260422 477418 296186 477654
rect 296422 477418 332186 477654
rect 332422 477418 368186 477654
rect 368422 477418 404186 477654
rect 404422 477418 440186 477654
rect 440422 477418 476186 477654
rect 476422 477418 512186 477654
rect 512422 477418 548186 477654
rect 548422 477418 589182 477654
rect 589418 477418 590520 477654
rect -6596 477334 590520 477418
rect -6596 477098 -5494 477334
rect -5258 477098 8186 477334
rect 8422 477098 44186 477334
rect 44422 477098 80186 477334
rect 80422 477098 116186 477334
rect 116422 477098 152186 477334
rect 152422 477098 188186 477334
rect 188422 477098 224186 477334
rect 224422 477098 260186 477334
rect 260422 477098 296186 477334
rect 296422 477098 332186 477334
rect 332422 477098 368186 477334
rect 368422 477098 404186 477334
rect 404422 477098 440186 477334
rect 440422 477098 476186 477334
rect 476422 477098 512186 477334
rect 512422 477098 548186 477334
rect 548422 477098 589182 477334
rect 589418 477098 590520 477334
rect -6596 477076 590520 477098
rect -5676 477074 -5076 477076
rect 8004 477074 8604 477076
rect 44004 477074 44604 477076
rect 80004 477074 80604 477076
rect 116004 477074 116604 477076
rect 152004 477074 152604 477076
rect 188004 477074 188604 477076
rect 224004 477074 224604 477076
rect 260004 477074 260604 477076
rect 296004 477074 296604 477076
rect 332004 477074 332604 477076
rect 368004 477074 368604 477076
rect 404004 477074 404604 477076
rect 440004 477074 440604 477076
rect 476004 477074 476604 477076
rect 512004 477074 512604 477076
rect 548004 477074 548604 477076
rect 589000 477074 589600 477076
rect -3836 474076 -3236 474078
rect 4404 474076 5004 474078
rect 40404 474076 41004 474078
rect 76404 474076 77004 474078
rect 112404 474076 113004 474078
rect 148404 474076 149004 474078
rect 184404 474076 185004 474078
rect 220404 474076 221004 474078
rect 256404 474076 257004 474078
rect 292404 474076 293004 474078
rect 328404 474076 329004 474078
rect 364404 474076 365004 474078
rect 400404 474076 401004 474078
rect 436404 474076 437004 474078
rect 472404 474076 473004 474078
rect 508404 474076 509004 474078
rect 544404 474076 545004 474078
rect 580404 474076 581004 474078
rect 587160 474076 587760 474078
rect -4756 474054 588680 474076
rect -4756 473818 -3654 474054
rect -3418 473818 4586 474054
rect 4822 473818 40586 474054
rect 40822 473818 76586 474054
rect 76822 473818 112586 474054
rect 112822 473818 148586 474054
rect 148822 473818 184586 474054
rect 184822 473818 220586 474054
rect 220822 473818 256586 474054
rect 256822 473818 292586 474054
rect 292822 473818 328586 474054
rect 328822 473818 364586 474054
rect 364822 473818 400586 474054
rect 400822 473818 436586 474054
rect 436822 473818 472586 474054
rect 472822 473818 508586 474054
rect 508822 473818 544586 474054
rect 544822 473818 580586 474054
rect 580822 473818 587342 474054
rect 587578 473818 588680 474054
rect -4756 473734 588680 473818
rect -4756 473498 -3654 473734
rect -3418 473498 4586 473734
rect 4822 473498 40586 473734
rect 40822 473498 76586 473734
rect 76822 473498 112586 473734
rect 112822 473498 148586 473734
rect 148822 473498 184586 473734
rect 184822 473498 220586 473734
rect 220822 473498 256586 473734
rect 256822 473498 292586 473734
rect 292822 473498 328586 473734
rect 328822 473498 364586 473734
rect 364822 473498 400586 473734
rect 400822 473498 436586 473734
rect 436822 473498 472586 473734
rect 472822 473498 508586 473734
rect 508822 473498 544586 473734
rect 544822 473498 580586 473734
rect 580822 473498 587342 473734
rect 587578 473498 588680 473734
rect -4756 473476 588680 473498
rect -3836 473474 -3236 473476
rect 4404 473474 5004 473476
rect 40404 473474 41004 473476
rect 76404 473474 77004 473476
rect 112404 473474 113004 473476
rect 148404 473474 149004 473476
rect 184404 473474 185004 473476
rect 220404 473474 221004 473476
rect 256404 473474 257004 473476
rect 292404 473474 293004 473476
rect 328404 473474 329004 473476
rect 364404 473474 365004 473476
rect 400404 473474 401004 473476
rect 436404 473474 437004 473476
rect 472404 473474 473004 473476
rect 508404 473474 509004 473476
rect 544404 473474 545004 473476
rect 580404 473474 581004 473476
rect 587160 473474 587760 473476
rect -1996 470476 -1396 470478
rect 804 470476 1404 470478
rect 36804 470476 37404 470478
rect 72804 470476 73404 470478
rect 108804 470476 109404 470478
rect 144804 470476 145404 470478
rect 180804 470476 181404 470478
rect 216804 470476 217404 470478
rect 252804 470476 253404 470478
rect 288804 470476 289404 470478
rect 324804 470476 325404 470478
rect 360804 470476 361404 470478
rect 396804 470476 397404 470478
rect 432804 470476 433404 470478
rect 468804 470476 469404 470478
rect 504804 470476 505404 470478
rect 540804 470476 541404 470478
rect 576804 470476 577404 470478
rect 585320 470476 585920 470478
rect -2916 470454 586840 470476
rect -2916 470218 -1814 470454
rect -1578 470218 986 470454
rect 1222 470218 36986 470454
rect 37222 470218 72986 470454
rect 73222 470218 108986 470454
rect 109222 470218 144986 470454
rect 145222 470218 180986 470454
rect 181222 470218 216986 470454
rect 217222 470218 252986 470454
rect 253222 470218 288986 470454
rect 289222 470218 324986 470454
rect 325222 470218 360986 470454
rect 361222 470218 396986 470454
rect 397222 470218 432986 470454
rect 433222 470218 468986 470454
rect 469222 470218 504986 470454
rect 505222 470218 540986 470454
rect 541222 470218 576986 470454
rect 577222 470218 585502 470454
rect 585738 470218 586840 470454
rect -2916 470134 586840 470218
rect -2916 469898 -1814 470134
rect -1578 469898 986 470134
rect 1222 469898 36986 470134
rect 37222 469898 72986 470134
rect 73222 469898 108986 470134
rect 109222 469898 144986 470134
rect 145222 469898 180986 470134
rect 181222 469898 216986 470134
rect 217222 469898 252986 470134
rect 253222 469898 288986 470134
rect 289222 469898 324986 470134
rect 325222 469898 360986 470134
rect 361222 469898 396986 470134
rect 397222 469898 432986 470134
rect 433222 469898 468986 470134
rect 469222 469898 504986 470134
rect 505222 469898 540986 470134
rect 541222 469898 576986 470134
rect 577222 469898 585502 470134
rect 585738 469898 586840 470134
rect -2916 469876 586840 469898
rect -1996 469874 -1396 469876
rect 804 469874 1404 469876
rect 36804 469874 37404 469876
rect 72804 469874 73404 469876
rect 108804 469874 109404 469876
rect 144804 469874 145404 469876
rect 180804 469874 181404 469876
rect 216804 469874 217404 469876
rect 252804 469874 253404 469876
rect 288804 469874 289404 469876
rect 324804 469874 325404 469876
rect 360804 469874 361404 469876
rect 396804 469874 397404 469876
rect 432804 469874 433404 469876
rect 468804 469874 469404 469876
rect 504804 469874 505404 469876
rect 540804 469874 541404 469876
rect 576804 469874 577404 469876
rect 585320 469874 585920 469876
rect -8436 463276 -7836 463278
rect 29604 463276 30204 463278
rect 65604 463276 66204 463278
rect 101604 463276 102204 463278
rect 137604 463276 138204 463278
rect 173604 463276 174204 463278
rect 209604 463276 210204 463278
rect 245604 463276 246204 463278
rect 281604 463276 282204 463278
rect 317604 463276 318204 463278
rect 353604 463276 354204 463278
rect 389604 463276 390204 463278
rect 425604 463276 426204 463278
rect 461604 463276 462204 463278
rect 497604 463276 498204 463278
rect 533604 463276 534204 463278
rect 569604 463276 570204 463278
rect 591760 463276 592360 463278
rect -8436 463254 592360 463276
rect -8436 463018 -8254 463254
rect -8018 463018 29786 463254
rect 30022 463018 65786 463254
rect 66022 463018 101786 463254
rect 102022 463018 137786 463254
rect 138022 463018 173786 463254
rect 174022 463018 209786 463254
rect 210022 463018 245786 463254
rect 246022 463018 281786 463254
rect 282022 463018 317786 463254
rect 318022 463018 353786 463254
rect 354022 463018 389786 463254
rect 390022 463018 425786 463254
rect 426022 463018 461786 463254
rect 462022 463018 497786 463254
rect 498022 463018 533786 463254
rect 534022 463018 569786 463254
rect 570022 463018 591942 463254
rect 592178 463018 592360 463254
rect -8436 462934 592360 463018
rect -8436 462698 -8254 462934
rect -8018 462698 29786 462934
rect 30022 462698 65786 462934
rect 66022 462698 101786 462934
rect 102022 462698 137786 462934
rect 138022 462698 173786 462934
rect 174022 462698 209786 462934
rect 210022 462698 245786 462934
rect 246022 462698 281786 462934
rect 282022 462698 317786 462934
rect 318022 462698 353786 462934
rect 354022 462698 389786 462934
rect 390022 462698 425786 462934
rect 426022 462698 461786 462934
rect 462022 462698 497786 462934
rect 498022 462698 533786 462934
rect 534022 462698 569786 462934
rect 570022 462698 591942 462934
rect 592178 462698 592360 462934
rect -8436 462676 592360 462698
rect -8436 462674 -7836 462676
rect 29604 462674 30204 462676
rect 65604 462674 66204 462676
rect 101604 462674 102204 462676
rect 137604 462674 138204 462676
rect 173604 462674 174204 462676
rect 209604 462674 210204 462676
rect 245604 462674 246204 462676
rect 281604 462674 282204 462676
rect 317604 462674 318204 462676
rect 353604 462674 354204 462676
rect 389604 462674 390204 462676
rect 425604 462674 426204 462676
rect 461604 462674 462204 462676
rect 497604 462674 498204 462676
rect 533604 462674 534204 462676
rect 569604 462674 570204 462676
rect 591760 462674 592360 462676
rect -6596 459676 -5996 459678
rect 26004 459676 26604 459678
rect 62004 459676 62604 459678
rect 98004 459676 98604 459678
rect 134004 459676 134604 459678
rect 170004 459676 170604 459678
rect 206004 459676 206604 459678
rect 242004 459676 242604 459678
rect 278004 459676 278604 459678
rect 314004 459676 314604 459678
rect 350004 459676 350604 459678
rect 386004 459676 386604 459678
rect 422004 459676 422604 459678
rect 458004 459676 458604 459678
rect 494004 459676 494604 459678
rect 530004 459676 530604 459678
rect 566004 459676 566604 459678
rect 589920 459676 590520 459678
rect -6596 459654 590520 459676
rect -6596 459418 -6414 459654
rect -6178 459418 26186 459654
rect 26422 459418 62186 459654
rect 62422 459418 98186 459654
rect 98422 459418 134186 459654
rect 134422 459418 170186 459654
rect 170422 459418 206186 459654
rect 206422 459418 242186 459654
rect 242422 459418 278186 459654
rect 278422 459418 314186 459654
rect 314422 459418 350186 459654
rect 350422 459418 386186 459654
rect 386422 459418 422186 459654
rect 422422 459418 458186 459654
rect 458422 459418 494186 459654
rect 494422 459418 530186 459654
rect 530422 459418 566186 459654
rect 566422 459418 590102 459654
rect 590338 459418 590520 459654
rect -6596 459334 590520 459418
rect -6596 459098 -6414 459334
rect -6178 459098 26186 459334
rect 26422 459098 62186 459334
rect 62422 459098 98186 459334
rect 98422 459098 134186 459334
rect 134422 459098 170186 459334
rect 170422 459098 206186 459334
rect 206422 459098 242186 459334
rect 242422 459098 278186 459334
rect 278422 459098 314186 459334
rect 314422 459098 350186 459334
rect 350422 459098 386186 459334
rect 386422 459098 422186 459334
rect 422422 459098 458186 459334
rect 458422 459098 494186 459334
rect 494422 459098 530186 459334
rect 530422 459098 566186 459334
rect 566422 459098 590102 459334
rect 590338 459098 590520 459334
rect -6596 459076 590520 459098
rect -6596 459074 -5996 459076
rect 26004 459074 26604 459076
rect 62004 459074 62604 459076
rect 98004 459074 98604 459076
rect 134004 459074 134604 459076
rect 170004 459074 170604 459076
rect 206004 459074 206604 459076
rect 242004 459074 242604 459076
rect 278004 459074 278604 459076
rect 314004 459074 314604 459076
rect 350004 459074 350604 459076
rect 386004 459074 386604 459076
rect 422004 459074 422604 459076
rect 458004 459074 458604 459076
rect 494004 459074 494604 459076
rect 530004 459074 530604 459076
rect 566004 459074 566604 459076
rect 589920 459074 590520 459076
rect -4756 456076 -4156 456078
rect 22404 456076 23004 456078
rect 58404 456076 59004 456078
rect 94404 456076 95004 456078
rect 130404 456076 131004 456078
rect 166404 456076 167004 456078
rect 202404 456076 203004 456078
rect 238404 456076 239004 456078
rect 274404 456076 275004 456078
rect 310404 456076 311004 456078
rect 346404 456076 347004 456078
rect 382404 456076 383004 456078
rect 418404 456076 419004 456078
rect 454404 456076 455004 456078
rect 490404 456076 491004 456078
rect 526404 456076 527004 456078
rect 562404 456076 563004 456078
rect 588080 456076 588680 456078
rect -4756 456054 588680 456076
rect -4756 455818 -4574 456054
rect -4338 455818 22586 456054
rect 22822 455818 58586 456054
rect 58822 455818 94586 456054
rect 94822 455818 130586 456054
rect 130822 455818 166586 456054
rect 166822 455818 202586 456054
rect 202822 455818 238586 456054
rect 238822 455818 274586 456054
rect 274822 455818 310586 456054
rect 310822 455818 346586 456054
rect 346822 455818 382586 456054
rect 382822 455818 418586 456054
rect 418822 455818 454586 456054
rect 454822 455818 490586 456054
rect 490822 455818 526586 456054
rect 526822 455818 562586 456054
rect 562822 455818 588262 456054
rect 588498 455818 588680 456054
rect -4756 455734 588680 455818
rect -4756 455498 -4574 455734
rect -4338 455498 22586 455734
rect 22822 455498 58586 455734
rect 58822 455498 94586 455734
rect 94822 455498 130586 455734
rect 130822 455498 166586 455734
rect 166822 455498 202586 455734
rect 202822 455498 238586 455734
rect 238822 455498 274586 455734
rect 274822 455498 310586 455734
rect 310822 455498 346586 455734
rect 346822 455498 382586 455734
rect 382822 455498 418586 455734
rect 418822 455498 454586 455734
rect 454822 455498 490586 455734
rect 490822 455498 526586 455734
rect 526822 455498 562586 455734
rect 562822 455498 588262 455734
rect 588498 455498 588680 455734
rect -4756 455476 588680 455498
rect -4756 455474 -4156 455476
rect 22404 455474 23004 455476
rect 58404 455474 59004 455476
rect 94404 455474 95004 455476
rect 130404 455474 131004 455476
rect 166404 455474 167004 455476
rect 202404 455474 203004 455476
rect 238404 455474 239004 455476
rect 274404 455474 275004 455476
rect 310404 455474 311004 455476
rect 346404 455474 347004 455476
rect 382404 455474 383004 455476
rect 418404 455474 419004 455476
rect 454404 455474 455004 455476
rect 490404 455474 491004 455476
rect 526404 455474 527004 455476
rect 562404 455474 563004 455476
rect 588080 455474 588680 455476
rect -2916 452476 -2316 452478
rect 18804 452476 19404 452478
rect 54804 452476 55404 452478
rect 90804 452476 91404 452478
rect 126804 452476 127404 452478
rect 162804 452476 163404 452478
rect 198804 452476 199404 452478
rect 234804 452476 235404 452478
rect 270804 452476 271404 452478
rect 306804 452476 307404 452478
rect 342804 452476 343404 452478
rect 378804 452476 379404 452478
rect 414804 452476 415404 452478
rect 450804 452476 451404 452478
rect 486804 452476 487404 452478
rect 522804 452476 523404 452478
rect 558804 452476 559404 452478
rect 586240 452476 586840 452478
rect -2916 452454 586840 452476
rect -2916 452218 -2734 452454
rect -2498 452218 18986 452454
rect 19222 452218 54986 452454
rect 55222 452218 90986 452454
rect 91222 452218 126986 452454
rect 127222 452218 162986 452454
rect 163222 452218 198986 452454
rect 199222 452218 234986 452454
rect 235222 452218 270986 452454
rect 271222 452218 306986 452454
rect 307222 452218 342986 452454
rect 343222 452218 378986 452454
rect 379222 452218 414986 452454
rect 415222 452218 450986 452454
rect 451222 452218 486986 452454
rect 487222 452218 522986 452454
rect 523222 452218 558986 452454
rect 559222 452218 586422 452454
rect 586658 452218 586840 452454
rect -2916 452134 586840 452218
rect -2916 451898 -2734 452134
rect -2498 451898 18986 452134
rect 19222 451898 54986 452134
rect 55222 451898 90986 452134
rect 91222 451898 126986 452134
rect 127222 451898 162986 452134
rect 163222 451898 198986 452134
rect 199222 451898 234986 452134
rect 235222 451898 270986 452134
rect 271222 451898 306986 452134
rect 307222 451898 342986 452134
rect 343222 451898 378986 452134
rect 379222 451898 414986 452134
rect 415222 451898 450986 452134
rect 451222 451898 486986 452134
rect 487222 451898 522986 452134
rect 523222 451898 558986 452134
rect 559222 451898 586422 452134
rect 586658 451898 586840 452134
rect -2916 451876 586840 451898
rect -2916 451874 -2316 451876
rect 18804 451874 19404 451876
rect 54804 451874 55404 451876
rect 90804 451874 91404 451876
rect 126804 451874 127404 451876
rect 162804 451874 163404 451876
rect 198804 451874 199404 451876
rect 234804 451874 235404 451876
rect 270804 451874 271404 451876
rect 306804 451874 307404 451876
rect 342804 451874 343404 451876
rect 378804 451874 379404 451876
rect 414804 451874 415404 451876
rect 450804 451874 451404 451876
rect 486804 451874 487404 451876
rect 522804 451874 523404 451876
rect 558804 451874 559404 451876
rect 586240 451874 586840 451876
rect -7516 445276 -6916 445278
rect 11604 445276 12204 445278
rect 47604 445276 48204 445278
rect 83604 445276 84204 445278
rect 119604 445276 120204 445278
rect 155604 445276 156204 445278
rect 191604 445276 192204 445278
rect 227604 445276 228204 445278
rect 263604 445276 264204 445278
rect 299604 445276 300204 445278
rect 335604 445276 336204 445278
rect 371604 445276 372204 445278
rect 407604 445276 408204 445278
rect 443604 445276 444204 445278
rect 479604 445276 480204 445278
rect 515604 445276 516204 445278
rect 551604 445276 552204 445278
rect 590840 445276 591440 445278
rect -8436 445254 592360 445276
rect -8436 445018 -7334 445254
rect -7098 445018 11786 445254
rect 12022 445018 47786 445254
rect 48022 445018 83786 445254
rect 84022 445018 119786 445254
rect 120022 445018 155786 445254
rect 156022 445018 191786 445254
rect 192022 445018 227786 445254
rect 228022 445018 263786 445254
rect 264022 445018 299786 445254
rect 300022 445018 335786 445254
rect 336022 445018 371786 445254
rect 372022 445018 407786 445254
rect 408022 445018 443786 445254
rect 444022 445018 479786 445254
rect 480022 445018 515786 445254
rect 516022 445018 551786 445254
rect 552022 445018 591022 445254
rect 591258 445018 592360 445254
rect -8436 444934 592360 445018
rect -8436 444698 -7334 444934
rect -7098 444698 11786 444934
rect 12022 444698 47786 444934
rect 48022 444698 83786 444934
rect 84022 444698 119786 444934
rect 120022 444698 155786 444934
rect 156022 444698 191786 444934
rect 192022 444698 227786 444934
rect 228022 444698 263786 444934
rect 264022 444698 299786 444934
rect 300022 444698 335786 444934
rect 336022 444698 371786 444934
rect 372022 444698 407786 444934
rect 408022 444698 443786 444934
rect 444022 444698 479786 444934
rect 480022 444698 515786 444934
rect 516022 444698 551786 444934
rect 552022 444698 591022 444934
rect 591258 444698 592360 444934
rect -8436 444676 592360 444698
rect -7516 444674 -6916 444676
rect 11604 444674 12204 444676
rect 47604 444674 48204 444676
rect 83604 444674 84204 444676
rect 119604 444674 120204 444676
rect 155604 444674 156204 444676
rect 191604 444674 192204 444676
rect 227604 444674 228204 444676
rect 263604 444674 264204 444676
rect 299604 444674 300204 444676
rect 335604 444674 336204 444676
rect 371604 444674 372204 444676
rect 407604 444674 408204 444676
rect 443604 444674 444204 444676
rect 479604 444674 480204 444676
rect 515604 444674 516204 444676
rect 551604 444674 552204 444676
rect 590840 444674 591440 444676
rect -5676 441676 -5076 441678
rect 8004 441676 8604 441678
rect 44004 441676 44604 441678
rect 80004 441676 80604 441678
rect 116004 441676 116604 441678
rect 152004 441676 152604 441678
rect 188004 441676 188604 441678
rect 224004 441676 224604 441678
rect 260004 441676 260604 441678
rect 296004 441676 296604 441678
rect 332004 441676 332604 441678
rect 368004 441676 368604 441678
rect 404004 441676 404604 441678
rect 440004 441676 440604 441678
rect 476004 441676 476604 441678
rect 512004 441676 512604 441678
rect 548004 441676 548604 441678
rect 589000 441676 589600 441678
rect -6596 441654 590520 441676
rect -6596 441418 -5494 441654
rect -5258 441418 8186 441654
rect 8422 441418 44186 441654
rect 44422 441418 80186 441654
rect 80422 441418 116186 441654
rect 116422 441418 152186 441654
rect 152422 441418 188186 441654
rect 188422 441418 224186 441654
rect 224422 441418 260186 441654
rect 260422 441418 296186 441654
rect 296422 441418 332186 441654
rect 332422 441418 368186 441654
rect 368422 441418 404186 441654
rect 404422 441418 440186 441654
rect 440422 441418 476186 441654
rect 476422 441418 512186 441654
rect 512422 441418 548186 441654
rect 548422 441418 589182 441654
rect 589418 441418 590520 441654
rect -6596 441334 590520 441418
rect -6596 441098 -5494 441334
rect -5258 441098 8186 441334
rect 8422 441098 44186 441334
rect 44422 441098 80186 441334
rect 80422 441098 116186 441334
rect 116422 441098 152186 441334
rect 152422 441098 188186 441334
rect 188422 441098 224186 441334
rect 224422 441098 260186 441334
rect 260422 441098 296186 441334
rect 296422 441098 332186 441334
rect 332422 441098 368186 441334
rect 368422 441098 404186 441334
rect 404422 441098 440186 441334
rect 440422 441098 476186 441334
rect 476422 441098 512186 441334
rect 512422 441098 548186 441334
rect 548422 441098 589182 441334
rect 589418 441098 590520 441334
rect -6596 441076 590520 441098
rect -5676 441074 -5076 441076
rect 8004 441074 8604 441076
rect 44004 441074 44604 441076
rect 80004 441074 80604 441076
rect 116004 441074 116604 441076
rect 152004 441074 152604 441076
rect 188004 441074 188604 441076
rect 224004 441074 224604 441076
rect 260004 441074 260604 441076
rect 296004 441074 296604 441076
rect 332004 441074 332604 441076
rect 368004 441074 368604 441076
rect 404004 441074 404604 441076
rect 440004 441074 440604 441076
rect 476004 441074 476604 441076
rect 512004 441074 512604 441076
rect 548004 441074 548604 441076
rect 589000 441074 589600 441076
rect -3836 438076 -3236 438078
rect 4404 438076 5004 438078
rect 40404 438076 41004 438078
rect 76404 438076 77004 438078
rect 112404 438076 113004 438078
rect 148404 438076 149004 438078
rect 184404 438076 185004 438078
rect 220404 438076 221004 438078
rect 256404 438076 257004 438078
rect 292404 438076 293004 438078
rect 328404 438076 329004 438078
rect 364404 438076 365004 438078
rect 400404 438076 401004 438078
rect 436404 438076 437004 438078
rect 472404 438076 473004 438078
rect 508404 438076 509004 438078
rect 544404 438076 545004 438078
rect 580404 438076 581004 438078
rect 587160 438076 587760 438078
rect -4756 438054 588680 438076
rect -4756 437818 -3654 438054
rect -3418 437818 4586 438054
rect 4822 437818 40586 438054
rect 40822 437818 76586 438054
rect 76822 437818 112586 438054
rect 112822 437818 148586 438054
rect 148822 437818 184586 438054
rect 184822 437818 220586 438054
rect 220822 437818 256586 438054
rect 256822 437818 292586 438054
rect 292822 437818 328586 438054
rect 328822 437818 364586 438054
rect 364822 437818 400586 438054
rect 400822 437818 436586 438054
rect 436822 437818 472586 438054
rect 472822 437818 508586 438054
rect 508822 437818 544586 438054
rect 544822 437818 580586 438054
rect 580822 437818 587342 438054
rect 587578 437818 588680 438054
rect -4756 437734 588680 437818
rect -4756 437498 -3654 437734
rect -3418 437498 4586 437734
rect 4822 437498 40586 437734
rect 40822 437498 76586 437734
rect 76822 437498 112586 437734
rect 112822 437498 148586 437734
rect 148822 437498 184586 437734
rect 184822 437498 220586 437734
rect 220822 437498 256586 437734
rect 256822 437498 292586 437734
rect 292822 437498 328586 437734
rect 328822 437498 364586 437734
rect 364822 437498 400586 437734
rect 400822 437498 436586 437734
rect 436822 437498 472586 437734
rect 472822 437498 508586 437734
rect 508822 437498 544586 437734
rect 544822 437498 580586 437734
rect 580822 437498 587342 437734
rect 587578 437498 588680 437734
rect -4756 437476 588680 437498
rect -3836 437474 -3236 437476
rect 4404 437474 5004 437476
rect 40404 437474 41004 437476
rect 76404 437474 77004 437476
rect 112404 437474 113004 437476
rect 148404 437474 149004 437476
rect 184404 437474 185004 437476
rect 220404 437474 221004 437476
rect 256404 437474 257004 437476
rect 292404 437474 293004 437476
rect 328404 437474 329004 437476
rect 364404 437474 365004 437476
rect 400404 437474 401004 437476
rect 436404 437474 437004 437476
rect 472404 437474 473004 437476
rect 508404 437474 509004 437476
rect 544404 437474 545004 437476
rect 580404 437474 581004 437476
rect 587160 437474 587760 437476
rect -1996 434476 -1396 434478
rect 804 434476 1404 434478
rect 36804 434476 37404 434478
rect 72804 434476 73404 434478
rect 108804 434476 109404 434478
rect 144804 434476 145404 434478
rect 180804 434476 181404 434478
rect 216804 434476 217404 434478
rect 252804 434476 253404 434478
rect 288804 434476 289404 434478
rect 324804 434476 325404 434478
rect 360804 434476 361404 434478
rect 396804 434476 397404 434478
rect 432804 434476 433404 434478
rect 468804 434476 469404 434478
rect 504804 434476 505404 434478
rect 540804 434476 541404 434478
rect 576804 434476 577404 434478
rect 585320 434476 585920 434478
rect -2916 434454 586840 434476
rect -2916 434218 -1814 434454
rect -1578 434218 986 434454
rect 1222 434218 36986 434454
rect 37222 434218 72986 434454
rect 73222 434218 108986 434454
rect 109222 434218 144986 434454
rect 145222 434218 180986 434454
rect 181222 434218 216986 434454
rect 217222 434218 252986 434454
rect 253222 434218 288986 434454
rect 289222 434218 324986 434454
rect 325222 434218 360986 434454
rect 361222 434218 396986 434454
rect 397222 434218 432986 434454
rect 433222 434218 468986 434454
rect 469222 434218 504986 434454
rect 505222 434218 540986 434454
rect 541222 434218 576986 434454
rect 577222 434218 585502 434454
rect 585738 434218 586840 434454
rect -2916 434134 586840 434218
rect -2916 433898 -1814 434134
rect -1578 433898 986 434134
rect 1222 433898 36986 434134
rect 37222 433898 72986 434134
rect 73222 433898 108986 434134
rect 109222 433898 144986 434134
rect 145222 433898 180986 434134
rect 181222 433898 216986 434134
rect 217222 433898 252986 434134
rect 253222 433898 288986 434134
rect 289222 433898 324986 434134
rect 325222 433898 360986 434134
rect 361222 433898 396986 434134
rect 397222 433898 432986 434134
rect 433222 433898 468986 434134
rect 469222 433898 504986 434134
rect 505222 433898 540986 434134
rect 541222 433898 576986 434134
rect 577222 433898 585502 434134
rect 585738 433898 586840 434134
rect -2916 433876 586840 433898
rect -1996 433874 -1396 433876
rect 804 433874 1404 433876
rect 36804 433874 37404 433876
rect 72804 433874 73404 433876
rect 108804 433874 109404 433876
rect 144804 433874 145404 433876
rect 180804 433874 181404 433876
rect 216804 433874 217404 433876
rect 252804 433874 253404 433876
rect 288804 433874 289404 433876
rect 324804 433874 325404 433876
rect 360804 433874 361404 433876
rect 396804 433874 397404 433876
rect 432804 433874 433404 433876
rect 468804 433874 469404 433876
rect 504804 433874 505404 433876
rect 540804 433874 541404 433876
rect 576804 433874 577404 433876
rect 585320 433874 585920 433876
rect -8436 427276 -7836 427278
rect 29604 427276 30204 427278
rect 65604 427276 66204 427278
rect 101604 427276 102204 427278
rect 137604 427276 138204 427278
rect 173604 427276 174204 427278
rect 209604 427276 210204 427278
rect 245604 427276 246204 427278
rect 281604 427276 282204 427278
rect 317604 427276 318204 427278
rect 353604 427276 354204 427278
rect 389604 427276 390204 427278
rect 425604 427276 426204 427278
rect 461604 427276 462204 427278
rect 497604 427276 498204 427278
rect 533604 427276 534204 427278
rect 569604 427276 570204 427278
rect 591760 427276 592360 427278
rect -8436 427254 592360 427276
rect -8436 427018 -8254 427254
rect -8018 427018 29786 427254
rect 30022 427018 65786 427254
rect 66022 427018 101786 427254
rect 102022 427018 137786 427254
rect 138022 427018 173786 427254
rect 174022 427018 209786 427254
rect 210022 427018 245786 427254
rect 246022 427018 281786 427254
rect 282022 427018 317786 427254
rect 318022 427018 353786 427254
rect 354022 427018 389786 427254
rect 390022 427018 425786 427254
rect 426022 427018 461786 427254
rect 462022 427018 497786 427254
rect 498022 427018 533786 427254
rect 534022 427018 569786 427254
rect 570022 427018 591942 427254
rect 592178 427018 592360 427254
rect -8436 426934 592360 427018
rect -8436 426698 -8254 426934
rect -8018 426698 29786 426934
rect 30022 426698 65786 426934
rect 66022 426698 101786 426934
rect 102022 426698 137786 426934
rect 138022 426698 173786 426934
rect 174022 426698 209786 426934
rect 210022 426698 245786 426934
rect 246022 426698 281786 426934
rect 282022 426698 317786 426934
rect 318022 426698 353786 426934
rect 354022 426698 389786 426934
rect 390022 426698 425786 426934
rect 426022 426698 461786 426934
rect 462022 426698 497786 426934
rect 498022 426698 533786 426934
rect 534022 426698 569786 426934
rect 570022 426698 591942 426934
rect 592178 426698 592360 426934
rect -8436 426676 592360 426698
rect -8436 426674 -7836 426676
rect 29604 426674 30204 426676
rect 65604 426674 66204 426676
rect 101604 426674 102204 426676
rect 137604 426674 138204 426676
rect 173604 426674 174204 426676
rect 209604 426674 210204 426676
rect 245604 426674 246204 426676
rect 281604 426674 282204 426676
rect 317604 426674 318204 426676
rect 353604 426674 354204 426676
rect 389604 426674 390204 426676
rect 425604 426674 426204 426676
rect 461604 426674 462204 426676
rect 497604 426674 498204 426676
rect 533604 426674 534204 426676
rect 569604 426674 570204 426676
rect 591760 426674 592360 426676
rect -6596 423676 -5996 423678
rect 26004 423676 26604 423678
rect 62004 423676 62604 423678
rect 98004 423676 98604 423678
rect 134004 423676 134604 423678
rect 170004 423676 170604 423678
rect 206004 423676 206604 423678
rect 242004 423676 242604 423678
rect 278004 423676 278604 423678
rect 314004 423676 314604 423678
rect 350004 423676 350604 423678
rect 386004 423676 386604 423678
rect 422004 423676 422604 423678
rect 458004 423676 458604 423678
rect 494004 423676 494604 423678
rect 530004 423676 530604 423678
rect 566004 423676 566604 423678
rect 589920 423676 590520 423678
rect -6596 423654 590520 423676
rect -6596 423418 -6414 423654
rect -6178 423418 26186 423654
rect 26422 423418 62186 423654
rect 62422 423418 98186 423654
rect 98422 423418 134186 423654
rect 134422 423418 170186 423654
rect 170422 423418 206186 423654
rect 206422 423418 242186 423654
rect 242422 423418 278186 423654
rect 278422 423418 314186 423654
rect 314422 423418 350186 423654
rect 350422 423418 386186 423654
rect 386422 423418 422186 423654
rect 422422 423418 458186 423654
rect 458422 423418 494186 423654
rect 494422 423418 530186 423654
rect 530422 423418 566186 423654
rect 566422 423418 590102 423654
rect 590338 423418 590520 423654
rect -6596 423334 590520 423418
rect -6596 423098 -6414 423334
rect -6178 423098 26186 423334
rect 26422 423098 62186 423334
rect 62422 423098 98186 423334
rect 98422 423098 134186 423334
rect 134422 423098 170186 423334
rect 170422 423098 206186 423334
rect 206422 423098 242186 423334
rect 242422 423098 278186 423334
rect 278422 423098 314186 423334
rect 314422 423098 350186 423334
rect 350422 423098 386186 423334
rect 386422 423098 422186 423334
rect 422422 423098 458186 423334
rect 458422 423098 494186 423334
rect 494422 423098 530186 423334
rect 530422 423098 566186 423334
rect 566422 423098 590102 423334
rect 590338 423098 590520 423334
rect -6596 423076 590520 423098
rect -6596 423074 -5996 423076
rect 26004 423074 26604 423076
rect 62004 423074 62604 423076
rect 98004 423074 98604 423076
rect 134004 423074 134604 423076
rect 170004 423074 170604 423076
rect 206004 423074 206604 423076
rect 242004 423074 242604 423076
rect 278004 423074 278604 423076
rect 314004 423074 314604 423076
rect 350004 423074 350604 423076
rect 386004 423074 386604 423076
rect 422004 423074 422604 423076
rect 458004 423074 458604 423076
rect 494004 423074 494604 423076
rect 530004 423074 530604 423076
rect 566004 423074 566604 423076
rect 589920 423074 590520 423076
rect -4756 420076 -4156 420078
rect 22404 420076 23004 420078
rect 58404 420076 59004 420078
rect 94404 420076 95004 420078
rect 130404 420076 131004 420078
rect 166404 420076 167004 420078
rect 202404 420076 203004 420078
rect 238404 420076 239004 420078
rect 274404 420076 275004 420078
rect 310404 420076 311004 420078
rect 346404 420076 347004 420078
rect 382404 420076 383004 420078
rect 418404 420076 419004 420078
rect 454404 420076 455004 420078
rect 490404 420076 491004 420078
rect 526404 420076 527004 420078
rect 562404 420076 563004 420078
rect 588080 420076 588680 420078
rect -4756 420054 588680 420076
rect -4756 419818 -4574 420054
rect -4338 419818 22586 420054
rect 22822 419818 58586 420054
rect 58822 419818 94586 420054
rect 94822 419818 130586 420054
rect 130822 419818 166586 420054
rect 166822 419818 202586 420054
rect 202822 419818 238586 420054
rect 238822 419818 274586 420054
rect 274822 419818 310586 420054
rect 310822 419818 346586 420054
rect 346822 419818 382586 420054
rect 382822 419818 418586 420054
rect 418822 419818 454586 420054
rect 454822 419818 490586 420054
rect 490822 419818 526586 420054
rect 526822 419818 562586 420054
rect 562822 419818 588262 420054
rect 588498 419818 588680 420054
rect -4756 419734 588680 419818
rect -4756 419498 -4574 419734
rect -4338 419498 22586 419734
rect 22822 419498 58586 419734
rect 58822 419498 94586 419734
rect 94822 419498 130586 419734
rect 130822 419498 166586 419734
rect 166822 419498 202586 419734
rect 202822 419498 238586 419734
rect 238822 419498 274586 419734
rect 274822 419498 310586 419734
rect 310822 419498 346586 419734
rect 346822 419498 382586 419734
rect 382822 419498 418586 419734
rect 418822 419498 454586 419734
rect 454822 419498 490586 419734
rect 490822 419498 526586 419734
rect 526822 419498 562586 419734
rect 562822 419498 588262 419734
rect 588498 419498 588680 419734
rect -4756 419476 588680 419498
rect -4756 419474 -4156 419476
rect 22404 419474 23004 419476
rect 58404 419474 59004 419476
rect 94404 419474 95004 419476
rect 130404 419474 131004 419476
rect 166404 419474 167004 419476
rect 202404 419474 203004 419476
rect 238404 419474 239004 419476
rect 274404 419474 275004 419476
rect 310404 419474 311004 419476
rect 346404 419474 347004 419476
rect 382404 419474 383004 419476
rect 418404 419474 419004 419476
rect 454404 419474 455004 419476
rect 490404 419474 491004 419476
rect 526404 419474 527004 419476
rect 562404 419474 563004 419476
rect 588080 419474 588680 419476
rect -2916 416476 -2316 416478
rect 18804 416476 19404 416478
rect 54804 416476 55404 416478
rect 90804 416476 91404 416478
rect 126804 416476 127404 416478
rect 162804 416476 163404 416478
rect 198804 416476 199404 416478
rect 234804 416476 235404 416478
rect 270804 416476 271404 416478
rect 306804 416476 307404 416478
rect 342804 416476 343404 416478
rect 378804 416476 379404 416478
rect 414804 416476 415404 416478
rect 450804 416476 451404 416478
rect 486804 416476 487404 416478
rect 522804 416476 523404 416478
rect 558804 416476 559404 416478
rect 586240 416476 586840 416478
rect -2916 416454 586840 416476
rect -2916 416218 -2734 416454
rect -2498 416218 18986 416454
rect 19222 416218 54986 416454
rect 55222 416218 90986 416454
rect 91222 416218 126986 416454
rect 127222 416218 162986 416454
rect 163222 416218 198986 416454
rect 199222 416218 234986 416454
rect 235222 416218 270986 416454
rect 271222 416218 306986 416454
rect 307222 416218 342986 416454
rect 343222 416218 378986 416454
rect 379222 416218 414986 416454
rect 415222 416218 450986 416454
rect 451222 416218 486986 416454
rect 487222 416218 522986 416454
rect 523222 416218 558986 416454
rect 559222 416218 586422 416454
rect 586658 416218 586840 416454
rect -2916 416134 586840 416218
rect -2916 415898 -2734 416134
rect -2498 415898 18986 416134
rect 19222 415898 54986 416134
rect 55222 415898 90986 416134
rect 91222 415898 126986 416134
rect 127222 415898 162986 416134
rect 163222 415898 198986 416134
rect 199222 415898 234986 416134
rect 235222 415898 270986 416134
rect 271222 415898 306986 416134
rect 307222 415898 342986 416134
rect 343222 415898 378986 416134
rect 379222 415898 414986 416134
rect 415222 415898 450986 416134
rect 451222 415898 486986 416134
rect 487222 415898 522986 416134
rect 523222 415898 558986 416134
rect 559222 415898 586422 416134
rect 586658 415898 586840 416134
rect -2916 415876 586840 415898
rect -2916 415874 -2316 415876
rect 18804 415874 19404 415876
rect 54804 415874 55404 415876
rect 90804 415874 91404 415876
rect 126804 415874 127404 415876
rect 162804 415874 163404 415876
rect 198804 415874 199404 415876
rect 234804 415874 235404 415876
rect 270804 415874 271404 415876
rect 306804 415874 307404 415876
rect 342804 415874 343404 415876
rect 378804 415874 379404 415876
rect 414804 415874 415404 415876
rect 450804 415874 451404 415876
rect 486804 415874 487404 415876
rect 522804 415874 523404 415876
rect 558804 415874 559404 415876
rect 586240 415874 586840 415876
rect -7516 409276 -6916 409278
rect 11604 409276 12204 409278
rect 47604 409276 48204 409278
rect 83604 409276 84204 409278
rect 119604 409276 120204 409278
rect 155604 409276 156204 409278
rect 191604 409276 192204 409278
rect 227604 409276 228204 409278
rect 263604 409276 264204 409278
rect 299604 409276 300204 409278
rect 335604 409276 336204 409278
rect 371604 409276 372204 409278
rect 407604 409276 408204 409278
rect 443604 409276 444204 409278
rect 479604 409276 480204 409278
rect 515604 409276 516204 409278
rect 551604 409276 552204 409278
rect 590840 409276 591440 409278
rect -8436 409254 592360 409276
rect -8436 409018 -7334 409254
rect -7098 409018 11786 409254
rect 12022 409018 47786 409254
rect 48022 409018 83786 409254
rect 84022 409018 119786 409254
rect 120022 409018 155786 409254
rect 156022 409018 191786 409254
rect 192022 409018 227786 409254
rect 228022 409018 263786 409254
rect 264022 409018 299786 409254
rect 300022 409018 335786 409254
rect 336022 409018 371786 409254
rect 372022 409018 407786 409254
rect 408022 409018 443786 409254
rect 444022 409018 479786 409254
rect 480022 409018 515786 409254
rect 516022 409018 551786 409254
rect 552022 409018 591022 409254
rect 591258 409018 592360 409254
rect -8436 408934 592360 409018
rect -8436 408698 -7334 408934
rect -7098 408698 11786 408934
rect 12022 408698 47786 408934
rect 48022 408698 83786 408934
rect 84022 408698 119786 408934
rect 120022 408698 155786 408934
rect 156022 408698 191786 408934
rect 192022 408698 227786 408934
rect 228022 408698 263786 408934
rect 264022 408698 299786 408934
rect 300022 408698 335786 408934
rect 336022 408698 371786 408934
rect 372022 408698 407786 408934
rect 408022 408698 443786 408934
rect 444022 408698 479786 408934
rect 480022 408698 515786 408934
rect 516022 408698 551786 408934
rect 552022 408698 591022 408934
rect 591258 408698 592360 408934
rect -8436 408676 592360 408698
rect -7516 408674 -6916 408676
rect 11604 408674 12204 408676
rect 47604 408674 48204 408676
rect 83604 408674 84204 408676
rect 119604 408674 120204 408676
rect 155604 408674 156204 408676
rect 191604 408674 192204 408676
rect 227604 408674 228204 408676
rect 263604 408674 264204 408676
rect 299604 408674 300204 408676
rect 335604 408674 336204 408676
rect 371604 408674 372204 408676
rect 407604 408674 408204 408676
rect 443604 408674 444204 408676
rect 479604 408674 480204 408676
rect 515604 408674 516204 408676
rect 551604 408674 552204 408676
rect 590840 408674 591440 408676
rect -5676 405676 -5076 405678
rect 8004 405676 8604 405678
rect 44004 405676 44604 405678
rect 80004 405676 80604 405678
rect 116004 405676 116604 405678
rect 152004 405676 152604 405678
rect 188004 405676 188604 405678
rect 224004 405676 224604 405678
rect 260004 405676 260604 405678
rect 296004 405676 296604 405678
rect 332004 405676 332604 405678
rect 368004 405676 368604 405678
rect 404004 405676 404604 405678
rect 440004 405676 440604 405678
rect 476004 405676 476604 405678
rect 512004 405676 512604 405678
rect 548004 405676 548604 405678
rect 589000 405676 589600 405678
rect -6596 405654 590520 405676
rect -6596 405418 -5494 405654
rect -5258 405418 8186 405654
rect 8422 405418 44186 405654
rect 44422 405418 80186 405654
rect 80422 405418 116186 405654
rect 116422 405418 152186 405654
rect 152422 405418 188186 405654
rect 188422 405418 224186 405654
rect 224422 405418 260186 405654
rect 260422 405418 296186 405654
rect 296422 405418 332186 405654
rect 332422 405418 368186 405654
rect 368422 405418 404186 405654
rect 404422 405418 440186 405654
rect 440422 405418 476186 405654
rect 476422 405418 512186 405654
rect 512422 405418 548186 405654
rect 548422 405418 589182 405654
rect 589418 405418 590520 405654
rect -6596 405334 590520 405418
rect -6596 405098 -5494 405334
rect -5258 405098 8186 405334
rect 8422 405098 44186 405334
rect 44422 405098 80186 405334
rect 80422 405098 116186 405334
rect 116422 405098 152186 405334
rect 152422 405098 188186 405334
rect 188422 405098 224186 405334
rect 224422 405098 260186 405334
rect 260422 405098 296186 405334
rect 296422 405098 332186 405334
rect 332422 405098 368186 405334
rect 368422 405098 404186 405334
rect 404422 405098 440186 405334
rect 440422 405098 476186 405334
rect 476422 405098 512186 405334
rect 512422 405098 548186 405334
rect 548422 405098 589182 405334
rect 589418 405098 590520 405334
rect -6596 405076 590520 405098
rect -5676 405074 -5076 405076
rect 8004 405074 8604 405076
rect 44004 405074 44604 405076
rect 80004 405074 80604 405076
rect 116004 405074 116604 405076
rect 152004 405074 152604 405076
rect 188004 405074 188604 405076
rect 224004 405074 224604 405076
rect 260004 405074 260604 405076
rect 296004 405074 296604 405076
rect 332004 405074 332604 405076
rect 368004 405074 368604 405076
rect 404004 405074 404604 405076
rect 440004 405074 440604 405076
rect 476004 405074 476604 405076
rect 512004 405074 512604 405076
rect 548004 405074 548604 405076
rect 589000 405074 589600 405076
rect -3836 402076 -3236 402078
rect 4404 402076 5004 402078
rect 40404 402076 41004 402078
rect 76404 402076 77004 402078
rect 112404 402076 113004 402078
rect 148404 402076 149004 402078
rect 184404 402076 185004 402078
rect 220404 402076 221004 402078
rect 256404 402076 257004 402078
rect 292404 402076 293004 402078
rect 328404 402076 329004 402078
rect 364404 402076 365004 402078
rect 400404 402076 401004 402078
rect 436404 402076 437004 402078
rect 472404 402076 473004 402078
rect 508404 402076 509004 402078
rect 544404 402076 545004 402078
rect 580404 402076 581004 402078
rect 587160 402076 587760 402078
rect -4756 402054 588680 402076
rect -4756 401818 -3654 402054
rect -3418 401818 4586 402054
rect 4822 401818 40586 402054
rect 40822 401818 76586 402054
rect 76822 401818 112586 402054
rect 112822 401818 148586 402054
rect 148822 401818 184586 402054
rect 184822 401818 220586 402054
rect 220822 401818 256586 402054
rect 256822 401818 292586 402054
rect 292822 401818 328586 402054
rect 328822 401818 364586 402054
rect 364822 401818 400586 402054
rect 400822 401818 436586 402054
rect 436822 401818 472586 402054
rect 472822 401818 508586 402054
rect 508822 401818 544586 402054
rect 544822 401818 580586 402054
rect 580822 401818 587342 402054
rect 587578 401818 588680 402054
rect -4756 401734 588680 401818
rect -4756 401498 -3654 401734
rect -3418 401498 4586 401734
rect 4822 401498 40586 401734
rect 40822 401498 76586 401734
rect 76822 401498 112586 401734
rect 112822 401498 148586 401734
rect 148822 401498 184586 401734
rect 184822 401498 220586 401734
rect 220822 401498 256586 401734
rect 256822 401498 292586 401734
rect 292822 401498 328586 401734
rect 328822 401498 364586 401734
rect 364822 401498 400586 401734
rect 400822 401498 436586 401734
rect 436822 401498 472586 401734
rect 472822 401498 508586 401734
rect 508822 401498 544586 401734
rect 544822 401498 580586 401734
rect 580822 401498 587342 401734
rect 587578 401498 588680 401734
rect -4756 401476 588680 401498
rect -3836 401474 -3236 401476
rect 4404 401474 5004 401476
rect 40404 401474 41004 401476
rect 76404 401474 77004 401476
rect 112404 401474 113004 401476
rect 148404 401474 149004 401476
rect 184404 401474 185004 401476
rect 220404 401474 221004 401476
rect 256404 401474 257004 401476
rect 292404 401474 293004 401476
rect 328404 401474 329004 401476
rect 364404 401474 365004 401476
rect 400404 401474 401004 401476
rect 436404 401474 437004 401476
rect 472404 401474 473004 401476
rect 508404 401474 509004 401476
rect 544404 401474 545004 401476
rect 580404 401474 581004 401476
rect 587160 401474 587760 401476
rect -1996 398476 -1396 398478
rect 804 398476 1404 398478
rect 36804 398476 37404 398478
rect 72804 398476 73404 398478
rect 108804 398476 109404 398478
rect 144804 398476 145404 398478
rect 180804 398476 181404 398478
rect 216804 398476 217404 398478
rect 252804 398476 253404 398478
rect 288804 398476 289404 398478
rect 324804 398476 325404 398478
rect 360804 398476 361404 398478
rect 396804 398476 397404 398478
rect 432804 398476 433404 398478
rect 468804 398476 469404 398478
rect 504804 398476 505404 398478
rect 540804 398476 541404 398478
rect 576804 398476 577404 398478
rect 585320 398476 585920 398478
rect -2916 398454 586840 398476
rect -2916 398218 -1814 398454
rect -1578 398218 986 398454
rect 1222 398218 36986 398454
rect 37222 398218 72986 398454
rect 73222 398218 108986 398454
rect 109222 398218 144986 398454
rect 145222 398218 180986 398454
rect 181222 398218 216986 398454
rect 217222 398218 252986 398454
rect 253222 398218 288986 398454
rect 289222 398218 324986 398454
rect 325222 398218 360986 398454
rect 361222 398218 396986 398454
rect 397222 398218 432986 398454
rect 433222 398218 468986 398454
rect 469222 398218 504986 398454
rect 505222 398218 540986 398454
rect 541222 398218 576986 398454
rect 577222 398218 585502 398454
rect 585738 398218 586840 398454
rect -2916 398134 586840 398218
rect -2916 397898 -1814 398134
rect -1578 397898 986 398134
rect 1222 397898 36986 398134
rect 37222 397898 72986 398134
rect 73222 397898 108986 398134
rect 109222 397898 144986 398134
rect 145222 397898 180986 398134
rect 181222 397898 216986 398134
rect 217222 397898 252986 398134
rect 253222 397898 288986 398134
rect 289222 397898 324986 398134
rect 325222 397898 360986 398134
rect 361222 397898 396986 398134
rect 397222 397898 432986 398134
rect 433222 397898 468986 398134
rect 469222 397898 504986 398134
rect 505222 397898 540986 398134
rect 541222 397898 576986 398134
rect 577222 397898 585502 398134
rect 585738 397898 586840 398134
rect -2916 397876 586840 397898
rect -1996 397874 -1396 397876
rect 804 397874 1404 397876
rect 36804 397874 37404 397876
rect 72804 397874 73404 397876
rect 108804 397874 109404 397876
rect 144804 397874 145404 397876
rect 180804 397874 181404 397876
rect 216804 397874 217404 397876
rect 252804 397874 253404 397876
rect 288804 397874 289404 397876
rect 324804 397874 325404 397876
rect 360804 397874 361404 397876
rect 396804 397874 397404 397876
rect 432804 397874 433404 397876
rect 468804 397874 469404 397876
rect 504804 397874 505404 397876
rect 540804 397874 541404 397876
rect 576804 397874 577404 397876
rect 585320 397874 585920 397876
rect -8436 391276 -7836 391278
rect 29604 391276 30204 391278
rect 65604 391276 66204 391278
rect 101604 391276 102204 391278
rect 137604 391276 138204 391278
rect 173604 391276 174204 391278
rect 209604 391276 210204 391278
rect 245604 391276 246204 391278
rect 281604 391276 282204 391278
rect 317604 391276 318204 391278
rect 353604 391276 354204 391278
rect 389604 391276 390204 391278
rect 425604 391276 426204 391278
rect 461604 391276 462204 391278
rect 497604 391276 498204 391278
rect 533604 391276 534204 391278
rect 569604 391276 570204 391278
rect 591760 391276 592360 391278
rect -8436 391254 592360 391276
rect -8436 391018 -8254 391254
rect -8018 391018 29786 391254
rect 30022 391018 65786 391254
rect 66022 391018 101786 391254
rect 102022 391018 137786 391254
rect 138022 391018 173786 391254
rect 174022 391018 209786 391254
rect 210022 391018 245786 391254
rect 246022 391018 281786 391254
rect 282022 391018 317786 391254
rect 318022 391018 353786 391254
rect 354022 391018 389786 391254
rect 390022 391018 425786 391254
rect 426022 391018 461786 391254
rect 462022 391018 497786 391254
rect 498022 391018 533786 391254
rect 534022 391018 569786 391254
rect 570022 391018 591942 391254
rect 592178 391018 592360 391254
rect -8436 390934 592360 391018
rect -8436 390698 -8254 390934
rect -8018 390698 29786 390934
rect 30022 390698 65786 390934
rect 66022 390698 101786 390934
rect 102022 390698 137786 390934
rect 138022 390698 173786 390934
rect 174022 390698 209786 390934
rect 210022 390698 245786 390934
rect 246022 390698 281786 390934
rect 282022 390698 317786 390934
rect 318022 390698 353786 390934
rect 354022 390698 389786 390934
rect 390022 390698 425786 390934
rect 426022 390698 461786 390934
rect 462022 390698 497786 390934
rect 498022 390698 533786 390934
rect 534022 390698 569786 390934
rect 570022 390698 591942 390934
rect 592178 390698 592360 390934
rect -8436 390676 592360 390698
rect -8436 390674 -7836 390676
rect 29604 390674 30204 390676
rect 65604 390674 66204 390676
rect 101604 390674 102204 390676
rect 137604 390674 138204 390676
rect 173604 390674 174204 390676
rect 209604 390674 210204 390676
rect 245604 390674 246204 390676
rect 281604 390674 282204 390676
rect 317604 390674 318204 390676
rect 353604 390674 354204 390676
rect 389604 390674 390204 390676
rect 425604 390674 426204 390676
rect 461604 390674 462204 390676
rect 497604 390674 498204 390676
rect 533604 390674 534204 390676
rect 569604 390674 570204 390676
rect 591760 390674 592360 390676
rect -6596 387676 -5996 387678
rect 26004 387676 26604 387678
rect 62004 387676 62604 387678
rect 98004 387676 98604 387678
rect 134004 387676 134604 387678
rect 170004 387676 170604 387678
rect 206004 387676 206604 387678
rect 242004 387676 242604 387678
rect 278004 387676 278604 387678
rect 314004 387676 314604 387678
rect 350004 387676 350604 387678
rect 386004 387676 386604 387678
rect 422004 387676 422604 387678
rect 458004 387676 458604 387678
rect 494004 387676 494604 387678
rect 530004 387676 530604 387678
rect 566004 387676 566604 387678
rect 589920 387676 590520 387678
rect -6596 387654 590520 387676
rect -6596 387418 -6414 387654
rect -6178 387418 26186 387654
rect 26422 387418 62186 387654
rect 62422 387418 98186 387654
rect 98422 387418 134186 387654
rect 134422 387418 170186 387654
rect 170422 387418 206186 387654
rect 206422 387418 242186 387654
rect 242422 387418 278186 387654
rect 278422 387418 314186 387654
rect 314422 387418 350186 387654
rect 350422 387418 386186 387654
rect 386422 387418 422186 387654
rect 422422 387418 458186 387654
rect 458422 387418 494186 387654
rect 494422 387418 530186 387654
rect 530422 387418 566186 387654
rect 566422 387418 590102 387654
rect 590338 387418 590520 387654
rect -6596 387334 590520 387418
rect -6596 387098 -6414 387334
rect -6178 387098 26186 387334
rect 26422 387098 62186 387334
rect 62422 387098 98186 387334
rect 98422 387098 134186 387334
rect 134422 387098 170186 387334
rect 170422 387098 206186 387334
rect 206422 387098 242186 387334
rect 242422 387098 278186 387334
rect 278422 387098 314186 387334
rect 314422 387098 350186 387334
rect 350422 387098 386186 387334
rect 386422 387098 422186 387334
rect 422422 387098 458186 387334
rect 458422 387098 494186 387334
rect 494422 387098 530186 387334
rect 530422 387098 566186 387334
rect 566422 387098 590102 387334
rect 590338 387098 590520 387334
rect -6596 387076 590520 387098
rect -6596 387074 -5996 387076
rect 26004 387074 26604 387076
rect 62004 387074 62604 387076
rect 98004 387074 98604 387076
rect 134004 387074 134604 387076
rect 170004 387074 170604 387076
rect 206004 387074 206604 387076
rect 242004 387074 242604 387076
rect 278004 387074 278604 387076
rect 314004 387074 314604 387076
rect 350004 387074 350604 387076
rect 386004 387074 386604 387076
rect 422004 387074 422604 387076
rect 458004 387074 458604 387076
rect 494004 387074 494604 387076
rect 530004 387074 530604 387076
rect 566004 387074 566604 387076
rect 589920 387074 590520 387076
rect -4756 384076 -4156 384078
rect 22404 384076 23004 384078
rect 58404 384076 59004 384078
rect 94404 384076 95004 384078
rect 130404 384076 131004 384078
rect 166404 384076 167004 384078
rect 202404 384076 203004 384078
rect 238404 384076 239004 384078
rect 274404 384076 275004 384078
rect 310404 384076 311004 384078
rect 346404 384076 347004 384078
rect 382404 384076 383004 384078
rect 418404 384076 419004 384078
rect 454404 384076 455004 384078
rect 490404 384076 491004 384078
rect 526404 384076 527004 384078
rect 562404 384076 563004 384078
rect 588080 384076 588680 384078
rect -4756 384054 588680 384076
rect -4756 383818 -4574 384054
rect -4338 383818 22586 384054
rect 22822 383818 58586 384054
rect 58822 383818 94586 384054
rect 94822 383818 130586 384054
rect 130822 383818 166586 384054
rect 166822 383818 202586 384054
rect 202822 383818 238586 384054
rect 238822 383818 274586 384054
rect 274822 383818 310586 384054
rect 310822 383818 346586 384054
rect 346822 383818 382586 384054
rect 382822 383818 418586 384054
rect 418822 383818 454586 384054
rect 454822 383818 490586 384054
rect 490822 383818 526586 384054
rect 526822 383818 562586 384054
rect 562822 383818 588262 384054
rect 588498 383818 588680 384054
rect -4756 383734 588680 383818
rect -4756 383498 -4574 383734
rect -4338 383498 22586 383734
rect 22822 383498 58586 383734
rect 58822 383498 94586 383734
rect 94822 383498 130586 383734
rect 130822 383498 166586 383734
rect 166822 383498 202586 383734
rect 202822 383498 238586 383734
rect 238822 383498 274586 383734
rect 274822 383498 310586 383734
rect 310822 383498 346586 383734
rect 346822 383498 382586 383734
rect 382822 383498 418586 383734
rect 418822 383498 454586 383734
rect 454822 383498 490586 383734
rect 490822 383498 526586 383734
rect 526822 383498 562586 383734
rect 562822 383498 588262 383734
rect 588498 383498 588680 383734
rect -4756 383476 588680 383498
rect -4756 383474 -4156 383476
rect 22404 383474 23004 383476
rect 58404 383474 59004 383476
rect 94404 383474 95004 383476
rect 130404 383474 131004 383476
rect 166404 383474 167004 383476
rect 202404 383474 203004 383476
rect 238404 383474 239004 383476
rect 274404 383474 275004 383476
rect 310404 383474 311004 383476
rect 346404 383474 347004 383476
rect 382404 383474 383004 383476
rect 418404 383474 419004 383476
rect 454404 383474 455004 383476
rect 490404 383474 491004 383476
rect 526404 383474 527004 383476
rect 562404 383474 563004 383476
rect 588080 383474 588680 383476
rect -2916 380476 -2316 380478
rect 18804 380476 19404 380478
rect 54804 380476 55404 380478
rect 90804 380476 91404 380478
rect 126804 380476 127404 380478
rect 162804 380476 163404 380478
rect 198804 380476 199404 380478
rect 234804 380476 235404 380478
rect 270804 380476 271404 380478
rect 306804 380476 307404 380478
rect 342804 380476 343404 380478
rect 378804 380476 379404 380478
rect 414804 380476 415404 380478
rect 450804 380476 451404 380478
rect 486804 380476 487404 380478
rect 522804 380476 523404 380478
rect 558804 380476 559404 380478
rect 586240 380476 586840 380478
rect -2916 380454 586840 380476
rect -2916 380218 -2734 380454
rect -2498 380218 18986 380454
rect 19222 380218 54986 380454
rect 55222 380218 90986 380454
rect 91222 380218 126986 380454
rect 127222 380218 162986 380454
rect 163222 380218 198986 380454
rect 199222 380218 234986 380454
rect 235222 380218 270986 380454
rect 271222 380218 306986 380454
rect 307222 380218 342986 380454
rect 343222 380218 378986 380454
rect 379222 380218 414986 380454
rect 415222 380218 450986 380454
rect 451222 380218 486986 380454
rect 487222 380218 522986 380454
rect 523222 380218 558986 380454
rect 559222 380218 586422 380454
rect 586658 380218 586840 380454
rect -2916 380134 586840 380218
rect -2916 379898 -2734 380134
rect -2498 379898 18986 380134
rect 19222 379898 54986 380134
rect 55222 379898 90986 380134
rect 91222 379898 126986 380134
rect 127222 379898 162986 380134
rect 163222 379898 198986 380134
rect 199222 379898 234986 380134
rect 235222 379898 270986 380134
rect 271222 379898 306986 380134
rect 307222 379898 342986 380134
rect 343222 379898 378986 380134
rect 379222 379898 414986 380134
rect 415222 379898 450986 380134
rect 451222 379898 486986 380134
rect 487222 379898 522986 380134
rect 523222 379898 558986 380134
rect 559222 379898 586422 380134
rect 586658 379898 586840 380134
rect -2916 379876 586840 379898
rect -2916 379874 -2316 379876
rect 18804 379874 19404 379876
rect 54804 379874 55404 379876
rect 90804 379874 91404 379876
rect 126804 379874 127404 379876
rect 162804 379874 163404 379876
rect 198804 379874 199404 379876
rect 234804 379874 235404 379876
rect 270804 379874 271404 379876
rect 306804 379874 307404 379876
rect 342804 379874 343404 379876
rect 378804 379874 379404 379876
rect 414804 379874 415404 379876
rect 450804 379874 451404 379876
rect 486804 379874 487404 379876
rect 522804 379874 523404 379876
rect 558804 379874 559404 379876
rect 586240 379874 586840 379876
rect -7516 373276 -6916 373278
rect 11604 373276 12204 373278
rect 47604 373276 48204 373278
rect 83604 373276 84204 373278
rect 119604 373276 120204 373278
rect 155604 373276 156204 373278
rect 191604 373276 192204 373278
rect 227604 373276 228204 373278
rect 263604 373276 264204 373278
rect 299604 373276 300204 373278
rect 335604 373276 336204 373278
rect 371604 373276 372204 373278
rect 407604 373276 408204 373278
rect 443604 373276 444204 373278
rect 479604 373276 480204 373278
rect 515604 373276 516204 373278
rect 551604 373276 552204 373278
rect 590840 373276 591440 373278
rect -8436 373254 592360 373276
rect -8436 373018 -7334 373254
rect -7098 373018 11786 373254
rect 12022 373018 47786 373254
rect 48022 373018 83786 373254
rect 84022 373018 119786 373254
rect 120022 373018 155786 373254
rect 156022 373018 191786 373254
rect 192022 373018 227786 373254
rect 228022 373018 263786 373254
rect 264022 373018 299786 373254
rect 300022 373018 335786 373254
rect 336022 373018 371786 373254
rect 372022 373018 407786 373254
rect 408022 373018 443786 373254
rect 444022 373018 479786 373254
rect 480022 373018 515786 373254
rect 516022 373018 551786 373254
rect 552022 373018 591022 373254
rect 591258 373018 592360 373254
rect -8436 372934 592360 373018
rect -8436 372698 -7334 372934
rect -7098 372698 11786 372934
rect 12022 372698 47786 372934
rect 48022 372698 83786 372934
rect 84022 372698 119786 372934
rect 120022 372698 155786 372934
rect 156022 372698 191786 372934
rect 192022 372698 227786 372934
rect 228022 372698 263786 372934
rect 264022 372698 299786 372934
rect 300022 372698 335786 372934
rect 336022 372698 371786 372934
rect 372022 372698 407786 372934
rect 408022 372698 443786 372934
rect 444022 372698 479786 372934
rect 480022 372698 515786 372934
rect 516022 372698 551786 372934
rect 552022 372698 591022 372934
rect 591258 372698 592360 372934
rect -8436 372676 592360 372698
rect -7516 372674 -6916 372676
rect 11604 372674 12204 372676
rect 47604 372674 48204 372676
rect 83604 372674 84204 372676
rect 119604 372674 120204 372676
rect 155604 372674 156204 372676
rect 191604 372674 192204 372676
rect 227604 372674 228204 372676
rect 263604 372674 264204 372676
rect 299604 372674 300204 372676
rect 335604 372674 336204 372676
rect 371604 372674 372204 372676
rect 407604 372674 408204 372676
rect 443604 372674 444204 372676
rect 479604 372674 480204 372676
rect 515604 372674 516204 372676
rect 551604 372674 552204 372676
rect 590840 372674 591440 372676
rect -5676 369676 -5076 369678
rect 8004 369676 8604 369678
rect 44004 369676 44604 369678
rect 80004 369676 80604 369678
rect 116004 369676 116604 369678
rect 152004 369676 152604 369678
rect 188004 369676 188604 369678
rect 224004 369676 224604 369678
rect 260004 369676 260604 369678
rect 296004 369676 296604 369678
rect 332004 369676 332604 369678
rect 368004 369676 368604 369678
rect 404004 369676 404604 369678
rect 440004 369676 440604 369678
rect 476004 369676 476604 369678
rect 512004 369676 512604 369678
rect 548004 369676 548604 369678
rect 589000 369676 589600 369678
rect -6596 369654 590520 369676
rect -6596 369418 -5494 369654
rect -5258 369418 8186 369654
rect 8422 369418 44186 369654
rect 44422 369418 80186 369654
rect 80422 369418 116186 369654
rect 116422 369418 152186 369654
rect 152422 369418 188186 369654
rect 188422 369418 224186 369654
rect 224422 369418 260186 369654
rect 260422 369418 296186 369654
rect 296422 369418 332186 369654
rect 332422 369418 368186 369654
rect 368422 369418 404186 369654
rect 404422 369418 440186 369654
rect 440422 369418 476186 369654
rect 476422 369418 512186 369654
rect 512422 369418 548186 369654
rect 548422 369418 589182 369654
rect 589418 369418 590520 369654
rect -6596 369334 590520 369418
rect -6596 369098 -5494 369334
rect -5258 369098 8186 369334
rect 8422 369098 44186 369334
rect 44422 369098 80186 369334
rect 80422 369098 116186 369334
rect 116422 369098 152186 369334
rect 152422 369098 188186 369334
rect 188422 369098 224186 369334
rect 224422 369098 260186 369334
rect 260422 369098 296186 369334
rect 296422 369098 332186 369334
rect 332422 369098 368186 369334
rect 368422 369098 404186 369334
rect 404422 369098 440186 369334
rect 440422 369098 476186 369334
rect 476422 369098 512186 369334
rect 512422 369098 548186 369334
rect 548422 369098 589182 369334
rect 589418 369098 590520 369334
rect -6596 369076 590520 369098
rect -5676 369074 -5076 369076
rect 8004 369074 8604 369076
rect 44004 369074 44604 369076
rect 80004 369074 80604 369076
rect 116004 369074 116604 369076
rect 152004 369074 152604 369076
rect 188004 369074 188604 369076
rect 224004 369074 224604 369076
rect 260004 369074 260604 369076
rect 296004 369074 296604 369076
rect 332004 369074 332604 369076
rect 368004 369074 368604 369076
rect 404004 369074 404604 369076
rect 440004 369074 440604 369076
rect 476004 369074 476604 369076
rect 512004 369074 512604 369076
rect 548004 369074 548604 369076
rect 589000 369074 589600 369076
rect -3836 366076 -3236 366078
rect 4404 366076 5004 366078
rect 40404 366076 41004 366078
rect 76404 366076 77004 366078
rect 112404 366076 113004 366078
rect 148404 366076 149004 366078
rect 184404 366076 185004 366078
rect 220404 366076 221004 366078
rect 256404 366076 257004 366078
rect 292404 366076 293004 366078
rect 328404 366076 329004 366078
rect 364404 366076 365004 366078
rect 400404 366076 401004 366078
rect 436404 366076 437004 366078
rect 472404 366076 473004 366078
rect 508404 366076 509004 366078
rect 544404 366076 545004 366078
rect 580404 366076 581004 366078
rect 587160 366076 587760 366078
rect -4756 366054 588680 366076
rect -4756 365818 -3654 366054
rect -3418 365818 4586 366054
rect 4822 365818 40586 366054
rect 40822 365818 76586 366054
rect 76822 365818 112586 366054
rect 112822 365818 148586 366054
rect 148822 365818 184586 366054
rect 184822 365818 220586 366054
rect 220822 365818 256586 366054
rect 256822 365818 292586 366054
rect 292822 365818 328586 366054
rect 328822 365818 364586 366054
rect 364822 365818 400586 366054
rect 400822 365818 436586 366054
rect 436822 365818 472586 366054
rect 472822 365818 508586 366054
rect 508822 365818 544586 366054
rect 544822 365818 580586 366054
rect 580822 365818 587342 366054
rect 587578 365818 588680 366054
rect -4756 365734 588680 365818
rect -4756 365498 -3654 365734
rect -3418 365498 4586 365734
rect 4822 365498 40586 365734
rect 40822 365498 76586 365734
rect 76822 365498 112586 365734
rect 112822 365498 148586 365734
rect 148822 365498 184586 365734
rect 184822 365498 220586 365734
rect 220822 365498 256586 365734
rect 256822 365498 292586 365734
rect 292822 365498 328586 365734
rect 328822 365498 364586 365734
rect 364822 365498 400586 365734
rect 400822 365498 436586 365734
rect 436822 365498 472586 365734
rect 472822 365498 508586 365734
rect 508822 365498 544586 365734
rect 544822 365498 580586 365734
rect 580822 365498 587342 365734
rect 587578 365498 588680 365734
rect -4756 365476 588680 365498
rect -3836 365474 -3236 365476
rect 4404 365474 5004 365476
rect 40404 365474 41004 365476
rect 76404 365474 77004 365476
rect 112404 365474 113004 365476
rect 148404 365474 149004 365476
rect 184404 365474 185004 365476
rect 220404 365474 221004 365476
rect 256404 365474 257004 365476
rect 292404 365474 293004 365476
rect 328404 365474 329004 365476
rect 364404 365474 365004 365476
rect 400404 365474 401004 365476
rect 436404 365474 437004 365476
rect 472404 365474 473004 365476
rect 508404 365474 509004 365476
rect 544404 365474 545004 365476
rect 580404 365474 581004 365476
rect 587160 365474 587760 365476
rect -1996 362476 -1396 362478
rect 804 362476 1404 362478
rect 36804 362476 37404 362478
rect 72804 362476 73404 362478
rect 108804 362476 109404 362478
rect 144804 362476 145404 362478
rect 180804 362476 181404 362478
rect 216804 362476 217404 362478
rect 252804 362476 253404 362478
rect 288804 362476 289404 362478
rect 324804 362476 325404 362478
rect 360804 362476 361404 362478
rect 396804 362476 397404 362478
rect 432804 362476 433404 362478
rect 468804 362476 469404 362478
rect 504804 362476 505404 362478
rect 540804 362476 541404 362478
rect 576804 362476 577404 362478
rect 585320 362476 585920 362478
rect -2916 362454 586840 362476
rect -2916 362218 -1814 362454
rect -1578 362218 986 362454
rect 1222 362218 36986 362454
rect 37222 362218 72986 362454
rect 73222 362218 108986 362454
rect 109222 362218 144986 362454
rect 145222 362218 180986 362454
rect 181222 362218 216986 362454
rect 217222 362218 252986 362454
rect 253222 362218 288986 362454
rect 289222 362218 324986 362454
rect 325222 362218 360986 362454
rect 361222 362218 396986 362454
rect 397222 362218 432986 362454
rect 433222 362218 468986 362454
rect 469222 362218 504986 362454
rect 505222 362218 540986 362454
rect 541222 362218 576986 362454
rect 577222 362218 585502 362454
rect 585738 362218 586840 362454
rect -2916 362134 586840 362218
rect -2916 361898 -1814 362134
rect -1578 361898 986 362134
rect 1222 361898 36986 362134
rect 37222 361898 72986 362134
rect 73222 361898 108986 362134
rect 109222 361898 144986 362134
rect 145222 361898 180986 362134
rect 181222 361898 216986 362134
rect 217222 361898 252986 362134
rect 253222 361898 288986 362134
rect 289222 361898 324986 362134
rect 325222 361898 360986 362134
rect 361222 361898 396986 362134
rect 397222 361898 432986 362134
rect 433222 361898 468986 362134
rect 469222 361898 504986 362134
rect 505222 361898 540986 362134
rect 541222 361898 576986 362134
rect 577222 361898 585502 362134
rect 585738 361898 586840 362134
rect -2916 361876 586840 361898
rect -1996 361874 -1396 361876
rect 804 361874 1404 361876
rect 36804 361874 37404 361876
rect 72804 361874 73404 361876
rect 108804 361874 109404 361876
rect 144804 361874 145404 361876
rect 180804 361874 181404 361876
rect 216804 361874 217404 361876
rect 252804 361874 253404 361876
rect 288804 361874 289404 361876
rect 324804 361874 325404 361876
rect 360804 361874 361404 361876
rect 396804 361874 397404 361876
rect 432804 361874 433404 361876
rect 468804 361874 469404 361876
rect 504804 361874 505404 361876
rect 540804 361874 541404 361876
rect 576804 361874 577404 361876
rect 585320 361874 585920 361876
rect -8436 355276 -7836 355278
rect 29604 355276 30204 355278
rect 65604 355276 66204 355278
rect 101604 355276 102204 355278
rect 137604 355276 138204 355278
rect 173604 355276 174204 355278
rect 209604 355276 210204 355278
rect 245604 355276 246204 355278
rect 281604 355276 282204 355278
rect 317604 355276 318204 355278
rect 353604 355276 354204 355278
rect 389604 355276 390204 355278
rect 425604 355276 426204 355278
rect 461604 355276 462204 355278
rect 497604 355276 498204 355278
rect 533604 355276 534204 355278
rect 569604 355276 570204 355278
rect 591760 355276 592360 355278
rect -8436 355254 592360 355276
rect -8436 355018 -8254 355254
rect -8018 355018 29786 355254
rect 30022 355018 65786 355254
rect 66022 355018 101786 355254
rect 102022 355018 137786 355254
rect 138022 355018 173786 355254
rect 174022 355018 209786 355254
rect 210022 355018 245786 355254
rect 246022 355018 281786 355254
rect 282022 355018 317786 355254
rect 318022 355018 353786 355254
rect 354022 355018 389786 355254
rect 390022 355018 425786 355254
rect 426022 355018 461786 355254
rect 462022 355018 497786 355254
rect 498022 355018 533786 355254
rect 534022 355018 569786 355254
rect 570022 355018 591942 355254
rect 592178 355018 592360 355254
rect -8436 354934 592360 355018
rect -8436 354698 -8254 354934
rect -8018 354698 29786 354934
rect 30022 354698 65786 354934
rect 66022 354698 101786 354934
rect 102022 354698 137786 354934
rect 138022 354698 173786 354934
rect 174022 354698 209786 354934
rect 210022 354698 245786 354934
rect 246022 354698 281786 354934
rect 282022 354698 317786 354934
rect 318022 354698 353786 354934
rect 354022 354698 389786 354934
rect 390022 354698 425786 354934
rect 426022 354698 461786 354934
rect 462022 354698 497786 354934
rect 498022 354698 533786 354934
rect 534022 354698 569786 354934
rect 570022 354698 591942 354934
rect 592178 354698 592360 354934
rect -8436 354676 592360 354698
rect -8436 354674 -7836 354676
rect 29604 354674 30204 354676
rect 65604 354674 66204 354676
rect 101604 354674 102204 354676
rect 137604 354674 138204 354676
rect 173604 354674 174204 354676
rect 209604 354674 210204 354676
rect 245604 354674 246204 354676
rect 281604 354674 282204 354676
rect 317604 354674 318204 354676
rect 353604 354674 354204 354676
rect 389604 354674 390204 354676
rect 425604 354674 426204 354676
rect 461604 354674 462204 354676
rect 497604 354674 498204 354676
rect 533604 354674 534204 354676
rect 569604 354674 570204 354676
rect 591760 354674 592360 354676
rect -6596 351676 -5996 351678
rect 26004 351676 26604 351678
rect 62004 351676 62604 351678
rect 98004 351676 98604 351678
rect 134004 351676 134604 351678
rect 170004 351676 170604 351678
rect 206004 351676 206604 351678
rect 242004 351676 242604 351678
rect 278004 351676 278604 351678
rect 314004 351676 314604 351678
rect 350004 351676 350604 351678
rect 386004 351676 386604 351678
rect 422004 351676 422604 351678
rect 458004 351676 458604 351678
rect 494004 351676 494604 351678
rect 530004 351676 530604 351678
rect 566004 351676 566604 351678
rect 589920 351676 590520 351678
rect -6596 351654 590520 351676
rect -6596 351418 -6414 351654
rect -6178 351418 26186 351654
rect 26422 351418 62186 351654
rect 62422 351418 98186 351654
rect 98422 351418 134186 351654
rect 134422 351418 170186 351654
rect 170422 351418 206186 351654
rect 206422 351418 242186 351654
rect 242422 351418 278186 351654
rect 278422 351418 314186 351654
rect 314422 351418 350186 351654
rect 350422 351418 386186 351654
rect 386422 351418 422186 351654
rect 422422 351418 458186 351654
rect 458422 351418 494186 351654
rect 494422 351418 530186 351654
rect 530422 351418 566186 351654
rect 566422 351418 590102 351654
rect 590338 351418 590520 351654
rect -6596 351334 590520 351418
rect -6596 351098 -6414 351334
rect -6178 351098 26186 351334
rect 26422 351098 62186 351334
rect 62422 351098 98186 351334
rect 98422 351098 134186 351334
rect 134422 351098 170186 351334
rect 170422 351098 206186 351334
rect 206422 351098 242186 351334
rect 242422 351098 278186 351334
rect 278422 351098 314186 351334
rect 314422 351098 350186 351334
rect 350422 351098 386186 351334
rect 386422 351098 422186 351334
rect 422422 351098 458186 351334
rect 458422 351098 494186 351334
rect 494422 351098 530186 351334
rect 530422 351098 566186 351334
rect 566422 351098 590102 351334
rect 590338 351098 590520 351334
rect -6596 351076 590520 351098
rect -6596 351074 -5996 351076
rect 26004 351074 26604 351076
rect 62004 351074 62604 351076
rect 98004 351074 98604 351076
rect 134004 351074 134604 351076
rect 170004 351074 170604 351076
rect 206004 351074 206604 351076
rect 242004 351074 242604 351076
rect 278004 351074 278604 351076
rect 314004 351074 314604 351076
rect 350004 351074 350604 351076
rect 386004 351074 386604 351076
rect 422004 351074 422604 351076
rect 458004 351074 458604 351076
rect 494004 351074 494604 351076
rect 530004 351074 530604 351076
rect 566004 351074 566604 351076
rect 589920 351074 590520 351076
rect -4756 348076 -4156 348078
rect 22404 348076 23004 348078
rect 58404 348076 59004 348078
rect 94404 348076 95004 348078
rect 130404 348076 131004 348078
rect 166404 348076 167004 348078
rect 202404 348076 203004 348078
rect 238404 348076 239004 348078
rect 274404 348076 275004 348078
rect 310404 348076 311004 348078
rect 346404 348076 347004 348078
rect 382404 348076 383004 348078
rect 418404 348076 419004 348078
rect 454404 348076 455004 348078
rect 490404 348076 491004 348078
rect 526404 348076 527004 348078
rect 562404 348076 563004 348078
rect 588080 348076 588680 348078
rect -4756 348054 588680 348076
rect -4756 347818 -4574 348054
rect -4338 347818 22586 348054
rect 22822 347818 58586 348054
rect 58822 347818 94586 348054
rect 94822 347818 130586 348054
rect 130822 347818 166586 348054
rect 166822 347818 202586 348054
rect 202822 347818 238586 348054
rect 238822 347818 274586 348054
rect 274822 347818 310586 348054
rect 310822 347818 346586 348054
rect 346822 347818 382586 348054
rect 382822 347818 418586 348054
rect 418822 347818 454586 348054
rect 454822 347818 490586 348054
rect 490822 347818 526586 348054
rect 526822 347818 562586 348054
rect 562822 347818 588262 348054
rect 588498 347818 588680 348054
rect -4756 347734 588680 347818
rect -4756 347498 -4574 347734
rect -4338 347498 22586 347734
rect 22822 347498 58586 347734
rect 58822 347498 94586 347734
rect 94822 347498 130586 347734
rect 130822 347498 166586 347734
rect 166822 347498 202586 347734
rect 202822 347498 238586 347734
rect 238822 347498 274586 347734
rect 274822 347498 310586 347734
rect 310822 347498 346586 347734
rect 346822 347498 382586 347734
rect 382822 347498 418586 347734
rect 418822 347498 454586 347734
rect 454822 347498 490586 347734
rect 490822 347498 526586 347734
rect 526822 347498 562586 347734
rect 562822 347498 588262 347734
rect 588498 347498 588680 347734
rect -4756 347476 588680 347498
rect -4756 347474 -4156 347476
rect 22404 347474 23004 347476
rect 58404 347474 59004 347476
rect 94404 347474 95004 347476
rect 130404 347474 131004 347476
rect 166404 347474 167004 347476
rect 202404 347474 203004 347476
rect 238404 347474 239004 347476
rect 274404 347474 275004 347476
rect 310404 347474 311004 347476
rect 346404 347474 347004 347476
rect 382404 347474 383004 347476
rect 418404 347474 419004 347476
rect 454404 347474 455004 347476
rect 490404 347474 491004 347476
rect 526404 347474 527004 347476
rect 562404 347474 563004 347476
rect 588080 347474 588680 347476
rect -2916 344476 -2316 344478
rect 18804 344476 19404 344478
rect 54804 344476 55404 344478
rect 90804 344476 91404 344478
rect 126804 344476 127404 344478
rect 162804 344476 163404 344478
rect 198804 344476 199404 344478
rect 234804 344476 235404 344478
rect 270804 344476 271404 344478
rect 306804 344476 307404 344478
rect 342804 344476 343404 344478
rect 378804 344476 379404 344478
rect 414804 344476 415404 344478
rect 450804 344476 451404 344478
rect 486804 344476 487404 344478
rect 522804 344476 523404 344478
rect 558804 344476 559404 344478
rect 586240 344476 586840 344478
rect -2916 344454 586840 344476
rect -2916 344218 -2734 344454
rect -2498 344218 18986 344454
rect 19222 344218 54986 344454
rect 55222 344218 90986 344454
rect 91222 344218 126986 344454
rect 127222 344218 162986 344454
rect 163222 344218 198986 344454
rect 199222 344218 234986 344454
rect 235222 344218 270986 344454
rect 271222 344218 306986 344454
rect 307222 344218 342986 344454
rect 343222 344218 378986 344454
rect 379222 344218 414986 344454
rect 415222 344218 450986 344454
rect 451222 344218 486986 344454
rect 487222 344218 522986 344454
rect 523222 344218 558986 344454
rect 559222 344218 586422 344454
rect 586658 344218 586840 344454
rect -2916 344134 586840 344218
rect -2916 343898 -2734 344134
rect -2498 343898 18986 344134
rect 19222 343898 54986 344134
rect 55222 343898 90986 344134
rect 91222 343898 126986 344134
rect 127222 343898 162986 344134
rect 163222 343898 198986 344134
rect 199222 343898 234986 344134
rect 235222 343898 270986 344134
rect 271222 343898 306986 344134
rect 307222 343898 342986 344134
rect 343222 343898 378986 344134
rect 379222 343898 414986 344134
rect 415222 343898 450986 344134
rect 451222 343898 486986 344134
rect 487222 343898 522986 344134
rect 523222 343898 558986 344134
rect 559222 343898 586422 344134
rect 586658 343898 586840 344134
rect -2916 343876 586840 343898
rect -2916 343874 -2316 343876
rect 18804 343874 19404 343876
rect 54804 343874 55404 343876
rect 90804 343874 91404 343876
rect 126804 343874 127404 343876
rect 162804 343874 163404 343876
rect 198804 343874 199404 343876
rect 234804 343874 235404 343876
rect 270804 343874 271404 343876
rect 306804 343874 307404 343876
rect 342804 343874 343404 343876
rect 378804 343874 379404 343876
rect 414804 343874 415404 343876
rect 450804 343874 451404 343876
rect 486804 343874 487404 343876
rect 522804 343874 523404 343876
rect 558804 343874 559404 343876
rect 586240 343874 586840 343876
rect -7516 337276 -6916 337278
rect 11604 337276 12204 337278
rect 47604 337276 48204 337278
rect 83604 337276 84204 337278
rect 119604 337276 120204 337278
rect 155604 337276 156204 337278
rect 191604 337276 192204 337278
rect 227604 337276 228204 337278
rect 263604 337276 264204 337278
rect 299604 337276 300204 337278
rect 335604 337276 336204 337278
rect 371604 337276 372204 337278
rect 407604 337276 408204 337278
rect 443604 337276 444204 337278
rect 479604 337276 480204 337278
rect 515604 337276 516204 337278
rect 551604 337276 552204 337278
rect 590840 337276 591440 337278
rect -8436 337254 592360 337276
rect -8436 337018 -7334 337254
rect -7098 337018 11786 337254
rect 12022 337018 47786 337254
rect 48022 337018 83786 337254
rect 84022 337018 119786 337254
rect 120022 337018 155786 337254
rect 156022 337018 191786 337254
rect 192022 337018 227786 337254
rect 228022 337018 263786 337254
rect 264022 337018 299786 337254
rect 300022 337018 335786 337254
rect 336022 337018 371786 337254
rect 372022 337018 407786 337254
rect 408022 337018 443786 337254
rect 444022 337018 479786 337254
rect 480022 337018 515786 337254
rect 516022 337018 551786 337254
rect 552022 337018 591022 337254
rect 591258 337018 592360 337254
rect -8436 336934 592360 337018
rect -8436 336698 -7334 336934
rect -7098 336698 11786 336934
rect 12022 336698 47786 336934
rect 48022 336698 83786 336934
rect 84022 336698 119786 336934
rect 120022 336698 155786 336934
rect 156022 336698 191786 336934
rect 192022 336698 227786 336934
rect 228022 336698 263786 336934
rect 264022 336698 299786 336934
rect 300022 336698 335786 336934
rect 336022 336698 371786 336934
rect 372022 336698 407786 336934
rect 408022 336698 443786 336934
rect 444022 336698 479786 336934
rect 480022 336698 515786 336934
rect 516022 336698 551786 336934
rect 552022 336698 591022 336934
rect 591258 336698 592360 336934
rect -8436 336676 592360 336698
rect -7516 336674 -6916 336676
rect 11604 336674 12204 336676
rect 47604 336674 48204 336676
rect 83604 336674 84204 336676
rect 119604 336674 120204 336676
rect 155604 336674 156204 336676
rect 191604 336674 192204 336676
rect 227604 336674 228204 336676
rect 263604 336674 264204 336676
rect 299604 336674 300204 336676
rect 335604 336674 336204 336676
rect 371604 336674 372204 336676
rect 407604 336674 408204 336676
rect 443604 336674 444204 336676
rect 479604 336674 480204 336676
rect 515604 336674 516204 336676
rect 551604 336674 552204 336676
rect 590840 336674 591440 336676
rect -5676 333676 -5076 333678
rect 8004 333676 8604 333678
rect 44004 333676 44604 333678
rect 80004 333676 80604 333678
rect 116004 333676 116604 333678
rect 152004 333676 152604 333678
rect 188004 333676 188604 333678
rect 224004 333676 224604 333678
rect 260004 333676 260604 333678
rect 296004 333676 296604 333678
rect 332004 333676 332604 333678
rect 368004 333676 368604 333678
rect 404004 333676 404604 333678
rect 440004 333676 440604 333678
rect 476004 333676 476604 333678
rect 512004 333676 512604 333678
rect 548004 333676 548604 333678
rect 589000 333676 589600 333678
rect -6596 333654 590520 333676
rect -6596 333418 -5494 333654
rect -5258 333418 8186 333654
rect 8422 333418 44186 333654
rect 44422 333418 80186 333654
rect 80422 333418 116186 333654
rect 116422 333418 152186 333654
rect 152422 333418 188186 333654
rect 188422 333418 224186 333654
rect 224422 333418 260186 333654
rect 260422 333418 296186 333654
rect 296422 333418 332186 333654
rect 332422 333418 368186 333654
rect 368422 333418 404186 333654
rect 404422 333418 440186 333654
rect 440422 333418 476186 333654
rect 476422 333418 512186 333654
rect 512422 333418 548186 333654
rect 548422 333418 589182 333654
rect 589418 333418 590520 333654
rect -6596 333334 590520 333418
rect -6596 333098 -5494 333334
rect -5258 333098 8186 333334
rect 8422 333098 44186 333334
rect 44422 333098 80186 333334
rect 80422 333098 116186 333334
rect 116422 333098 152186 333334
rect 152422 333098 188186 333334
rect 188422 333098 224186 333334
rect 224422 333098 260186 333334
rect 260422 333098 296186 333334
rect 296422 333098 332186 333334
rect 332422 333098 368186 333334
rect 368422 333098 404186 333334
rect 404422 333098 440186 333334
rect 440422 333098 476186 333334
rect 476422 333098 512186 333334
rect 512422 333098 548186 333334
rect 548422 333098 589182 333334
rect 589418 333098 590520 333334
rect -6596 333076 590520 333098
rect -5676 333074 -5076 333076
rect 8004 333074 8604 333076
rect 44004 333074 44604 333076
rect 80004 333074 80604 333076
rect 116004 333074 116604 333076
rect 152004 333074 152604 333076
rect 188004 333074 188604 333076
rect 224004 333074 224604 333076
rect 260004 333074 260604 333076
rect 296004 333074 296604 333076
rect 332004 333074 332604 333076
rect 368004 333074 368604 333076
rect 404004 333074 404604 333076
rect 440004 333074 440604 333076
rect 476004 333074 476604 333076
rect 512004 333074 512604 333076
rect 548004 333074 548604 333076
rect 589000 333074 589600 333076
rect -3836 330076 -3236 330078
rect 4404 330076 5004 330078
rect 40404 330076 41004 330078
rect 76404 330076 77004 330078
rect 112404 330076 113004 330078
rect 148404 330076 149004 330078
rect 184404 330076 185004 330078
rect 220404 330076 221004 330078
rect 256404 330076 257004 330078
rect 292404 330076 293004 330078
rect 328404 330076 329004 330078
rect 364404 330076 365004 330078
rect 400404 330076 401004 330078
rect 436404 330076 437004 330078
rect 472404 330076 473004 330078
rect 508404 330076 509004 330078
rect 544404 330076 545004 330078
rect 580404 330076 581004 330078
rect 587160 330076 587760 330078
rect -4756 330054 588680 330076
rect -4756 329818 -3654 330054
rect -3418 329818 4586 330054
rect 4822 329818 40586 330054
rect 40822 329818 76586 330054
rect 76822 329818 112586 330054
rect 112822 329818 148586 330054
rect 148822 329818 184586 330054
rect 184822 329818 220586 330054
rect 220822 329818 256586 330054
rect 256822 329818 292586 330054
rect 292822 329818 328586 330054
rect 328822 329818 364586 330054
rect 364822 329818 400586 330054
rect 400822 329818 436586 330054
rect 436822 329818 472586 330054
rect 472822 329818 508586 330054
rect 508822 329818 544586 330054
rect 544822 329818 580586 330054
rect 580822 329818 587342 330054
rect 587578 329818 588680 330054
rect -4756 329734 588680 329818
rect -4756 329498 -3654 329734
rect -3418 329498 4586 329734
rect 4822 329498 40586 329734
rect 40822 329498 76586 329734
rect 76822 329498 112586 329734
rect 112822 329498 148586 329734
rect 148822 329498 184586 329734
rect 184822 329498 220586 329734
rect 220822 329498 256586 329734
rect 256822 329498 292586 329734
rect 292822 329498 328586 329734
rect 328822 329498 364586 329734
rect 364822 329498 400586 329734
rect 400822 329498 436586 329734
rect 436822 329498 472586 329734
rect 472822 329498 508586 329734
rect 508822 329498 544586 329734
rect 544822 329498 580586 329734
rect 580822 329498 587342 329734
rect 587578 329498 588680 329734
rect -4756 329476 588680 329498
rect -3836 329474 -3236 329476
rect 4404 329474 5004 329476
rect 40404 329474 41004 329476
rect 76404 329474 77004 329476
rect 112404 329474 113004 329476
rect 148404 329474 149004 329476
rect 184404 329474 185004 329476
rect 220404 329474 221004 329476
rect 256404 329474 257004 329476
rect 292404 329474 293004 329476
rect 328404 329474 329004 329476
rect 364404 329474 365004 329476
rect 400404 329474 401004 329476
rect 436404 329474 437004 329476
rect 472404 329474 473004 329476
rect 508404 329474 509004 329476
rect 544404 329474 545004 329476
rect 580404 329474 581004 329476
rect 587160 329474 587760 329476
rect -1996 326476 -1396 326478
rect 804 326476 1404 326478
rect 36804 326476 37404 326478
rect 72804 326476 73404 326478
rect 108804 326476 109404 326478
rect 144804 326476 145404 326478
rect 180804 326476 181404 326478
rect 216804 326476 217404 326478
rect 252804 326476 253404 326478
rect 288804 326476 289404 326478
rect 324804 326476 325404 326478
rect 360804 326476 361404 326478
rect 396804 326476 397404 326478
rect 432804 326476 433404 326478
rect 468804 326476 469404 326478
rect 504804 326476 505404 326478
rect 540804 326476 541404 326478
rect 576804 326476 577404 326478
rect 585320 326476 585920 326478
rect -2916 326454 586840 326476
rect -2916 326218 -1814 326454
rect -1578 326218 986 326454
rect 1222 326218 36986 326454
rect 37222 326218 72986 326454
rect 73222 326218 108986 326454
rect 109222 326218 144986 326454
rect 145222 326218 180986 326454
rect 181222 326218 216986 326454
rect 217222 326218 252986 326454
rect 253222 326218 288986 326454
rect 289222 326218 324986 326454
rect 325222 326218 360986 326454
rect 361222 326218 396986 326454
rect 397222 326218 432986 326454
rect 433222 326218 468986 326454
rect 469222 326218 504986 326454
rect 505222 326218 540986 326454
rect 541222 326218 576986 326454
rect 577222 326218 585502 326454
rect 585738 326218 586840 326454
rect -2916 326134 586840 326218
rect -2916 325898 -1814 326134
rect -1578 325898 986 326134
rect 1222 325898 36986 326134
rect 37222 325898 72986 326134
rect 73222 325898 108986 326134
rect 109222 325898 144986 326134
rect 145222 325898 180986 326134
rect 181222 325898 216986 326134
rect 217222 325898 252986 326134
rect 253222 325898 288986 326134
rect 289222 325898 324986 326134
rect 325222 325898 360986 326134
rect 361222 325898 396986 326134
rect 397222 325898 432986 326134
rect 433222 325898 468986 326134
rect 469222 325898 504986 326134
rect 505222 325898 540986 326134
rect 541222 325898 576986 326134
rect 577222 325898 585502 326134
rect 585738 325898 586840 326134
rect -2916 325876 586840 325898
rect -1996 325874 -1396 325876
rect 804 325874 1404 325876
rect 36804 325874 37404 325876
rect 72804 325874 73404 325876
rect 108804 325874 109404 325876
rect 144804 325874 145404 325876
rect 180804 325874 181404 325876
rect 216804 325874 217404 325876
rect 252804 325874 253404 325876
rect 288804 325874 289404 325876
rect 324804 325874 325404 325876
rect 360804 325874 361404 325876
rect 396804 325874 397404 325876
rect 432804 325874 433404 325876
rect 468804 325874 469404 325876
rect 504804 325874 505404 325876
rect 540804 325874 541404 325876
rect 576804 325874 577404 325876
rect 585320 325874 585920 325876
rect -8436 319276 -7836 319278
rect 29604 319276 30204 319278
rect 65604 319276 66204 319278
rect 101604 319276 102204 319278
rect 137604 319276 138204 319278
rect 173604 319276 174204 319278
rect 209604 319276 210204 319278
rect 245604 319276 246204 319278
rect 281604 319276 282204 319278
rect 317604 319276 318204 319278
rect 353604 319276 354204 319278
rect 389604 319276 390204 319278
rect 425604 319276 426204 319278
rect 461604 319276 462204 319278
rect 497604 319276 498204 319278
rect 533604 319276 534204 319278
rect 569604 319276 570204 319278
rect 591760 319276 592360 319278
rect -8436 319254 592360 319276
rect -8436 319018 -8254 319254
rect -8018 319018 29786 319254
rect 30022 319018 65786 319254
rect 66022 319018 101786 319254
rect 102022 319018 137786 319254
rect 138022 319018 173786 319254
rect 174022 319018 209786 319254
rect 210022 319018 245786 319254
rect 246022 319018 281786 319254
rect 282022 319018 317786 319254
rect 318022 319018 353786 319254
rect 354022 319018 389786 319254
rect 390022 319018 425786 319254
rect 426022 319018 461786 319254
rect 462022 319018 497786 319254
rect 498022 319018 533786 319254
rect 534022 319018 569786 319254
rect 570022 319018 591942 319254
rect 592178 319018 592360 319254
rect -8436 318934 592360 319018
rect -8436 318698 -8254 318934
rect -8018 318698 29786 318934
rect 30022 318698 65786 318934
rect 66022 318698 101786 318934
rect 102022 318698 137786 318934
rect 138022 318698 173786 318934
rect 174022 318698 209786 318934
rect 210022 318698 245786 318934
rect 246022 318698 281786 318934
rect 282022 318698 317786 318934
rect 318022 318698 353786 318934
rect 354022 318698 389786 318934
rect 390022 318698 425786 318934
rect 426022 318698 461786 318934
rect 462022 318698 497786 318934
rect 498022 318698 533786 318934
rect 534022 318698 569786 318934
rect 570022 318698 591942 318934
rect 592178 318698 592360 318934
rect -8436 318676 592360 318698
rect -8436 318674 -7836 318676
rect 29604 318674 30204 318676
rect 65604 318674 66204 318676
rect 101604 318674 102204 318676
rect 137604 318674 138204 318676
rect 173604 318674 174204 318676
rect 209604 318674 210204 318676
rect 245604 318674 246204 318676
rect 281604 318674 282204 318676
rect 317604 318674 318204 318676
rect 353604 318674 354204 318676
rect 389604 318674 390204 318676
rect 425604 318674 426204 318676
rect 461604 318674 462204 318676
rect 497604 318674 498204 318676
rect 533604 318674 534204 318676
rect 569604 318674 570204 318676
rect 591760 318674 592360 318676
rect -6596 315676 -5996 315678
rect 26004 315676 26604 315678
rect 62004 315676 62604 315678
rect 98004 315676 98604 315678
rect 134004 315676 134604 315678
rect 170004 315676 170604 315678
rect 206004 315676 206604 315678
rect 242004 315676 242604 315678
rect 278004 315676 278604 315678
rect 314004 315676 314604 315678
rect 350004 315676 350604 315678
rect 386004 315676 386604 315678
rect 422004 315676 422604 315678
rect 458004 315676 458604 315678
rect 494004 315676 494604 315678
rect 530004 315676 530604 315678
rect 566004 315676 566604 315678
rect 589920 315676 590520 315678
rect -6596 315654 590520 315676
rect -6596 315418 -6414 315654
rect -6178 315418 26186 315654
rect 26422 315418 62186 315654
rect 62422 315418 98186 315654
rect 98422 315418 134186 315654
rect 134422 315418 170186 315654
rect 170422 315418 206186 315654
rect 206422 315418 242186 315654
rect 242422 315418 278186 315654
rect 278422 315418 314186 315654
rect 314422 315418 350186 315654
rect 350422 315418 386186 315654
rect 386422 315418 422186 315654
rect 422422 315418 458186 315654
rect 458422 315418 494186 315654
rect 494422 315418 530186 315654
rect 530422 315418 566186 315654
rect 566422 315418 590102 315654
rect 590338 315418 590520 315654
rect -6596 315334 590520 315418
rect -6596 315098 -6414 315334
rect -6178 315098 26186 315334
rect 26422 315098 62186 315334
rect 62422 315098 98186 315334
rect 98422 315098 134186 315334
rect 134422 315098 170186 315334
rect 170422 315098 206186 315334
rect 206422 315098 242186 315334
rect 242422 315098 278186 315334
rect 278422 315098 314186 315334
rect 314422 315098 350186 315334
rect 350422 315098 386186 315334
rect 386422 315098 422186 315334
rect 422422 315098 458186 315334
rect 458422 315098 494186 315334
rect 494422 315098 530186 315334
rect 530422 315098 566186 315334
rect 566422 315098 590102 315334
rect 590338 315098 590520 315334
rect -6596 315076 590520 315098
rect -6596 315074 -5996 315076
rect 26004 315074 26604 315076
rect 62004 315074 62604 315076
rect 98004 315074 98604 315076
rect 134004 315074 134604 315076
rect 170004 315074 170604 315076
rect 206004 315074 206604 315076
rect 242004 315074 242604 315076
rect 278004 315074 278604 315076
rect 314004 315074 314604 315076
rect 350004 315074 350604 315076
rect 386004 315074 386604 315076
rect 422004 315074 422604 315076
rect 458004 315074 458604 315076
rect 494004 315074 494604 315076
rect 530004 315074 530604 315076
rect 566004 315074 566604 315076
rect 589920 315074 590520 315076
rect -4756 312076 -4156 312078
rect 22404 312076 23004 312078
rect 58404 312076 59004 312078
rect 94404 312076 95004 312078
rect 130404 312076 131004 312078
rect 166404 312076 167004 312078
rect 202404 312076 203004 312078
rect 238404 312076 239004 312078
rect 274404 312076 275004 312078
rect 310404 312076 311004 312078
rect 346404 312076 347004 312078
rect 382404 312076 383004 312078
rect 418404 312076 419004 312078
rect 454404 312076 455004 312078
rect 490404 312076 491004 312078
rect 526404 312076 527004 312078
rect 562404 312076 563004 312078
rect 588080 312076 588680 312078
rect -4756 312054 588680 312076
rect -4756 311818 -4574 312054
rect -4338 311818 22586 312054
rect 22822 311818 58586 312054
rect 58822 311818 94586 312054
rect 94822 311818 130586 312054
rect 130822 311818 166586 312054
rect 166822 311818 202586 312054
rect 202822 311818 238586 312054
rect 238822 311818 274586 312054
rect 274822 311818 310586 312054
rect 310822 311818 346586 312054
rect 346822 311818 382586 312054
rect 382822 311818 418586 312054
rect 418822 311818 454586 312054
rect 454822 311818 490586 312054
rect 490822 311818 526586 312054
rect 526822 311818 562586 312054
rect 562822 311818 588262 312054
rect 588498 311818 588680 312054
rect -4756 311734 588680 311818
rect -4756 311498 -4574 311734
rect -4338 311498 22586 311734
rect 22822 311498 58586 311734
rect 58822 311498 94586 311734
rect 94822 311498 130586 311734
rect 130822 311498 166586 311734
rect 166822 311498 202586 311734
rect 202822 311498 238586 311734
rect 238822 311498 274586 311734
rect 274822 311498 310586 311734
rect 310822 311498 346586 311734
rect 346822 311498 382586 311734
rect 382822 311498 418586 311734
rect 418822 311498 454586 311734
rect 454822 311498 490586 311734
rect 490822 311498 526586 311734
rect 526822 311498 562586 311734
rect 562822 311498 588262 311734
rect 588498 311498 588680 311734
rect -4756 311476 588680 311498
rect -4756 311474 -4156 311476
rect 22404 311474 23004 311476
rect 58404 311474 59004 311476
rect 94404 311474 95004 311476
rect 130404 311474 131004 311476
rect 166404 311474 167004 311476
rect 202404 311474 203004 311476
rect 238404 311474 239004 311476
rect 274404 311474 275004 311476
rect 310404 311474 311004 311476
rect 346404 311474 347004 311476
rect 382404 311474 383004 311476
rect 418404 311474 419004 311476
rect 454404 311474 455004 311476
rect 490404 311474 491004 311476
rect 526404 311474 527004 311476
rect 562404 311474 563004 311476
rect 588080 311474 588680 311476
rect -2916 308476 -2316 308478
rect 18804 308476 19404 308478
rect 54804 308476 55404 308478
rect 90804 308476 91404 308478
rect 126804 308476 127404 308478
rect 162804 308476 163404 308478
rect 198804 308476 199404 308478
rect 234804 308476 235404 308478
rect 270804 308476 271404 308478
rect 306804 308476 307404 308478
rect 342804 308476 343404 308478
rect 378804 308476 379404 308478
rect 414804 308476 415404 308478
rect 450804 308476 451404 308478
rect 486804 308476 487404 308478
rect 522804 308476 523404 308478
rect 558804 308476 559404 308478
rect 586240 308476 586840 308478
rect -2916 308454 586840 308476
rect -2916 308218 -2734 308454
rect -2498 308218 18986 308454
rect 19222 308218 54986 308454
rect 55222 308218 90986 308454
rect 91222 308218 126986 308454
rect 127222 308218 162986 308454
rect 163222 308218 198986 308454
rect 199222 308218 234986 308454
rect 235222 308218 270986 308454
rect 271222 308218 306986 308454
rect 307222 308218 342986 308454
rect 343222 308218 378986 308454
rect 379222 308218 414986 308454
rect 415222 308218 450986 308454
rect 451222 308218 486986 308454
rect 487222 308218 522986 308454
rect 523222 308218 558986 308454
rect 559222 308218 586422 308454
rect 586658 308218 586840 308454
rect -2916 308134 586840 308218
rect -2916 307898 -2734 308134
rect -2498 307898 18986 308134
rect 19222 307898 54986 308134
rect 55222 307898 90986 308134
rect 91222 307898 126986 308134
rect 127222 307898 162986 308134
rect 163222 307898 198986 308134
rect 199222 307898 234986 308134
rect 235222 307898 270986 308134
rect 271222 307898 306986 308134
rect 307222 307898 342986 308134
rect 343222 307898 378986 308134
rect 379222 307898 414986 308134
rect 415222 307898 450986 308134
rect 451222 307898 486986 308134
rect 487222 307898 522986 308134
rect 523222 307898 558986 308134
rect 559222 307898 586422 308134
rect 586658 307898 586840 308134
rect -2916 307876 586840 307898
rect -2916 307874 -2316 307876
rect 18804 307874 19404 307876
rect 54804 307874 55404 307876
rect 90804 307874 91404 307876
rect 126804 307874 127404 307876
rect 162804 307874 163404 307876
rect 198804 307874 199404 307876
rect 234804 307874 235404 307876
rect 270804 307874 271404 307876
rect 306804 307874 307404 307876
rect 342804 307874 343404 307876
rect 378804 307874 379404 307876
rect 414804 307874 415404 307876
rect 450804 307874 451404 307876
rect 486804 307874 487404 307876
rect 522804 307874 523404 307876
rect 558804 307874 559404 307876
rect 586240 307874 586840 307876
rect -7516 301276 -6916 301278
rect 11604 301276 12204 301278
rect 47604 301276 48204 301278
rect 83604 301276 84204 301278
rect 119604 301276 120204 301278
rect 155604 301276 156204 301278
rect 191604 301276 192204 301278
rect 227604 301276 228204 301278
rect 263604 301276 264204 301278
rect 299604 301276 300204 301278
rect 335604 301276 336204 301278
rect 371604 301276 372204 301278
rect 407604 301276 408204 301278
rect 443604 301276 444204 301278
rect 479604 301276 480204 301278
rect 515604 301276 516204 301278
rect 551604 301276 552204 301278
rect 590840 301276 591440 301278
rect -8436 301254 592360 301276
rect -8436 301018 -7334 301254
rect -7098 301018 11786 301254
rect 12022 301018 47786 301254
rect 48022 301018 83786 301254
rect 84022 301018 119786 301254
rect 120022 301018 155786 301254
rect 156022 301018 191786 301254
rect 192022 301018 227786 301254
rect 228022 301018 263786 301254
rect 264022 301018 299786 301254
rect 300022 301018 335786 301254
rect 336022 301018 371786 301254
rect 372022 301018 407786 301254
rect 408022 301018 443786 301254
rect 444022 301018 479786 301254
rect 480022 301018 515786 301254
rect 516022 301018 551786 301254
rect 552022 301018 591022 301254
rect 591258 301018 592360 301254
rect -8436 300934 592360 301018
rect -8436 300698 -7334 300934
rect -7098 300698 11786 300934
rect 12022 300698 47786 300934
rect 48022 300698 83786 300934
rect 84022 300698 119786 300934
rect 120022 300698 155786 300934
rect 156022 300698 191786 300934
rect 192022 300698 227786 300934
rect 228022 300698 263786 300934
rect 264022 300698 299786 300934
rect 300022 300698 335786 300934
rect 336022 300698 371786 300934
rect 372022 300698 407786 300934
rect 408022 300698 443786 300934
rect 444022 300698 479786 300934
rect 480022 300698 515786 300934
rect 516022 300698 551786 300934
rect 552022 300698 591022 300934
rect 591258 300698 592360 300934
rect -8436 300676 592360 300698
rect -7516 300674 -6916 300676
rect 11604 300674 12204 300676
rect 47604 300674 48204 300676
rect 83604 300674 84204 300676
rect 119604 300674 120204 300676
rect 155604 300674 156204 300676
rect 191604 300674 192204 300676
rect 227604 300674 228204 300676
rect 263604 300674 264204 300676
rect 299604 300674 300204 300676
rect 335604 300674 336204 300676
rect 371604 300674 372204 300676
rect 407604 300674 408204 300676
rect 443604 300674 444204 300676
rect 479604 300674 480204 300676
rect 515604 300674 516204 300676
rect 551604 300674 552204 300676
rect 590840 300674 591440 300676
rect -5676 297676 -5076 297678
rect 8004 297676 8604 297678
rect 44004 297676 44604 297678
rect 80004 297676 80604 297678
rect 116004 297676 116604 297678
rect 152004 297676 152604 297678
rect 188004 297676 188604 297678
rect 224004 297676 224604 297678
rect 260004 297676 260604 297678
rect 296004 297676 296604 297678
rect 332004 297676 332604 297678
rect 368004 297676 368604 297678
rect 404004 297676 404604 297678
rect 440004 297676 440604 297678
rect 476004 297676 476604 297678
rect 512004 297676 512604 297678
rect 548004 297676 548604 297678
rect 589000 297676 589600 297678
rect -6596 297654 590520 297676
rect -6596 297418 -5494 297654
rect -5258 297418 8186 297654
rect 8422 297418 44186 297654
rect 44422 297418 80186 297654
rect 80422 297418 116186 297654
rect 116422 297418 152186 297654
rect 152422 297418 188186 297654
rect 188422 297418 224186 297654
rect 224422 297418 260186 297654
rect 260422 297418 296186 297654
rect 296422 297418 332186 297654
rect 332422 297418 368186 297654
rect 368422 297418 404186 297654
rect 404422 297418 440186 297654
rect 440422 297418 476186 297654
rect 476422 297418 512186 297654
rect 512422 297418 548186 297654
rect 548422 297418 589182 297654
rect 589418 297418 590520 297654
rect -6596 297334 590520 297418
rect -6596 297098 -5494 297334
rect -5258 297098 8186 297334
rect 8422 297098 44186 297334
rect 44422 297098 80186 297334
rect 80422 297098 116186 297334
rect 116422 297098 152186 297334
rect 152422 297098 188186 297334
rect 188422 297098 224186 297334
rect 224422 297098 260186 297334
rect 260422 297098 296186 297334
rect 296422 297098 332186 297334
rect 332422 297098 368186 297334
rect 368422 297098 404186 297334
rect 404422 297098 440186 297334
rect 440422 297098 476186 297334
rect 476422 297098 512186 297334
rect 512422 297098 548186 297334
rect 548422 297098 589182 297334
rect 589418 297098 590520 297334
rect -6596 297076 590520 297098
rect -5676 297074 -5076 297076
rect 8004 297074 8604 297076
rect 44004 297074 44604 297076
rect 80004 297074 80604 297076
rect 116004 297074 116604 297076
rect 152004 297074 152604 297076
rect 188004 297074 188604 297076
rect 224004 297074 224604 297076
rect 260004 297074 260604 297076
rect 296004 297074 296604 297076
rect 332004 297074 332604 297076
rect 368004 297074 368604 297076
rect 404004 297074 404604 297076
rect 440004 297074 440604 297076
rect 476004 297074 476604 297076
rect 512004 297074 512604 297076
rect 548004 297074 548604 297076
rect 589000 297074 589600 297076
rect -3836 294076 -3236 294078
rect 4404 294076 5004 294078
rect 40404 294076 41004 294078
rect 76404 294076 77004 294078
rect 112404 294076 113004 294078
rect 148404 294076 149004 294078
rect 184404 294076 185004 294078
rect 220404 294076 221004 294078
rect 256404 294076 257004 294078
rect 292404 294076 293004 294078
rect 328404 294076 329004 294078
rect 364404 294076 365004 294078
rect 400404 294076 401004 294078
rect 436404 294076 437004 294078
rect 472404 294076 473004 294078
rect 508404 294076 509004 294078
rect 544404 294076 545004 294078
rect 580404 294076 581004 294078
rect 587160 294076 587760 294078
rect -4756 294054 588680 294076
rect -4756 293818 -3654 294054
rect -3418 293818 4586 294054
rect 4822 293818 40586 294054
rect 40822 293818 76586 294054
rect 76822 293818 112586 294054
rect 112822 293818 148586 294054
rect 148822 293818 184586 294054
rect 184822 293818 220586 294054
rect 220822 293818 256586 294054
rect 256822 293818 292586 294054
rect 292822 293818 328586 294054
rect 328822 293818 364586 294054
rect 364822 293818 400586 294054
rect 400822 293818 436586 294054
rect 436822 293818 472586 294054
rect 472822 293818 508586 294054
rect 508822 293818 544586 294054
rect 544822 293818 580586 294054
rect 580822 293818 587342 294054
rect 587578 293818 588680 294054
rect -4756 293734 588680 293818
rect -4756 293498 -3654 293734
rect -3418 293498 4586 293734
rect 4822 293498 40586 293734
rect 40822 293498 76586 293734
rect 76822 293498 112586 293734
rect 112822 293498 148586 293734
rect 148822 293498 184586 293734
rect 184822 293498 220586 293734
rect 220822 293498 256586 293734
rect 256822 293498 292586 293734
rect 292822 293498 328586 293734
rect 328822 293498 364586 293734
rect 364822 293498 400586 293734
rect 400822 293498 436586 293734
rect 436822 293498 472586 293734
rect 472822 293498 508586 293734
rect 508822 293498 544586 293734
rect 544822 293498 580586 293734
rect 580822 293498 587342 293734
rect 587578 293498 588680 293734
rect -4756 293476 588680 293498
rect -3836 293474 -3236 293476
rect 4404 293474 5004 293476
rect 40404 293474 41004 293476
rect 76404 293474 77004 293476
rect 112404 293474 113004 293476
rect 148404 293474 149004 293476
rect 184404 293474 185004 293476
rect 220404 293474 221004 293476
rect 256404 293474 257004 293476
rect 292404 293474 293004 293476
rect 328404 293474 329004 293476
rect 364404 293474 365004 293476
rect 400404 293474 401004 293476
rect 436404 293474 437004 293476
rect 472404 293474 473004 293476
rect 508404 293474 509004 293476
rect 544404 293474 545004 293476
rect 580404 293474 581004 293476
rect 587160 293474 587760 293476
rect -1996 290476 -1396 290478
rect 804 290476 1404 290478
rect 36804 290476 37404 290478
rect 72804 290476 73404 290478
rect 108804 290476 109404 290478
rect 144804 290476 145404 290478
rect 180804 290476 181404 290478
rect 216804 290476 217404 290478
rect 252804 290476 253404 290478
rect 288804 290476 289404 290478
rect 324804 290476 325404 290478
rect 360804 290476 361404 290478
rect 396804 290476 397404 290478
rect 432804 290476 433404 290478
rect 468804 290476 469404 290478
rect 504804 290476 505404 290478
rect 540804 290476 541404 290478
rect 576804 290476 577404 290478
rect 585320 290476 585920 290478
rect -2916 290454 586840 290476
rect -2916 290218 -1814 290454
rect -1578 290218 986 290454
rect 1222 290218 36986 290454
rect 37222 290218 72986 290454
rect 73222 290218 108986 290454
rect 109222 290218 144986 290454
rect 145222 290218 180986 290454
rect 181222 290218 216986 290454
rect 217222 290218 252986 290454
rect 253222 290218 288986 290454
rect 289222 290218 324986 290454
rect 325222 290218 360986 290454
rect 361222 290218 396986 290454
rect 397222 290218 432986 290454
rect 433222 290218 468986 290454
rect 469222 290218 504986 290454
rect 505222 290218 540986 290454
rect 541222 290218 576986 290454
rect 577222 290218 585502 290454
rect 585738 290218 586840 290454
rect -2916 290134 586840 290218
rect -2916 289898 -1814 290134
rect -1578 289898 986 290134
rect 1222 289898 36986 290134
rect 37222 289898 72986 290134
rect 73222 289898 108986 290134
rect 109222 289898 144986 290134
rect 145222 289898 180986 290134
rect 181222 289898 216986 290134
rect 217222 289898 252986 290134
rect 253222 289898 288986 290134
rect 289222 289898 324986 290134
rect 325222 289898 360986 290134
rect 361222 289898 396986 290134
rect 397222 289898 432986 290134
rect 433222 289898 468986 290134
rect 469222 289898 504986 290134
rect 505222 289898 540986 290134
rect 541222 289898 576986 290134
rect 577222 289898 585502 290134
rect 585738 289898 586840 290134
rect -2916 289876 586840 289898
rect -1996 289874 -1396 289876
rect 804 289874 1404 289876
rect 36804 289874 37404 289876
rect 72804 289874 73404 289876
rect 108804 289874 109404 289876
rect 144804 289874 145404 289876
rect 180804 289874 181404 289876
rect 216804 289874 217404 289876
rect 252804 289874 253404 289876
rect 288804 289874 289404 289876
rect 324804 289874 325404 289876
rect 360804 289874 361404 289876
rect 396804 289874 397404 289876
rect 432804 289874 433404 289876
rect 468804 289874 469404 289876
rect 504804 289874 505404 289876
rect 540804 289874 541404 289876
rect 576804 289874 577404 289876
rect 585320 289874 585920 289876
rect -8436 283276 -7836 283278
rect 29604 283276 30204 283278
rect 65604 283276 66204 283278
rect 101604 283276 102204 283278
rect 137604 283276 138204 283278
rect 173604 283276 174204 283278
rect 209604 283276 210204 283278
rect 245604 283276 246204 283278
rect 281604 283276 282204 283278
rect 317604 283276 318204 283278
rect 353604 283276 354204 283278
rect 389604 283276 390204 283278
rect 425604 283276 426204 283278
rect 461604 283276 462204 283278
rect 497604 283276 498204 283278
rect 533604 283276 534204 283278
rect 569604 283276 570204 283278
rect 591760 283276 592360 283278
rect -8436 283254 592360 283276
rect -8436 283018 -8254 283254
rect -8018 283018 29786 283254
rect 30022 283018 65786 283254
rect 66022 283018 101786 283254
rect 102022 283018 137786 283254
rect 138022 283018 173786 283254
rect 174022 283018 209786 283254
rect 210022 283018 245786 283254
rect 246022 283018 281786 283254
rect 282022 283018 317786 283254
rect 318022 283018 353786 283254
rect 354022 283018 389786 283254
rect 390022 283018 425786 283254
rect 426022 283018 461786 283254
rect 462022 283018 497786 283254
rect 498022 283018 533786 283254
rect 534022 283018 569786 283254
rect 570022 283018 591942 283254
rect 592178 283018 592360 283254
rect -8436 282934 592360 283018
rect -8436 282698 -8254 282934
rect -8018 282698 29786 282934
rect 30022 282698 65786 282934
rect 66022 282698 101786 282934
rect 102022 282698 137786 282934
rect 138022 282698 173786 282934
rect 174022 282698 209786 282934
rect 210022 282698 245786 282934
rect 246022 282698 281786 282934
rect 282022 282698 317786 282934
rect 318022 282698 353786 282934
rect 354022 282698 389786 282934
rect 390022 282698 425786 282934
rect 426022 282698 461786 282934
rect 462022 282698 497786 282934
rect 498022 282698 533786 282934
rect 534022 282698 569786 282934
rect 570022 282698 591942 282934
rect 592178 282698 592360 282934
rect -8436 282676 592360 282698
rect -8436 282674 -7836 282676
rect 29604 282674 30204 282676
rect 65604 282674 66204 282676
rect 101604 282674 102204 282676
rect 137604 282674 138204 282676
rect 173604 282674 174204 282676
rect 209604 282674 210204 282676
rect 245604 282674 246204 282676
rect 281604 282674 282204 282676
rect 317604 282674 318204 282676
rect 353604 282674 354204 282676
rect 389604 282674 390204 282676
rect 425604 282674 426204 282676
rect 461604 282674 462204 282676
rect 497604 282674 498204 282676
rect 533604 282674 534204 282676
rect 569604 282674 570204 282676
rect 591760 282674 592360 282676
rect -6596 279676 -5996 279678
rect 26004 279676 26604 279678
rect 62004 279676 62604 279678
rect 98004 279676 98604 279678
rect 134004 279676 134604 279678
rect 170004 279676 170604 279678
rect 206004 279676 206604 279678
rect 242004 279676 242604 279678
rect 278004 279676 278604 279678
rect 314004 279676 314604 279678
rect 350004 279676 350604 279678
rect 386004 279676 386604 279678
rect 422004 279676 422604 279678
rect 458004 279676 458604 279678
rect 494004 279676 494604 279678
rect 530004 279676 530604 279678
rect 566004 279676 566604 279678
rect 589920 279676 590520 279678
rect -6596 279654 590520 279676
rect -6596 279418 -6414 279654
rect -6178 279418 26186 279654
rect 26422 279418 62186 279654
rect 62422 279418 98186 279654
rect 98422 279418 134186 279654
rect 134422 279418 170186 279654
rect 170422 279418 206186 279654
rect 206422 279418 242186 279654
rect 242422 279418 278186 279654
rect 278422 279418 314186 279654
rect 314422 279418 350186 279654
rect 350422 279418 386186 279654
rect 386422 279418 422186 279654
rect 422422 279418 458186 279654
rect 458422 279418 494186 279654
rect 494422 279418 530186 279654
rect 530422 279418 566186 279654
rect 566422 279418 590102 279654
rect 590338 279418 590520 279654
rect -6596 279334 590520 279418
rect -6596 279098 -6414 279334
rect -6178 279098 26186 279334
rect 26422 279098 62186 279334
rect 62422 279098 98186 279334
rect 98422 279098 134186 279334
rect 134422 279098 170186 279334
rect 170422 279098 206186 279334
rect 206422 279098 242186 279334
rect 242422 279098 278186 279334
rect 278422 279098 314186 279334
rect 314422 279098 350186 279334
rect 350422 279098 386186 279334
rect 386422 279098 422186 279334
rect 422422 279098 458186 279334
rect 458422 279098 494186 279334
rect 494422 279098 530186 279334
rect 530422 279098 566186 279334
rect 566422 279098 590102 279334
rect 590338 279098 590520 279334
rect -6596 279076 590520 279098
rect -6596 279074 -5996 279076
rect 26004 279074 26604 279076
rect 62004 279074 62604 279076
rect 98004 279074 98604 279076
rect 134004 279074 134604 279076
rect 170004 279074 170604 279076
rect 206004 279074 206604 279076
rect 242004 279074 242604 279076
rect 278004 279074 278604 279076
rect 314004 279074 314604 279076
rect 350004 279074 350604 279076
rect 386004 279074 386604 279076
rect 422004 279074 422604 279076
rect 458004 279074 458604 279076
rect 494004 279074 494604 279076
rect 530004 279074 530604 279076
rect 566004 279074 566604 279076
rect 589920 279074 590520 279076
rect -4756 276076 -4156 276078
rect 22404 276076 23004 276078
rect 58404 276076 59004 276078
rect 94404 276076 95004 276078
rect 130404 276076 131004 276078
rect 166404 276076 167004 276078
rect 202404 276076 203004 276078
rect 238404 276076 239004 276078
rect 274404 276076 275004 276078
rect 310404 276076 311004 276078
rect 346404 276076 347004 276078
rect 382404 276076 383004 276078
rect 418404 276076 419004 276078
rect 454404 276076 455004 276078
rect 490404 276076 491004 276078
rect 526404 276076 527004 276078
rect 562404 276076 563004 276078
rect 588080 276076 588680 276078
rect -4756 276054 588680 276076
rect -4756 275818 -4574 276054
rect -4338 275818 22586 276054
rect 22822 275818 58586 276054
rect 58822 275818 94586 276054
rect 94822 275818 130586 276054
rect 130822 275818 166586 276054
rect 166822 275818 202586 276054
rect 202822 275818 238586 276054
rect 238822 275818 274586 276054
rect 274822 275818 310586 276054
rect 310822 275818 346586 276054
rect 346822 275818 382586 276054
rect 382822 275818 418586 276054
rect 418822 275818 454586 276054
rect 454822 275818 490586 276054
rect 490822 275818 526586 276054
rect 526822 275818 562586 276054
rect 562822 275818 588262 276054
rect 588498 275818 588680 276054
rect -4756 275734 588680 275818
rect -4756 275498 -4574 275734
rect -4338 275498 22586 275734
rect 22822 275498 58586 275734
rect 58822 275498 94586 275734
rect 94822 275498 130586 275734
rect 130822 275498 166586 275734
rect 166822 275498 202586 275734
rect 202822 275498 238586 275734
rect 238822 275498 274586 275734
rect 274822 275498 310586 275734
rect 310822 275498 346586 275734
rect 346822 275498 382586 275734
rect 382822 275498 418586 275734
rect 418822 275498 454586 275734
rect 454822 275498 490586 275734
rect 490822 275498 526586 275734
rect 526822 275498 562586 275734
rect 562822 275498 588262 275734
rect 588498 275498 588680 275734
rect -4756 275476 588680 275498
rect -4756 275474 -4156 275476
rect 22404 275474 23004 275476
rect 58404 275474 59004 275476
rect 94404 275474 95004 275476
rect 130404 275474 131004 275476
rect 166404 275474 167004 275476
rect 202404 275474 203004 275476
rect 238404 275474 239004 275476
rect 274404 275474 275004 275476
rect 310404 275474 311004 275476
rect 346404 275474 347004 275476
rect 382404 275474 383004 275476
rect 418404 275474 419004 275476
rect 454404 275474 455004 275476
rect 490404 275474 491004 275476
rect 526404 275474 527004 275476
rect 562404 275474 563004 275476
rect 588080 275474 588680 275476
rect -2916 272476 -2316 272478
rect 18804 272476 19404 272478
rect 54804 272476 55404 272478
rect 90804 272476 91404 272478
rect 126804 272476 127404 272478
rect 162804 272476 163404 272478
rect 198804 272476 199404 272478
rect 234804 272476 235404 272478
rect 270804 272476 271404 272478
rect 306804 272476 307404 272478
rect 342804 272476 343404 272478
rect 378804 272476 379404 272478
rect 414804 272476 415404 272478
rect 450804 272476 451404 272478
rect 486804 272476 487404 272478
rect 522804 272476 523404 272478
rect 558804 272476 559404 272478
rect 586240 272476 586840 272478
rect -2916 272454 586840 272476
rect -2916 272218 -2734 272454
rect -2498 272218 18986 272454
rect 19222 272218 54986 272454
rect 55222 272218 90986 272454
rect 91222 272218 126986 272454
rect 127222 272218 162986 272454
rect 163222 272218 198986 272454
rect 199222 272218 234986 272454
rect 235222 272218 270986 272454
rect 271222 272218 306986 272454
rect 307222 272218 342986 272454
rect 343222 272218 378986 272454
rect 379222 272218 414986 272454
rect 415222 272218 450986 272454
rect 451222 272218 486986 272454
rect 487222 272218 522986 272454
rect 523222 272218 558986 272454
rect 559222 272218 586422 272454
rect 586658 272218 586840 272454
rect -2916 272134 586840 272218
rect -2916 271898 -2734 272134
rect -2498 271898 18986 272134
rect 19222 271898 54986 272134
rect 55222 271898 90986 272134
rect 91222 271898 126986 272134
rect 127222 271898 162986 272134
rect 163222 271898 198986 272134
rect 199222 271898 234986 272134
rect 235222 271898 270986 272134
rect 271222 271898 306986 272134
rect 307222 271898 342986 272134
rect 343222 271898 378986 272134
rect 379222 271898 414986 272134
rect 415222 271898 450986 272134
rect 451222 271898 486986 272134
rect 487222 271898 522986 272134
rect 523222 271898 558986 272134
rect 559222 271898 586422 272134
rect 586658 271898 586840 272134
rect -2916 271876 586840 271898
rect -2916 271874 -2316 271876
rect 18804 271874 19404 271876
rect 54804 271874 55404 271876
rect 90804 271874 91404 271876
rect 126804 271874 127404 271876
rect 162804 271874 163404 271876
rect 198804 271874 199404 271876
rect 234804 271874 235404 271876
rect 270804 271874 271404 271876
rect 306804 271874 307404 271876
rect 342804 271874 343404 271876
rect 378804 271874 379404 271876
rect 414804 271874 415404 271876
rect 450804 271874 451404 271876
rect 486804 271874 487404 271876
rect 522804 271874 523404 271876
rect 558804 271874 559404 271876
rect 586240 271874 586840 271876
rect -7516 265276 -6916 265278
rect 11604 265276 12204 265278
rect 47604 265276 48204 265278
rect 83604 265276 84204 265278
rect 119604 265276 120204 265278
rect 155604 265276 156204 265278
rect 191604 265276 192204 265278
rect 227604 265276 228204 265278
rect 263604 265276 264204 265278
rect 299604 265276 300204 265278
rect 335604 265276 336204 265278
rect 371604 265276 372204 265278
rect 407604 265276 408204 265278
rect 443604 265276 444204 265278
rect 479604 265276 480204 265278
rect 515604 265276 516204 265278
rect 551604 265276 552204 265278
rect 590840 265276 591440 265278
rect -8436 265254 592360 265276
rect -8436 265018 -7334 265254
rect -7098 265018 11786 265254
rect 12022 265018 47786 265254
rect 48022 265018 83786 265254
rect 84022 265018 119786 265254
rect 120022 265018 155786 265254
rect 156022 265018 191786 265254
rect 192022 265018 227786 265254
rect 228022 265018 263786 265254
rect 264022 265018 299786 265254
rect 300022 265018 335786 265254
rect 336022 265018 371786 265254
rect 372022 265018 407786 265254
rect 408022 265018 443786 265254
rect 444022 265018 479786 265254
rect 480022 265018 515786 265254
rect 516022 265018 551786 265254
rect 552022 265018 591022 265254
rect 591258 265018 592360 265254
rect -8436 264934 592360 265018
rect -8436 264698 -7334 264934
rect -7098 264698 11786 264934
rect 12022 264698 47786 264934
rect 48022 264698 83786 264934
rect 84022 264698 119786 264934
rect 120022 264698 155786 264934
rect 156022 264698 191786 264934
rect 192022 264698 227786 264934
rect 228022 264698 263786 264934
rect 264022 264698 299786 264934
rect 300022 264698 335786 264934
rect 336022 264698 371786 264934
rect 372022 264698 407786 264934
rect 408022 264698 443786 264934
rect 444022 264698 479786 264934
rect 480022 264698 515786 264934
rect 516022 264698 551786 264934
rect 552022 264698 591022 264934
rect 591258 264698 592360 264934
rect -8436 264676 592360 264698
rect -7516 264674 -6916 264676
rect 11604 264674 12204 264676
rect 47604 264674 48204 264676
rect 83604 264674 84204 264676
rect 119604 264674 120204 264676
rect 155604 264674 156204 264676
rect 191604 264674 192204 264676
rect 227604 264674 228204 264676
rect 263604 264674 264204 264676
rect 299604 264674 300204 264676
rect 335604 264674 336204 264676
rect 371604 264674 372204 264676
rect 407604 264674 408204 264676
rect 443604 264674 444204 264676
rect 479604 264674 480204 264676
rect 515604 264674 516204 264676
rect 551604 264674 552204 264676
rect 590840 264674 591440 264676
rect -5676 261676 -5076 261678
rect 8004 261676 8604 261678
rect 44004 261676 44604 261678
rect 80004 261676 80604 261678
rect 116004 261676 116604 261678
rect 152004 261676 152604 261678
rect 188004 261676 188604 261678
rect 224004 261676 224604 261678
rect 260004 261676 260604 261678
rect 296004 261676 296604 261678
rect 332004 261676 332604 261678
rect 368004 261676 368604 261678
rect 404004 261676 404604 261678
rect 440004 261676 440604 261678
rect 476004 261676 476604 261678
rect 512004 261676 512604 261678
rect 548004 261676 548604 261678
rect 589000 261676 589600 261678
rect -6596 261654 590520 261676
rect -6596 261418 -5494 261654
rect -5258 261418 8186 261654
rect 8422 261418 44186 261654
rect 44422 261418 80186 261654
rect 80422 261418 116186 261654
rect 116422 261418 152186 261654
rect 152422 261418 188186 261654
rect 188422 261418 224186 261654
rect 224422 261418 260186 261654
rect 260422 261418 296186 261654
rect 296422 261418 332186 261654
rect 332422 261418 368186 261654
rect 368422 261418 404186 261654
rect 404422 261418 440186 261654
rect 440422 261418 476186 261654
rect 476422 261418 512186 261654
rect 512422 261418 548186 261654
rect 548422 261418 589182 261654
rect 589418 261418 590520 261654
rect -6596 261334 590520 261418
rect -6596 261098 -5494 261334
rect -5258 261098 8186 261334
rect 8422 261098 44186 261334
rect 44422 261098 80186 261334
rect 80422 261098 116186 261334
rect 116422 261098 152186 261334
rect 152422 261098 188186 261334
rect 188422 261098 224186 261334
rect 224422 261098 260186 261334
rect 260422 261098 296186 261334
rect 296422 261098 332186 261334
rect 332422 261098 368186 261334
rect 368422 261098 404186 261334
rect 404422 261098 440186 261334
rect 440422 261098 476186 261334
rect 476422 261098 512186 261334
rect 512422 261098 548186 261334
rect 548422 261098 589182 261334
rect 589418 261098 590520 261334
rect -6596 261076 590520 261098
rect -5676 261074 -5076 261076
rect 8004 261074 8604 261076
rect 44004 261074 44604 261076
rect 80004 261074 80604 261076
rect 116004 261074 116604 261076
rect 152004 261074 152604 261076
rect 188004 261074 188604 261076
rect 224004 261074 224604 261076
rect 260004 261074 260604 261076
rect 296004 261074 296604 261076
rect 332004 261074 332604 261076
rect 368004 261074 368604 261076
rect 404004 261074 404604 261076
rect 440004 261074 440604 261076
rect 476004 261074 476604 261076
rect 512004 261074 512604 261076
rect 548004 261074 548604 261076
rect 589000 261074 589600 261076
rect -3836 258076 -3236 258078
rect 4404 258076 5004 258078
rect 40404 258076 41004 258078
rect 76404 258076 77004 258078
rect 112404 258076 113004 258078
rect 148404 258076 149004 258078
rect 184404 258076 185004 258078
rect 220404 258076 221004 258078
rect 256404 258076 257004 258078
rect 292404 258076 293004 258078
rect 328404 258076 329004 258078
rect 364404 258076 365004 258078
rect 400404 258076 401004 258078
rect 436404 258076 437004 258078
rect 472404 258076 473004 258078
rect 508404 258076 509004 258078
rect 544404 258076 545004 258078
rect 580404 258076 581004 258078
rect 587160 258076 587760 258078
rect -4756 258054 588680 258076
rect -4756 257818 -3654 258054
rect -3418 257818 4586 258054
rect 4822 257818 40586 258054
rect 40822 257818 76586 258054
rect 76822 257818 112586 258054
rect 112822 257818 148586 258054
rect 148822 257818 184586 258054
rect 184822 257818 220586 258054
rect 220822 257818 256586 258054
rect 256822 257818 292586 258054
rect 292822 257818 328586 258054
rect 328822 257818 364586 258054
rect 364822 257818 400586 258054
rect 400822 257818 436586 258054
rect 436822 257818 472586 258054
rect 472822 257818 508586 258054
rect 508822 257818 544586 258054
rect 544822 257818 580586 258054
rect 580822 257818 587342 258054
rect 587578 257818 588680 258054
rect -4756 257734 588680 257818
rect -4756 257498 -3654 257734
rect -3418 257498 4586 257734
rect 4822 257498 40586 257734
rect 40822 257498 76586 257734
rect 76822 257498 112586 257734
rect 112822 257498 148586 257734
rect 148822 257498 184586 257734
rect 184822 257498 220586 257734
rect 220822 257498 256586 257734
rect 256822 257498 292586 257734
rect 292822 257498 328586 257734
rect 328822 257498 364586 257734
rect 364822 257498 400586 257734
rect 400822 257498 436586 257734
rect 436822 257498 472586 257734
rect 472822 257498 508586 257734
rect 508822 257498 544586 257734
rect 544822 257498 580586 257734
rect 580822 257498 587342 257734
rect 587578 257498 588680 257734
rect -4756 257476 588680 257498
rect -3836 257474 -3236 257476
rect 4404 257474 5004 257476
rect 40404 257474 41004 257476
rect 76404 257474 77004 257476
rect 112404 257474 113004 257476
rect 148404 257474 149004 257476
rect 184404 257474 185004 257476
rect 220404 257474 221004 257476
rect 256404 257474 257004 257476
rect 292404 257474 293004 257476
rect 328404 257474 329004 257476
rect 364404 257474 365004 257476
rect 400404 257474 401004 257476
rect 436404 257474 437004 257476
rect 472404 257474 473004 257476
rect 508404 257474 509004 257476
rect 544404 257474 545004 257476
rect 580404 257474 581004 257476
rect 587160 257474 587760 257476
rect -1996 254476 -1396 254478
rect 804 254476 1404 254478
rect 36804 254476 37404 254478
rect 72804 254476 73404 254478
rect 108804 254476 109404 254478
rect 144804 254476 145404 254478
rect 180804 254476 181404 254478
rect 216804 254476 217404 254478
rect 252804 254476 253404 254478
rect 288804 254476 289404 254478
rect 324804 254476 325404 254478
rect 360804 254476 361404 254478
rect 396804 254476 397404 254478
rect 432804 254476 433404 254478
rect 468804 254476 469404 254478
rect 504804 254476 505404 254478
rect 540804 254476 541404 254478
rect 576804 254476 577404 254478
rect 585320 254476 585920 254478
rect -2916 254454 586840 254476
rect -2916 254218 -1814 254454
rect -1578 254218 986 254454
rect 1222 254218 36986 254454
rect 37222 254218 72986 254454
rect 73222 254218 108986 254454
rect 109222 254218 144986 254454
rect 145222 254218 180986 254454
rect 181222 254218 216986 254454
rect 217222 254218 252986 254454
rect 253222 254218 288986 254454
rect 289222 254218 324986 254454
rect 325222 254218 360986 254454
rect 361222 254218 396986 254454
rect 397222 254218 432986 254454
rect 433222 254218 468986 254454
rect 469222 254218 504986 254454
rect 505222 254218 540986 254454
rect 541222 254218 576986 254454
rect 577222 254218 585502 254454
rect 585738 254218 586840 254454
rect -2916 254134 586840 254218
rect -2916 253898 -1814 254134
rect -1578 253898 986 254134
rect 1222 253898 36986 254134
rect 37222 253898 72986 254134
rect 73222 253898 108986 254134
rect 109222 253898 144986 254134
rect 145222 253898 180986 254134
rect 181222 253898 216986 254134
rect 217222 253898 252986 254134
rect 253222 253898 288986 254134
rect 289222 253898 324986 254134
rect 325222 253898 360986 254134
rect 361222 253898 396986 254134
rect 397222 253898 432986 254134
rect 433222 253898 468986 254134
rect 469222 253898 504986 254134
rect 505222 253898 540986 254134
rect 541222 253898 576986 254134
rect 577222 253898 585502 254134
rect 585738 253898 586840 254134
rect -2916 253876 586840 253898
rect -1996 253874 -1396 253876
rect 804 253874 1404 253876
rect 36804 253874 37404 253876
rect 72804 253874 73404 253876
rect 108804 253874 109404 253876
rect 144804 253874 145404 253876
rect 180804 253874 181404 253876
rect 216804 253874 217404 253876
rect 252804 253874 253404 253876
rect 288804 253874 289404 253876
rect 324804 253874 325404 253876
rect 360804 253874 361404 253876
rect 396804 253874 397404 253876
rect 432804 253874 433404 253876
rect 468804 253874 469404 253876
rect 504804 253874 505404 253876
rect 540804 253874 541404 253876
rect 576804 253874 577404 253876
rect 585320 253874 585920 253876
rect -8436 247276 -7836 247278
rect 29604 247276 30204 247278
rect 65604 247276 66204 247278
rect 101604 247276 102204 247278
rect 137604 247276 138204 247278
rect 173604 247276 174204 247278
rect 209604 247276 210204 247278
rect 245604 247276 246204 247278
rect 281604 247276 282204 247278
rect 317604 247276 318204 247278
rect 353604 247276 354204 247278
rect 389604 247276 390204 247278
rect 425604 247276 426204 247278
rect 461604 247276 462204 247278
rect 497604 247276 498204 247278
rect 533604 247276 534204 247278
rect 569604 247276 570204 247278
rect 591760 247276 592360 247278
rect -8436 247254 592360 247276
rect -8436 247018 -8254 247254
rect -8018 247018 29786 247254
rect 30022 247018 65786 247254
rect 66022 247018 101786 247254
rect 102022 247018 137786 247254
rect 138022 247018 173786 247254
rect 174022 247018 209786 247254
rect 210022 247018 245786 247254
rect 246022 247018 281786 247254
rect 282022 247018 317786 247254
rect 318022 247018 353786 247254
rect 354022 247018 389786 247254
rect 390022 247018 425786 247254
rect 426022 247018 461786 247254
rect 462022 247018 497786 247254
rect 498022 247018 533786 247254
rect 534022 247018 569786 247254
rect 570022 247018 591942 247254
rect 592178 247018 592360 247254
rect -8436 246934 592360 247018
rect -8436 246698 -8254 246934
rect -8018 246698 29786 246934
rect 30022 246698 65786 246934
rect 66022 246698 101786 246934
rect 102022 246698 137786 246934
rect 138022 246698 173786 246934
rect 174022 246698 209786 246934
rect 210022 246698 245786 246934
rect 246022 246698 281786 246934
rect 282022 246698 317786 246934
rect 318022 246698 353786 246934
rect 354022 246698 389786 246934
rect 390022 246698 425786 246934
rect 426022 246698 461786 246934
rect 462022 246698 497786 246934
rect 498022 246698 533786 246934
rect 534022 246698 569786 246934
rect 570022 246698 591942 246934
rect 592178 246698 592360 246934
rect -8436 246676 592360 246698
rect -8436 246674 -7836 246676
rect 29604 246674 30204 246676
rect 65604 246674 66204 246676
rect 101604 246674 102204 246676
rect 137604 246674 138204 246676
rect 173604 246674 174204 246676
rect 209604 246674 210204 246676
rect 245604 246674 246204 246676
rect 281604 246674 282204 246676
rect 317604 246674 318204 246676
rect 353604 246674 354204 246676
rect 389604 246674 390204 246676
rect 425604 246674 426204 246676
rect 461604 246674 462204 246676
rect 497604 246674 498204 246676
rect 533604 246674 534204 246676
rect 569604 246674 570204 246676
rect 591760 246674 592360 246676
rect -6596 243676 -5996 243678
rect 26004 243676 26604 243678
rect 62004 243676 62604 243678
rect 98004 243676 98604 243678
rect 134004 243676 134604 243678
rect 170004 243676 170604 243678
rect 206004 243676 206604 243678
rect 242004 243676 242604 243678
rect 278004 243676 278604 243678
rect 314004 243676 314604 243678
rect 350004 243676 350604 243678
rect 386004 243676 386604 243678
rect 422004 243676 422604 243678
rect 458004 243676 458604 243678
rect 494004 243676 494604 243678
rect 530004 243676 530604 243678
rect 566004 243676 566604 243678
rect 589920 243676 590520 243678
rect -6596 243654 590520 243676
rect -6596 243418 -6414 243654
rect -6178 243418 26186 243654
rect 26422 243418 62186 243654
rect 62422 243418 98186 243654
rect 98422 243418 134186 243654
rect 134422 243418 170186 243654
rect 170422 243418 206186 243654
rect 206422 243418 242186 243654
rect 242422 243418 278186 243654
rect 278422 243418 314186 243654
rect 314422 243418 350186 243654
rect 350422 243418 386186 243654
rect 386422 243418 422186 243654
rect 422422 243418 458186 243654
rect 458422 243418 494186 243654
rect 494422 243418 530186 243654
rect 530422 243418 566186 243654
rect 566422 243418 590102 243654
rect 590338 243418 590520 243654
rect -6596 243334 590520 243418
rect -6596 243098 -6414 243334
rect -6178 243098 26186 243334
rect 26422 243098 62186 243334
rect 62422 243098 98186 243334
rect 98422 243098 134186 243334
rect 134422 243098 170186 243334
rect 170422 243098 206186 243334
rect 206422 243098 242186 243334
rect 242422 243098 278186 243334
rect 278422 243098 314186 243334
rect 314422 243098 350186 243334
rect 350422 243098 386186 243334
rect 386422 243098 422186 243334
rect 422422 243098 458186 243334
rect 458422 243098 494186 243334
rect 494422 243098 530186 243334
rect 530422 243098 566186 243334
rect 566422 243098 590102 243334
rect 590338 243098 590520 243334
rect -6596 243076 590520 243098
rect -6596 243074 -5996 243076
rect 26004 243074 26604 243076
rect 62004 243074 62604 243076
rect 98004 243074 98604 243076
rect 134004 243074 134604 243076
rect 170004 243074 170604 243076
rect 206004 243074 206604 243076
rect 242004 243074 242604 243076
rect 278004 243074 278604 243076
rect 314004 243074 314604 243076
rect 350004 243074 350604 243076
rect 386004 243074 386604 243076
rect 422004 243074 422604 243076
rect 458004 243074 458604 243076
rect 494004 243074 494604 243076
rect 530004 243074 530604 243076
rect 566004 243074 566604 243076
rect 589920 243074 590520 243076
rect -4756 240076 -4156 240078
rect 22404 240076 23004 240078
rect 58404 240076 59004 240078
rect 94404 240076 95004 240078
rect 130404 240076 131004 240078
rect 166404 240076 167004 240078
rect 202404 240076 203004 240078
rect 238404 240076 239004 240078
rect 274404 240076 275004 240078
rect 310404 240076 311004 240078
rect 346404 240076 347004 240078
rect 382404 240076 383004 240078
rect 418404 240076 419004 240078
rect 454404 240076 455004 240078
rect 490404 240076 491004 240078
rect 526404 240076 527004 240078
rect 562404 240076 563004 240078
rect 588080 240076 588680 240078
rect -4756 240054 588680 240076
rect -4756 239818 -4574 240054
rect -4338 239818 22586 240054
rect 22822 239818 58586 240054
rect 58822 239818 94586 240054
rect 94822 239818 130586 240054
rect 130822 239818 166586 240054
rect 166822 239818 202586 240054
rect 202822 239818 238586 240054
rect 238822 239818 274586 240054
rect 274822 239818 310586 240054
rect 310822 239818 346586 240054
rect 346822 239818 382586 240054
rect 382822 239818 418586 240054
rect 418822 239818 454586 240054
rect 454822 239818 490586 240054
rect 490822 239818 526586 240054
rect 526822 239818 562586 240054
rect 562822 239818 588262 240054
rect 588498 239818 588680 240054
rect -4756 239734 588680 239818
rect -4756 239498 -4574 239734
rect -4338 239498 22586 239734
rect 22822 239498 58586 239734
rect 58822 239498 94586 239734
rect 94822 239498 130586 239734
rect 130822 239498 166586 239734
rect 166822 239498 202586 239734
rect 202822 239498 238586 239734
rect 238822 239498 274586 239734
rect 274822 239498 310586 239734
rect 310822 239498 346586 239734
rect 346822 239498 382586 239734
rect 382822 239498 418586 239734
rect 418822 239498 454586 239734
rect 454822 239498 490586 239734
rect 490822 239498 526586 239734
rect 526822 239498 562586 239734
rect 562822 239498 588262 239734
rect 588498 239498 588680 239734
rect -4756 239476 588680 239498
rect -4756 239474 -4156 239476
rect 22404 239474 23004 239476
rect 58404 239474 59004 239476
rect 94404 239474 95004 239476
rect 130404 239474 131004 239476
rect 166404 239474 167004 239476
rect 202404 239474 203004 239476
rect 238404 239474 239004 239476
rect 274404 239474 275004 239476
rect 310404 239474 311004 239476
rect 346404 239474 347004 239476
rect 382404 239474 383004 239476
rect 418404 239474 419004 239476
rect 454404 239474 455004 239476
rect 490404 239474 491004 239476
rect 526404 239474 527004 239476
rect 562404 239474 563004 239476
rect 588080 239474 588680 239476
rect -2916 236476 -2316 236478
rect 18804 236476 19404 236478
rect 54804 236476 55404 236478
rect 90804 236476 91404 236478
rect 126804 236476 127404 236478
rect 162804 236476 163404 236478
rect 198804 236476 199404 236478
rect 234804 236476 235404 236478
rect 270804 236476 271404 236478
rect 306804 236476 307404 236478
rect 342804 236476 343404 236478
rect 378804 236476 379404 236478
rect 414804 236476 415404 236478
rect 450804 236476 451404 236478
rect 486804 236476 487404 236478
rect 522804 236476 523404 236478
rect 558804 236476 559404 236478
rect 586240 236476 586840 236478
rect -2916 236454 586840 236476
rect -2916 236218 -2734 236454
rect -2498 236218 18986 236454
rect 19222 236218 54986 236454
rect 55222 236218 90986 236454
rect 91222 236218 126986 236454
rect 127222 236218 162986 236454
rect 163222 236218 198986 236454
rect 199222 236218 234986 236454
rect 235222 236218 270986 236454
rect 271222 236218 306986 236454
rect 307222 236218 342986 236454
rect 343222 236218 378986 236454
rect 379222 236218 414986 236454
rect 415222 236218 450986 236454
rect 451222 236218 486986 236454
rect 487222 236218 522986 236454
rect 523222 236218 558986 236454
rect 559222 236218 586422 236454
rect 586658 236218 586840 236454
rect -2916 236134 586840 236218
rect -2916 235898 -2734 236134
rect -2498 235898 18986 236134
rect 19222 235898 54986 236134
rect 55222 235898 90986 236134
rect 91222 235898 126986 236134
rect 127222 235898 162986 236134
rect 163222 235898 198986 236134
rect 199222 235898 234986 236134
rect 235222 235898 270986 236134
rect 271222 235898 306986 236134
rect 307222 235898 342986 236134
rect 343222 235898 378986 236134
rect 379222 235898 414986 236134
rect 415222 235898 450986 236134
rect 451222 235898 486986 236134
rect 487222 235898 522986 236134
rect 523222 235898 558986 236134
rect 559222 235898 586422 236134
rect 586658 235898 586840 236134
rect -2916 235876 586840 235898
rect -2916 235874 -2316 235876
rect 18804 235874 19404 235876
rect 54804 235874 55404 235876
rect 90804 235874 91404 235876
rect 126804 235874 127404 235876
rect 162804 235874 163404 235876
rect 198804 235874 199404 235876
rect 234804 235874 235404 235876
rect 270804 235874 271404 235876
rect 306804 235874 307404 235876
rect 342804 235874 343404 235876
rect 378804 235874 379404 235876
rect 414804 235874 415404 235876
rect 450804 235874 451404 235876
rect 486804 235874 487404 235876
rect 522804 235874 523404 235876
rect 558804 235874 559404 235876
rect 586240 235874 586840 235876
rect -7516 229276 -6916 229278
rect 11604 229276 12204 229278
rect 47604 229276 48204 229278
rect 83604 229276 84204 229278
rect 119604 229276 120204 229278
rect 155604 229276 156204 229278
rect 191604 229276 192204 229278
rect 227604 229276 228204 229278
rect 263604 229276 264204 229278
rect 299604 229276 300204 229278
rect 335604 229276 336204 229278
rect 371604 229276 372204 229278
rect 407604 229276 408204 229278
rect 443604 229276 444204 229278
rect 479604 229276 480204 229278
rect 515604 229276 516204 229278
rect 551604 229276 552204 229278
rect 590840 229276 591440 229278
rect -8436 229254 592360 229276
rect -8436 229018 -7334 229254
rect -7098 229018 11786 229254
rect 12022 229018 47786 229254
rect 48022 229018 83786 229254
rect 84022 229018 119786 229254
rect 120022 229018 155786 229254
rect 156022 229018 191786 229254
rect 192022 229018 227786 229254
rect 228022 229018 263786 229254
rect 264022 229018 299786 229254
rect 300022 229018 335786 229254
rect 336022 229018 371786 229254
rect 372022 229018 407786 229254
rect 408022 229018 443786 229254
rect 444022 229018 479786 229254
rect 480022 229018 515786 229254
rect 516022 229018 551786 229254
rect 552022 229018 591022 229254
rect 591258 229018 592360 229254
rect -8436 228934 592360 229018
rect -8436 228698 -7334 228934
rect -7098 228698 11786 228934
rect 12022 228698 47786 228934
rect 48022 228698 83786 228934
rect 84022 228698 119786 228934
rect 120022 228698 155786 228934
rect 156022 228698 191786 228934
rect 192022 228698 227786 228934
rect 228022 228698 263786 228934
rect 264022 228698 299786 228934
rect 300022 228698 335786 228934
rect 336022 228698 371786 228934
rect 372022 228698 407786 228934
rect 408022 228698 443786 228934
rect 444022 228698 479786 228934
rect 480022 228698 515786 228934
rect 516022 228698 551786 228934
rect 552022 228698 591022 228934
rect 591258 228698 592360 228934
rect -8436 228676 592360 228698
rect -7516 228674 -6916 228676
rect 11604 228674 12204 228676
rect 47604 228674 48204 228676
rect 83604 228674 84204 228676
rect 119604 228674 120204 228676
rect 155604 228674 156204 228676
rect 191604 228674 192204 228676
rect 227604 228674 228204 228676
rect 263604 228674 264204 228676
rect 299604 228674 300204 228676
rect 335604 228674 336204 228676
rect 371604 228674 372204 228676
rect 407604 228674 408204 228676
rect 443604 228674 444204 228676
rect 479604 228674 480204 228676
rect 515604 228674 516204 228676
rect 551604 228674 552204 228676
rect 590840 228674 591440 228676
rect -5676 225676 -5076 225678
rect 8004 225676 8604 225678
rect 44004 225676 44604 225678
rect 80004 225676 80604 225678
rect 116004 225676 116604 225678
rect 152004 225676 152604 225678
rect 188004 225676 188604 225678
rect 224004 225676 224604 225678
rect 260004 225676 260604 225678
rect 296004 225676 296604 225678
rect 332004 225676 332604 225678
rect 368004 225676 368604 225678
rect 404004 225676 404604 225678
rect 440004 225676 440604 225678
rect 476004 225676 476604 225678
rect 512004 225676 512604 225678
rect 548004 225676 548604 225678
rect 589000 225676 589600 225678
rect -6596 225654 590520 225676
rect -6596 225418 -5494 225654
rect -5258 225418 8186 225654
rect 8422 225418 44186 225654
rect 44422 225418 80186 225654
rect 80422 225418 116186 225654
rect 116422 225418 152186 225654
rect 152422 225418 188186 225654
rect 188422 225418 224186 225654
rect 224422 225418 260186 225654
rect 260422 225418 296186 225654
rect 296422 225418 332186 225654
rect 332422 225418 368186 225654
rect 368422 225418 404186 225654
rect 404422 225418 440186 225654
rect 440422 225418 476186 225654
rect 476422 225418 512186 225654
rect 512422 225418 548186 225654
rect 548422 225418 589182 225654
rect 589418 225418 590520 225654
rect -6596 225334 590520 225418
rect -6596 225098 -5494 225334
rect -5258 225098 8186 225334
rect 8422 225098 44186 225334
rect 44422 225098 80186 225334
rect 80422 225098 116186 225334
rect 116422 225098 152186 225334
rect 152422 225098 188186 225334
rect 188422 225098 224186 225334
rect 224422 225098 260186 225334
rect 260422 225098 296186 225334
rect 296422 225098 332186 225334
rect 332422 225098 368186 225334
rect 368422 225098 404186 225334
rect 404422 225098 440186 225334
rect 440422 225098 476186 225334
rect 476422 225098 512186 225334
rect 512422 225098 548186 225334
rect 548422 225098 589182 225334
rect 589418 225098 590520 225334
rect -6596 225076 590520 225098
rect -5676 225074 -5076 225076
rect 8004 225074 8604 225076
rect 44004 225074 44604 225076
rect 80004 225074 80604 225076
rect 116004 225074 116604 225076
rect 152004 225074 152604 225076
rect 188004 225074 188604 225076
rect 224004 225074 224604 225076
rect 260004 225074 260604 225076
rect 296004 225074 296604 225076
rect 332004 225074 332604 225076
rect 368004 225074 368604 225076
rect 404004 225074 404604 225076
rect 440004 225074 440604 225076
rect 476004 225074 476604 225076
rect 512004 225074 512604 225076
rect 548004 225074 548604 225076
rect 589000 225074 589600 225076
rect -3836 222076 -3236 222078
rect 4404 222076 5004 222078
rect 40404 222076 41004 222078
rect 76404 222076 77004 222078
rect 112404 222076 113004 222078
rect 148404 222076 149004 222078
rect 184404 222076 185004 222078
rect 220404 222076 221004 222078
rect 256404 222076 257004 222078
rect 292404 222076 293004 222078
rect 328404 222076 329004 222078
rect 364404 222076 365004 222078
rect 400404 222076 401004 222078
rect 436404 222076 437004 222078
rect 472404 222076 473004 222078
rect 508404 222076 509004 222078
rect 544404 222076 545004 222078
rect 580404 222076 581004 222078
rect 587160 222076 587760 222078
rect -4756 222054 588680 222076
rect -4756 221818 -3654 222054
rect -3418 221818 4586 222054
rect 4822 221818 40586 222054
rect 40822 221818 76586 222054
rect 76822 221818 112586 222054
rect 112822 221818 148586 222054
rect 148822 221818 184586 222054
rect 184822 221818 220586 222054
rect 220822 221818 256586 222054
rect 256822 221818 292586 222054
rect 292822 221818 328586 222054
rect 328822 221818 364586 222054
rect 364822 221818 400586 222054
rect 400822 221818 436586 222054
rect 436822 221818 472586 222054
rect 472822 221818 508586 222054
rect 508822 221818 544586 222054
rect 544822 221818 580586 222054
rect 580822 221818 587342 222054
rect 587578 221818 588680 222054
rect -4756 221734 588680 221818
rect -4756 221498 -3654 221734
rect -3418 221498 4586 221734
rect 4822 221498 40586 221734
rect 40822 221498 76586 221734
rect 76822 221498 112586 221734
rect 112822 221498 148586 221734
rect 148822 221498 184586 221734
rect 184822 221498 220586 221734
rect 220822 221498 256586 221734
rect 256822 221498 292586 221734
rect 292822 221498 328586 221734
rect 328822 221498 364586 221734
rect 364822 221498 400586 221734
rect 400822 221498 436586 221734
rect 436822 221498 472586 221734
rect 472822 221498 508586 221734
rect 508822 221498 544586 221734
rect 544822 221498 580586 221734
rect 580822 221498 587342 221734
rect 587578 221498 588680 221734
rect -4756 221476 588680 221498
rect -3836 221474 -3236 221476
rect 4404 221474 5004 221476
rect 40404 221474 41004 221476
rect 76404 221474 77004 221476
rect 112404 221474 113004 221476
rect 148404 221474 149004 221476
rect 184404 221474 185004 221476
rect 220404 221474 221004 221476
rect 256404 221474 257004 221476
rect 292404 221474 293004 221476
rect 328404 221474 329004 221476
rect 364404 221474 365004 221476
rect 400404 221474 401004 221476
rect 436404 221474 437004 221476
rect 472404 221474 473004 221476
rect 508404 221474 509004 221476
rect 544404 221474 545004 221476
rect 580404 221474 581004 221476
rect 587160 221474 587760 221476
rect -1996 218476 -1396 218478
rect 804 218476 1404 218478
rect 36804 218476 37404 218478
rect 72804 218476 73404 218478
rect 108804 218476 109404 218478
rect 144804 218476 145404 218478
rect 180804 218476 181404 218478
rect 216804 218476 217404 218478
rect 252804 218476 253404 218478
rect 288804 218476 289404 218478
rect 324804 218476 325404 218478
rect 360804 218476 361404 218478
rect 396804 218476 397404 218478
rect 432804 218476 433404 218478
rect 468804 218476 469404 218478
rect 504804 218476 505404 218478
rect 540804 218476 541404 218478
rect 576804 218476 577404 218478
rect 585320 218476 585920 218478
rect -2916 218454 586840 218476
rect -2916 218218 -1814 218454
rect -1578 218218 986 218454
rect 1222 218218 36986 218454
rect 37222 218218 72986 218454
rect 73222 218218 108986 218454
rect 109222 218218 144986 218454
rect 145222 218218 180986 218454
rect 181222 218218 216986 218454
rect 217222 218218 252986 218454
rect 253222 218218 288986 218454
rect 289222 218218 324986 218454
rect 325222 218218 360986 218454
rect 361222 218218 396986 218454
rect 397222 218218 432986 218454
rect 433222 218218 468986 218454
rect 469222 218218 504986 218454
rect 505222 218218 540986 218454
rect 541222 218218 576986 218454
rect 577222 218218 585502 218454
rect 585738 218218 586840 218454
rect -2916 218134 586840 218218
rect -2916 217898 -1814 218134
rect -1578 217898 986 218134
rect 1222 217898 36986 218134
rect 37222 217898 72986 218134
rect 73222 217898 108986 218134
rect 109222 217898 144986 218134
rect 145222 217898 180986 218134
rect 181222 217898 216986 218134
rect 217222 217898 252986 218134
rect 253222 217898 288986 218134
rect 289222 217898 324986 218134
rect 325222 217898 360986 218134
rect 361222 217898 396986 218134
rect 397222 217898 432986 218134
rect 433222 217898 468986 218134
rect 469222 217898 504986 218134
rect 505222 217898 540986 218134
rect 541222 217898 576986 218134
rect 577222 217898 585502 218134
rect 585738 217898 586840 218134
rect -2916 217876 586840 217898
rect -1996 217874 -1396 217876
rect 804 217874 1404 217876
rect 36804 217874 37404 217876
rect 72804 217874 73404 217876
rect 108804 217874 109404 217876
rect 144804 217874 145404 217876
rect 180804 217874 181404 217876
rect 216804 217874 217404 217876
rect 252804 217874 253404 217876
rect 288804 217874 289404 217876
rect 324804 217874 325404 217876
rect 360804 217874 361404 217876
rect 396804 217874 397404 217876
rect 432804 217874 433404 217876
rect 468804 217874 469404 217876
rect 504804 217874 505404 217876
rect 540804 217874 541404 217876
rect 576804 217874 577404 217876
rect 585320 217874 585920 217876
rect -8436 211276 -7836 211278
rect 29604 211276 30204 211278
rect 65604 211276 66204 211278
rect 101604 211276 102204 211278
rect 137604 211276 138204 211278
rect 173604 211276 174204 211278
rect 209604 211276 210204 211278
rect 245604 211276 246204 211278
rect 281604 211276 282204 211278
rect 317604 211276 318204 211278
rect 353604 211276 354204 211278
rect 389604 211276 390204 211278
rect 425604 211276 426204 211278
rect 461604 211276 462204 211278
rect 497604 211276 498204 211278
rect 533604 211276 534204 211278
rect 569604 211276 570204 211278
rect 591760 211276 592360 211278
rect -8436 211254 592360 211276
rect -8436 211018 -8254 211254
rect -8018 211018 29786 211254
rect 30022 211018 65786 211254
rect 66022 211018 101786 211254
rect 102022 211018 137786 211254
rect 138022 211018 173786 211254
rect 174022 211018 209786 211254
rect 210022 211018 245786 211254
rect 246022 211018 281786 211254
rect 282022 211018 317786 211254
rect 318022 211018 353786 211254
rect 354022 211018 389786 211254
rect 390022 211018 425786 211254
rect 426022 211018 461786 211254
rect 462022 211018 497786 211254
rect 498022 211018 533786 211254
rect 534022 211018 569786 211254
rect 570022 211018 591942 211254
rect 592178 211018 592360 211254
rect -8436 210934 592360 211018
rect -8436 210698 -8254 210934
rect -8018 210698 29786 210934
rect 30022 210698 65786 210934
rect 66022 210698 101786 210934
rect 102022 210698 137786 210934
rect 138022 210698 173786 210934
rect 174022 210698 209786 210934
rect 210022 210698 245786 210934
rect 246022 210698 281786 210934
rect 282022 210698 317786 210934
rect 318022 210698 353786 210934
rect 354022 210698 389786 210934
rect 390022 210698 425786 210934
rect 426022 210698 461786 210934
rect 462022 210698 497786 210934
rect 498022 210698 533786 210934
rect 534022 210698 569786 210934
rect 570022 210698 591942 210934
rect 592178 210698 592360 210934
rect -8436 210676 592360 210698
rect -8436 210674 -7836 210676
rect 29604 210674 30204 210676
rect 65604 210674 66204 210676
rect 101604 210674 102204 210676
rect 137604 210674 138204 210676
rect 173604 210674 174204 210676
rect 209604 210674 210204 210676
rect 245604 210674 246204 210676
rect 281604 210674 282204 210676
rect 317604 210674 318204 210676
rect 353604 210674 354204 210676
rect 389604 210674 390204 210676
rect 425604 210674 426204 210676
rect 461604 210674 462204 210676
rect 497604 210674 498204 210676
rect 533604 210674 534204 210676
rect 569604 210674 570204 210676
rect 591760 210674 592360 210676
rect -6596 207676 -5996 207678
rect 26004 207676 26604 207678
rect 62004 207676 62604 207678
rect 98004 207676 98604 207678
rect 134004 207676 134604 207678
rect 170004 207676 170604 207678
rect 206004 207676 206604 207678
rect 242004 207676 242604 207678
rect 278004 207676 278604 207678
rect 314004 207676 314604 207678
rect 350004 207676 350604 207678
rect 386004 207676 386604 207678
rect 422004 207676 422604 207678
rect 458004 207676 458604 207678
rect 494004 207676 494604 207678
rect 530004 207676 530604 207678
rect 566004 207676 566604 207678
rect 589920 207676 590520 207678
rect -6596 207654 590520 207676
rect -6596 207418 -6414 207654
rect -6178 207418 26186 207654
rect 26422 207418 62186 207654
rect 62422 207418 98186 207654
rect 98422 207418 134186 207654
rect 134422 207418 170186 207654
rect 170422 207418 206186 207654
rect 206422 207418 242186 207654
rect 242422 207418 278186 207654
rect 278422 207418 314186 207654
rect 314422 207418 350186 207654
rect 350422 207418 386186 207654
rect 386422 207418 422186 207654
rect 422422 207418 458186 207654
rect 458422 207418 494186 207654
rect 494422 207418 530186 207654
rect 530422 207418 566186 207654
rect 566422 207418 590102 207654
rect 590338 207418 590520 207654
rect -6596 207334 590520 207418
rect -6596 207098 -6414 207334
rect -6178 207098 26186 207334
rect 26422 207098 62186 207334
rect 62422 207098 98186 207334
rect 98422 207098 134186 207334
rect 134422 207098 170186 207334
rect 170422 207098 206186 207334
rect 206422 207098 242186 207334
rect 242422 207098 278186 207334
rect 278422 207098 314186 207334
rect 314422 207098 350186 207334
rect 350422 207098 386186 207334
rect 386422 207098 422186 207334
rect 422422 207098 458186 207334
rect 458422 207098 494186 207334
rect 494422 207098 530186 207334
rect 530422 207098 566186 207334
rect 566422 207098 590102 207334
rect 590338 207098 590520 207334
rect -6596 207076 590520 207098
rect -6596 207074 -5996 207076
rect 26004 207074 26604 207076
rect 62004 207074 62604 207076
rect 98004 207074 98604 207076
rect 134004 207074 134604 207076
rect 170004 207074 170604 207076
rect 206004 207074 206604 207076
rect 242004 207074 242604 207076
rect 278004 207074 278604 207076
rect 314004 207074 314604 207076
rect 350004 207074 350604 207076
rect 386004 207074 386604 207076
rect 422004 207074 422604 207076
rect 458004 207074 458604 207076
rect 494004 207074 494604 207076
rect 530004 207074 530604 207076
rect 566004 207074 566604 207076
rect 589920 207074 590520 207076
rect -4756 204076 -4156 204078
rect 22404 204076 23004 204078
rect 58404 204076 59004 204078
rect 94404 204076 95004 204078
rect 130404 204076 131004 204078
rect 166404 204076 167004 204078
rect 202404 204076 203004 204078
rect 238404 204076 239004 204078
rect 274404 204076 275004 204078
rect 310404 204076 311004 204078
rect 346404 204076 347004 204078
rect 382404 204076 383004 204078
rect 418404 204076 419004 204078
rect 454404 204076 455004 204078
rect 490404 204076 491004 204078
rect 526404 204076 527004 204078
rect 562404 204076 563004 204078
rect 588080 204076 588680 204078
rect -4756 204054 588680 204076
rect -4756 203818 -4574 204054
rect -4338 203818 22586 204054
rect 22822 203818 58586 204054
rect 58822 203818 94586 204054
rect 94822 203818 130586 204054
rect 130822 203818 166586 204054
rect 166822 203818 202586 204054
rect 202822 203818 238586 204054
rect 238822 203818 274586 204054
rect 274822 203818 310586 204054
rect 310822 203818 346586 204054
rect 346822 203818 382586 204054
rect 382822 203818 418586 204054
rect 418822 203818 454586 204054
rect 454822 203818 490586 204054
rect 490822 203818 526586 204054
rect 526822 203818 562586 204054
rect 562822 203818 588262 204054
rect 588498 203818 588680 204054
rect -4756 203734 588680 203818
rect -4756 203498 -4574 203734
rect -4338 203498 22586 203734
rect 22822 203498 58586 203734
rect 58822 203498 94586 203734
rect 94822 203498 130586 203734
rect 130822 203498 166586 203734
rect 166822 203498 202586 203734
rect 202822 203498 238586 203734
rect 238822 203498 274586 203734
rect 274822 203498 310586 203734
rect 310822 203498 346586 203734
rect 346822 203498 382586 203734
rect 382822 203498 418586 203734
rect 418822 203498 454586 203734
rect 454822 203498 490586 203734
rect 490822 203498 526586 203734
rect 526822 203498 562586 203734
rect 562822 203498 588262 203734
rect 588498 203498 588680 203734
rect -4756 203476 588680 203498
rect -4756 203474 -4156 203476
rect 22404 203474 23004 203476
rect 58404 203474 59004 203476
rect 94404 203474 95004 203476
rect 130404 203474 131004 203476
rect 166404 203474 167004 203476
rect 202404 203474 203004 203476
rect 238404 203474 239004 203476
rect 274404 203474 275004 203476
rect 310404 203474 311004 203476
rect 346404 203474 347004 203476
rect 382404 203474 383004 203476
rect 418404 203474 419004 203476
rect 454404 203474 455004 203476
rect 490404 203474 491004 203476
rect 526404 203474 527004 203476
rect 562404 203474 563004 203476
rect 588080 203474 588680 203476
rect -2916 200476 -2316 200478
rect 18804 200476 19404 200478
rect 54804 200476 55404 200478
rect 90804 200476 91404 200478
rect 126804 200476 127404 200478
rect 162804 200476 163404 200478
rect 198804 200476 199404 200478
rect 234804 200476 235404 200478
rect 270804 200476 271404 200478
rect 306804 200476 307404 200478
rect 342804 200476 343404 200478
rect 378804 200476 379404 200478
rect 414804 200476 415404 200478
rect 450804 200476 451404 200478
rect 486804 200476 487404 200478
rect 522804 200476 523404 200478
rect 558804 200476 559404 200478
rect 586240 200476 586840 200478
rect -2916 200454 586840 200476
rect -2916 200218 -2734 200454
rect -2498 200218 18986 200454
rect 19222 200218 54986 200454
rect 55222 200218 90986 200454
rect 91222 200218 126986 200454
rect 127222 200218 162986 200454
rect 163222 200218 198986 200454
rect 199222 200218 234986 200454
rect 235222 200218 270986 200454
rect 271222 200218 306986 200454
rect 307222 200218 342986 200454
rect 343222 200218 378986 200454
rect 379222 200218 414986 200454
rect 415222 200218 450986 200454
rect 451222 200218 486986 200454
rect 487222 200218 522986 200454
rect 523222 200218 558986 200454
rect 559222 200218 586422 200454
rect 586658 200218 586840 200454
rect -2916 200134 586840 200218
rect -2916 199898 -2734 200134
rect -2498 199898 18986 200134
rect 19222 199898 54986 200134
rect 55222 199898 90986 200134
rect 91222 199898 126986 200134
rect 127222 199898 162986 200134
rect 163222 199898 198986 200134
rect 199222 199898 234986 200134
rect 235222 199898 270986 200134
rect 271222 199898 306986 200134
rect 307222 199898 342986 200134
rect 343222 199898 378986 200134
rect 379222 199898 414986 200134
rect 415222 199898 450986 200134
rect 451222 199898 486986 200134
rect 487222 199898 522986 200134
rect 523222 199898 558986 200134
rect 559222 199898 586422 200134
rect 586658 199898 586840 200134
rect -2916 199876 586840 199898
rect -2916 199874 -2316 199876
rect 18804 199874 19404 199876
rect 54804 199874 55404 199876
rect 90804 199874 91404 199876
rect 126804 199874 127404 199876
rect 162804 199874 163404 199876
rect 198804 199874 199404 199876
rect 234804 199874 235404 199876
rect 270804 199874 271404 199876
rect 306804 199874 307404 199876
rect 342804 199874 343404 199876
rect 378804 199874 379404 199876
rect 414804 199874 415404 199876
rect 450804 199874 451404 199876
rect 486804 199874 487404 199876
rect 522804 199874 523404 199876
rect 558804 199874 559404 199876
rect 586240 199874 586840 199876
rect -7516 193276 -6916 193278
rect 11604 193276 12204 193278
rect 47604 193276 48204 193278
rect 83604 193276 84204 193278
rect 119604 193276 120204 193278
rect 155604 193276 156204 193278
rect 191604 193276 192204 193278
rect 227604 193276 228204 193278
rect 263604 193276 264204 193278
rect 299604 193276 300204 193278
rect 335604 193276 336204 193278
rect 371604 193276 372204 193278
rect 407604 193276 408204 193278
rect 443604 193276 444204 193278
rect 479604 193276 480204 193278
rect 515604 193276 516204 193278
rect 551604 193276 552204 193278
rect 590840 193276 591440 193278
rect -8436 193254 592360 193276
rect -8436 193018 -7334 193254
rect -7098 193018 11786 193254
rect 12022 193018 47786 193254
rect 48022 193018 83786 193254
rect 84022 193018 119786 193254
rect 120022 193018 155786 193254
rect 156022 193018 191786 193254
rect 192022 193018 227786 193254
rect 228022 193018 263786 193254
rect 264022 193018 299786 193254
rect 300022 193018 335786 193254
rect 336022 193018 371786 193254
rect 372022 193018 407786 193254
rect 408022 193018 443786 193254
rect 444022 193018 479786 193254
rect 480022 193018 515786 193254
rect 516022 193018 551786 193254
rect 552022 193018 591022 193254
rect 591258 193018 592360 193254
rect -8436 192934 592360 193018
rect -8436 192698 -7334 192934
rect -7098 192698 11786 192934
rect 12022 192698 47786 192934
rect 48022 192698 83786 192934
rect 84022 192698 119786 192934
rect 120022 192698 155786 192934
rect 156022 192698 191786 192934
rect 192022 192698 227786 192934
rect 228022 192698 263786 192934
rect 264022 192698 299786 192934
rect 300022 192698 335786 192934
rect 336022 192698 371786 192934
rect 372022 192698 407786 192934
rect 408022 192698 443786 192934
rect 444022 192698 479786 192934
rect 480022 192698 515786 192934
rect 516022 192698 551786 192934
rect 552022 192698 591022 192934
rect 591258 192698 592360 192934
rect -8436 192676 592360 192698
rect -7516 192674 -6916 192676
rect 11604 192674 12204 192676
rect 47604 192674 48204 192676
rect 83604 192674 84204 192676
rect 119604 192674 120204 192676
rect 155604 192674 156204 192676
rect 191604 192674 192204 192676
rect 227604 192674 228204 192676
rect 263604 192674 264204 192676
rect 299604 192674 300204 192676
rect 335604 192674 336204 192676
rect 371604 192674 372204 192676
rect 407604 192674 408204 192676
rect 443604 192674 444204 192676
rect 479604 192674 480204 192676
rect 515604 192674 516204 192676
rect 551604 192674 552204 192676
rect 590840 192674 591440 192676
rect -5676 189676 -5076 189678
rect 8004 189676 8604 189678
rect 44004 189676 44604 189678
rect 80004 189676 80604 189678
rect 116004 189676 116604 189678
rect 152004 189676 152604 189678
rect 188004 189676 188604 189678
rect 224004 189676 224604 189678
rect 260004 189676 260604 189678
rect 296004 189676 296604 189678
rect 332004 189676 332604 189678
rect 368004 189676 368604 189678
rect 404004 189676 404604 189678
rect 440004 189676 440604 189678
rect 476004 189676 476604 189678
rect 512004 189676 512604 189678
rect 548004 189676 548604 189678
rect 589000 189676 589600 189678
rect -6596 189654 590520 189676
rect -6596 189418 -5494 189654
rect -5258 189418 8186 189654
rect 8422 189418 44186 189654
rect 44422 189418 80186 189654
rect 80422 189418 116186 189654
rect 116422 189418 152186 189654
rect 152422 189418 188186 189654
rect 188422 189418 224186 189654
rect 224422 189418 260186 189654
rect 260422 189418 296186 189654
rect 296422 189418 332186 189654
rect 332422 189418 368186 189654
rect 368422 189418 404186 189654
rect 404422 189418 440186 189654
rect 440422 189418 476186 189654
rect 476422 189418 512186 189654
rect 512422 189418 548186 189654
rect 548422 189418 589182 189654
rect 589418 189418 590520 189654
rect -6596 189334 590520 189418
rect -6596 189098 -5494 189334
rect -5258 189098 8186 189334
rect 8422 189098 44186 189334
rect 44422 189098 80186 189334
rect 80422 189098 116186 189334
rect 116422 189098 152186 189334
rect 152422 189098 188186 189334
rect 188422 189098 224186 189334
rect 224422 189098 260186 189334
rect 260422 189098 296186 189334
rect 296422 189098 332186 189334
rect 332422 189098 368186 189334
rect 368422 189098 404186 189334
rect 404422 189098 440186 189334
rect 440422 189098 476186 189334
rect 476422 189098 512186 189334
rect 512422 189098 548186 189334
rect 548422 189098 589182 189334
rect 589418 189098 590520 189334
rect -6596 189076 590520 189098
rect -5676 189074 -5076 189076
rect 8004 189074 8604 189076
rect 44004 189074 44604 189076
rect 80004 189074 80604 189076
rect 116004 189074 116604 189076
rect 152004 189074 152604 189076
rect 188004 189074 188604 189076
rect 224004 189074 224604 189076
rect 260004 189074 260604 189076
rect 296004 189074 296604 189076
rect 332004 189074 332604 189076
rect 368004 189074 368604 189076
rect 404004 189074 404604 189076
rect 440004 189074 440604 189076
rect 476004 189074 476604 189076
rect 512004 189074 512604 189076
rect 548004 189074 548604 189076
rect 589000 189074 589600 189076
rect -3836 186076 -3236 186078
rect 4404 186076 5004 186078
rect 40404 186076 41004 186078
rect 76404 186076 77004 186078
rect 112404 186076 113004 186078
rect 148404 186076 149004 186078
rect 184404 186076 185004 186078
rect 220404 186076 221004 186078
rect 256404 186076 257004 186078
rect 292404 186076 293004 186078
rect 328404 186076 329004 186078
rect 364404 186076 365004 186078
rect 400404 186076 401004 186078
rect 436404 186076 437004 186078
rect 472404 186076 473004 186078
rect 508404 186076 509004 186078
rect 544404 186076 545004 186078
rect 580404 186076 581004 186078
rect 587160 186076 587760 186078
rect -4756 186054 588680 186076
rect -4756 185818 -3654 186054
rect -3418 185818 4586 186054
rect 4822 185818 40586 186054
rect 40822 185818 76586 186054
rect 76822 185818 112586 186054
rect 112822 185818 148586 186054
rect 148822 185818 184586 186054
rect 184822 185818 220586 186054
rect 220822 185818 256586 186054
rect 256822 185818 292586 186054
rect 292822 185818 328586 186054
rect 328822 185818 364586 186054
rect 364822 185818 400586 186054
rect 400822 185818 436586 186054
rect 436822 185818 472586 186054
rect 472822 185818 508586 186054
rect 508822 185818 544586 186054
rect 544822 185818 580586 186054
rect 580822 185818 587342 186054
rect 587578 185818 588680 186054
rect -4756 185734 588680 185818
rect -4756 185498 -3654 185734
rect -3418 185498 4586 185734
rect 4822 185498 40586 185734
rect 40822 185498 76586 185734
rect 76822 185498 112586 185734
rect 112822 185498 148586 185734
rect 148822 185498 184586 185734
rect 184822 185498 220586 185734
rect 220822 185498 256586 185734
rect 256822 185498 292586 185734
rect 292822 185498 328586 185734
rect 328822 185498 364586 185734
rect 364822 185498 400586 185734
rect 400822 185498 436586 185734
rect 436822 185498 472586 185734
rect 472822 185498 508586 185734
rect 508822 185498 544586 185734
rect 544822 185498 580586 185734
rect 580822 185498 587342 185734
rect 587578 185498 588680 185734
rect -4756 185476 588680 185498
rect -3836 185474 -3236 185476
rect 4404 185474 5004 185476
rect 40404 185474 41004 185476
rect 76404 185474 77004 185476
rect 112404 185474 113004 185476
rect 148404 185474 149004 185476
rect 184404 185474 185004 185476
rect 220404 185474 221004 185476
rect 256404 185474 257004 185476
rect 292404 185474 293004 185476
rect 328404 185474 329004 185476
rect 364404 185474 365004 185476
rect 400404 185474 401004 185476
rect 436404 185474 437004 185476
rect 472404 185474 473004 185476
rect 508404 185474 509004 185476
rect 544404 185474 545004 185476
rect 580404 185474 581004 185476
rect 587160 185474 587760 185476
rect -1996 182476 -1396 182478
rect 804 182476 1404 182478
rect 36804 182476 37404 182478
rect 72804 182476 73404 182478
rect 108804 182476 109404 182478
rect 144804 182476 145404 182478
rect 180804 182476 181404 182478
rect 216804 182476 217404 182478
rect 252804 182476 253404 182478
rect 288804 182476 289404 182478
rect 324804 182476 325404 182478
rect 360804 182476 361404 182478
rect 396804 182476 397404 182478
rect 432804 182476 433404 182478
rect 468804 182476 469404 182478
rect 504804 182476 505404 182478
rect 540804 182476 541404 182478
rect 576804 182476 577404 182478
rect 585320 182476 585920 182478
rect -2916 182454 586840 182476
rect -2916 182218 -1814 182454
rect -1578 182218 986 182454
rect 1222 182218 36986 182454
rect 37222 182218 72986 182454
rect 73222 182218 108986 182454
rect 109222 182218 144986 182454
rect 145222 182218 180986 182454
rect 181222 182218 216986 182454
rect 217222 182218 252986 182454
rect 253222 182218 288986 182454
rect 289222 182218 324986 182454
rect 325222 182218 360986 182454
rect 361222 182218 396986 182454
rect 397222 182218 432986 182454
rect 433222 182218 468986 182454
rect 469222 182218 504986 182454
rect 505222 182218 540986 182454
rect 541222 182218 576986 182454
rect 577222 182218 585502 182454
rect 585738 182218 586840 182454
rect -2916 182134 586840 182218
rect -2916 181898 -1814 182134
rect -1578 181898 986 182134
rect 1222 181898 36986 182134
rect 37222 181898 72986 182134
rect 73222 181898 108986 182134
rect 109222 181898 144986 182134
rect 145222 181898 180986 182134
rect 181222 181898 216986 182134
rect 217222 181898 252986 182134
rect 253222 181898 288986 182134
rect 289222 181898 324986 182134
rect 325222 181898 360986 182134
rect 361222 181898 396986 182134
rect 397222 181898 432986 182134
rect 433222 181898 468986 182134
rect 469222 181898 504986 182134
rect 505222 181898 540986 182134
rect 541222 181898 576986 182134
rect 577222 181898 585502 182134
rect 585738 181898 586840 182134
rect -2916 181876 586840 181898
rect -1996 181874 -1396 181876
rect 804 181874 1404 181876
rect 36804 181874 37404 181876
rect 72804 181874 73404 181876
rect 108804 181874 109404 181876
rect 144804 181874 145404 181876
rect 180804 181874 181404 181876
rect 216804 181874 217404 181876
rect 252804 181874 253404 181876
rect 288804 181874 289404 181876
rect 324804 181874 325404 181876
rect 360804 181874 361404 181876
rect 396804 181874 397404 181876
rect 432804 181874 433404 181876
rect 468804 181874 469404 181876
rect 504804 181874 505404 181876
rect 540804 181874 541404 181876
rect 576804 181874 577404 181876
rect 585320 181874 585920 181876
rect -8436 175276 -7836 175278
rect 29604 175276 30204 175278
rect 65604 175276 66204 175278
rect 101604 175276 102204 175278
rect 137604 175276 138204 175278
rect 173604 175276 174204 175278
rect 209604 175276 210204 175278
rect 245604 175276 246204 175278
rect 281604 175276 282204 175278
rect 317604 175276 318204 175278
rect 353604 175276 354204 175278
rect 389604 175276 390204 175278
rect 425604 175276 426204 175278
rect 461604 175276 462204 175278
rect 497604 175276 498204 175278
rect 533604 175276 534204 175278
rect 569604 175276 570204 175278
rect 591760 175276 592360 175278
rect -8436 175254 592360 175276
rect -8436 175018 -8254 175254
rect -8018 175018 29786 175254
rect 30022 175018 65786 175254
rect 66022 175018 101786 175254
rect 102022 175018 137786 175254
rect 138022 175018 173786 175254
rect 174022 175018 209786 175254
rect 210022 175018 245786 175254
rect 246022 175018 281786 175254
rect 282022 175018 317786 175254
rect 318022 175018 353786 175254
rect 354022 175018 389786 175254
rect 390022 175018 425786 175254
rect 426022 175018 461786 175254
rect 462022 175018 497786 175254
rect 498022 175018 533786 175254
rect 534022 175018 569786 175254
rect 570022 175018 591942 175254
rect 592178 175018 592360 175254
rect -8436 174934 592360 175018
rect -8436 174698 -8254 174934
rect -8018 174698 29786 174934
rect 30022 174698 65786 174934
rect 66022 174698 101786 174934
rect 102022 174698 137786 174934
rect 138022 174698 173786 174934
rect 174022 174698 209786 174934
rect 210022 174698 245786 174934
rect 246022 174698 281786 174934
rect 282022 174698 317786 174934
rect 318022 174698 353786 174934
rect 354022 174698 389786 174934
rect 390022 174698 425786 174934
rect 426022 174698 461786 174934
rect 462022 174698 497786 174934
rect 498022 174698 533786 174934
rect 534022 174698 569786 174934
rect 570022 174698 591942 174934
rect 592178 174698 592360 174934
rect -8436 174676 592360 174698
rect -8436 174674 -7836 174676
rect 29604 174674 30204 174676
rect 65604 174674 66204 174676
rect 101604 174674 102204 174676
rect 137604 174674 138204 174676
rect 173604 174674 174204 174676
rect 209604 174674 210204 174676
rect 245604 174674 246204 174676
rect 281604 174674 282204 174676
rect 317604 174674 318204 174676
rect 353604 174674 354204 174676
rect 389604 174674 390204 174676
rect 425604 174674 426204 174676
rect 461604 174674 462204 174676
rect 497604 174674 498204 174676
rect 533604 174674 534204 174676
rect 569604 174674 570204 174676
rect 591760 174674 592360 174676
rect -6596 171676 -5996 171678
rect 26004 171676 26604 171678
rect 62004 171676 62604 171678
rect 98004 171676 98604 171678
rect 134004 171676 134604 171678
rect 170004 171676 170604 171678
rect 206004 171676 206604 171678
rect 242004 171676 242604 171678
rect 278004 171676 278604 171678
rect 314004 171676 314604 171678
rect 350004 171676 350604 171678
rect 386004 171676 386604 171678
rect 422004 171676 422604 171678
rect 458004 171676 458604 171678
rect 494004 171676 494604 171678
rect 530004 171676 530604 171678
rect 566004 171676 566604 171678
rect 589920 171676 590520 171678
rect -6596 171654 590520 171676
rect -6596 171418 -6414 171654
rect -6178 171418 26186 171654
rect 26422 171418 62186 171654
rect 62422 171418 98186 171654
rect 98422 171418 134186 171654
rect 134422 171418 170186 171654
rect 170422 171418 206186 171654
rect 206422 171418 242186 171654
rect 242422 171418 278186 171654
rect 278422 171418 314186 171654
rect 314422 171418 350186 171654
rect 350422 171418 386186 171654
rect 386422 171418 422186 171654
rect 422422 171418 458186 171654
rect 458422 171418 494186 171654
rect 494422 171418 530186 171654
rect 530422 171418 566186 171654
rect 566422 171418 590102 171654
rect 590338 171418 590520 171654
rect -6596 171334 590520 171418
rect -6596 171098 -6414 171334
rect -6178 171098 26186 171334
rect 26422 171098 62186 171334
rect 62422 171098 98186 171334
rect 98422 171098 134186 171334
rect 134422 171098 170186 171334
rect 170422 171098 206186 171334
rect 206422 171098 242186 171334
rect 242422 171098 278186 171334
rect 278422 171098 314186 171334
rect 314422 171098 350186 171334
rect 350422 171098 386186 171334
rect 386422 171098 422186 171334
rect 422422 171098 458186 171334
rect 458422 171098 494186 171334
rect 494422 171098 530186 171334
rect 530422 171098 566186 171334
rect 566422 171098 590102 171334
rect 590338 171098 590520 171334
rect -6596 171076 590520 171098
rect -6596 171074 -5996 171076
rect 26004 171074 26604 171076
rect 62004 171074 62604 171076
rect 98004 171074 98604 171076
rect 134004 171074 134604 171076
rect 170004 171074 170604 171076
rect 206004 171074 206604 171076
rect 242004 171074 242604 171076
rect 278004 171074 278604 171076
rect 314004 171074 314604 171076
rect 350004 171074 350604 171076
rect 386004 171074 386604 171076
rect 422004 171074 422604 171076
rect 458004 171074 458604 171076
rect 494004 171074 494604 171076
rect 530004 171074 530604 171076
rect 566004 171074 566604 171076
rect 589920 171074 590520 171076
rect -4756 168076 -4156 168078
rect 22404 168076 23004 168078
rect 58404 168076 59004 168078
rect 94404 168076 95004 168078
rect 130404 168076 131004 168078
rect 166404 168076 167004 168078
rect 202404 168076 203004 168078
rect 238404 168076 239004 168078
rect 274404 168076 275004 168078
rect 310404 168076 311004 168078
rect 346404 168076 347004 168078
rect 382404 168076 383004 168078
rect 418404 168076 419004 168078
rect 454404 168076 455004 168078
rect 490404 168076 491004 168078
rect 526404 168076 527004 168078
rect 562404 168076 563004 168078
rect 588080 168076 588680 168078
rect -4756 168054 588680 168076
rect -4756 167818 -4574 168054
rect -4338 167818 22586 168054
rect 22822 167818 58586 168054
rect 58822 167818 94586 168054
rect 94822 167818 130586 168054
rect 130822 167818 166586 168054
rect 166822 167818 202586 168054
rect 202822 167818 238586 168054
rect 238822 167818 274586 168054
rect 274822 167818 310586 168054
rect 310822 167818 346586 168054
rect 346822 167818 382586 168054
rect 382822 167818 418586 168054
rect 418822 167818 454586 168054
rect 454822 167818 490586 168054
rect 490822 167818 526586 168054
rect 526822 167818 562586 168054
rect 562822 167818 588262 168054
rect 588498 167818 588680 168054
rect -4756 167734 588680 167818
rect -4756 167498 -4574 167734
rect -4338 167498 22586 167734
rect 22822 167498 58586 167734
rect 58822 167498 94586 167734
rect 94822 167498 130586 167734
rect 130822 167498 166586 167734
rect 166822 167498 202586 167734
rect 202822 167498 238586 167734
rect 238822 167498 274586 167734
rect 274822 167498 310586 167734
rect 310822 167498 346586 167734
rect 346822 167498 382586 167734
rect 382822 167498 418586 167734
rect 418822 167498 454586 167734
rect 454822 167498 490586 167734
rect 490822 167498 526586 167734
rect 526822 167498 562586 167734
rect 562822 167498 588262 167734
rect 588498 167498 588680 167734
rect -4756 167476 588680 167498
rect -4756 167474 -4156 167476
rect 22404 167474 23004 167476
rect 58404 167474 59004 167476
rect 94404 167474 95004 167476
rect 130404 167474 131004 167476
rect 166404 167474 167004 167476
rect 202404 167474 203004 167476
rect 238404 167474 239004 167476
rect 274404 167474 275004 167476
rect 310404 167474 311004 167476
rect 346404 167474 347004 167476
rect 382404 167474 383004 167476
rect 418404 167474 419004 167476
rect 454404 167474 455004 167476
rect 490404 167474 491004 167476
rect 526404 167474 527004 167476
rect 562404 167474 563004 167476
rect 588080 167474 588680 167476
rect -2916 164476 -2316 164478
rect 18804 164476 19404 164478
rect 54804 164476 55404 164478
rect 90804 164476 91404 164478
rect 126804 164476 127404 164478
rect 162804 164476 163404 164478
rect 198804 164476 199404 164478
rect 234804 164476 235404 164478
rect 270804 164476 271404 164478
rect 306804 164476 307404 164478
rect 342804 164476 343404 164478
rect 378804 164476 379404 164478
rect 414804 164476 415404 164478
rect 450804 164476 451404 164478
rect 486804 164476 487404 164478
rect 522804 164476 523404 164478
rect 558804 164476 559404 164478
rect 586240 164476 586840 164478
rect -2916 164454 586840 164476
rect -2916 164218 -2734 164454
rect -2498 164218 18986 164454
rect 19222 164218 54986 164454
rect 55222 164218 90986 164454
rect 91222 164218 126986 164454
rect 127222 164218 162986 164454
rect 163222 164218 198986 164454
rect 199222 164218 234986 164454
rect 235222 164218 270986 164454
rect 271222 164218 306986 164454
rect 307222 164218 342986 164454
rect 343222 164218 378986 164454
rect 379222 164218 414986 164454
rect 415222 164218 450986 164454
rect 451222 164218 486986 164454
rect 487222 164218 522986 164454
rect 523222 164218 558986 164454
rect 559222 164218 586422 164454
rect 586658 164218 586840 164454
rect -2916 164134 586840 164218
rect -2916 163898 -2734 164134
rect -2498 163898 18986 164134
rect 19222 163898 54986 164134
rect 55222 163898 90986 164134
rect 91222 163898 126986 164134
rect 127222 163898 162986 164134
rect 163222 163898 198986 164134
rect 199222 163898 234986 164134
rect 235222 163898 270986 164134
rect 271222 163898 306986 164134
rect 307222 163898 342986 164134
rect 343222 163898 378986 164134
rect 379222 163898 414986 164134
rect 415222 163898 450986 164134
rect 451222 163898 486986 164134
rect 487222 163898 522986 164134
rect 523222 163898 558986 164134
rect 559222 163898 586422 164134
rect 586658 163898 586840 164134
rect -2916 163876 586840 163898
rect -2916 163874 -2316 163876
rect 18804 163874 19404 163876
rect 54804 163874 55404 163876
rect 90804 163874 91404 163876
rect 126804 163874 127404 163876
rect 162804 163874 163404 163876
rect 198804 163874 199404 163876
rect 234804 163874 235404 163876
rect 270804 163874 271404 163876
rect 306804 163874 307404 163876
rect 342804 163874 343404 163876
rect 378804 163874 379404 163876
rect 414804 163874 415404 163876
rect 450804 163874 451404 163876
rect 486804 163874 487404 163876
rect 522804 163874 523404 163876
rect 558804 163874 559404 163876
rect 586240 163874 586840 163876
rect -7516 157276 -6916 157278
rect 11604 157276 12204 157278
rect 47604 157276 48204 157278
rect 83604 157276 84204 157278
rect 119604 157276 120204 157278
rect 155604 157276 156204 157278
rect 191604 157276 192204 157278
rect 227604 157276 228204 157278
rect 263604 157276 264204 157278
rect 299604 157276 300204 157278
rect 335604 157276 336204 157278
rect 371604 157276 372204 157278
rect 407604 157276 408204 157278
rect 443604 157276 444204 157278
rect 479604 157276 480204 157278
rect 515604 157276 516204 157278
rect 551604 157276 552204 157278
rect 590840 157276 591440 157278
rect -8436 157254 592360 157276
rect -8436 157018 -7334 157254
rect -7098 157018 11786 157254
rect 12022 157018 47786 157254
rect 48022 157018 83786 157254
rect 84022 157018 119786 157254
rect 120022 157018 155786 157254
rect 156022 157018 191786 157254
rect 192022 157018 227786 157254
rect 228022 157018 263786 157254
rect 264022 157018 299786 157254
rect 300022 157018 335786 157254
rect 336022 157018 371786 157254
rect 372022 157018 407786 157254
rect 408022 157018 443786 157254
rect 444022 157018 479786 157254
rect 480022 157018 515786 157254
rect 516022 157018 551786 157254
rect 552022 157018 591022 157254
rect 591258 157018 592360 157254
rect -8436 156934 592360 157018
rect -8436 156698 -7334 156934
rect -7098 156698 11786 156934
rect 12022 156698 47786 156934
rect 48022 156698 83786 156934
rect 84022 156698 119786 156934
rect 120022 156698 155786 156934
rect 156022 156698 191786 156934
rect 192022 156698 227786 156934
rect 228022 156698 263786 156934
rect 264022 156698 299786 156934
rect 300022 156698 335786 156934
rect 336022 156698 371786 156934
rect 372022 156698 407786 156934
rect 408022 156698 443786 156934
rect 444022 156698 479786 156934
rect 480022 156698 515786 156934
rect 516022 156698 551786 156934
rect 552022 156698 591022 156934
rect 591258 156698 592360 156934
rect -8436 156676 592360 156698
rect -7516 156674 -6916 156676
rect 11604 156674 12204 156676
rect 47604 156674 48204 156676
rect 83604 156674 84204 156676
rect 119604 156674 120204 156676
rect 155604 156674 156204 156676
rect 191604 156674 192204 156676
rect 227604 156674 228204 156676
rect 263604 156674 264204 156676
rect 299604 156674 300204 156676
rect 335604 156674 336204 156676
rect 371604 156674 372204 156676
rect 407604 156674 408204 156676
rect 443604 156674 444204 156676
rect 479604 156674 480204 156676
rect 515604 156674 516204 156676
rect 551604 156674 552204 156676
rect 590840 156674 591440 156676
rect -5676 153676 -5076 153678
rect 8004 153676 8604 153678
rect 44004 153676 44604 153678
rect 80004 153676 80604 153678
rect 116004 153676 116604 153678
rect 152004 153676 152604 153678
rect 188004 153676 188604 153678
rect 224004 153676 224604 153678
rect 260004 153676 260604 153678
rect 296004 153676 296604 153678
rect 332004 153676 332604 153678
rect 368004 153676 368604 153678
rect 404004 153676 404604 153678
rect 440004 153676 440604 153678
rect 476004 153676 476604 153678
rect 512004 153676 512604 153678
rect 548004 153676 548604 153678
rect 589000 153676 589600 153678
rect -6596 153654 590520 153676
rect -6596 153418 -5494 153654
rect -5258 153418 8186 153654
rect 8422 153418 44186 153654
rect 44422 153418 80186 153654
rect 80422 153418 116186 153654
rect 116422 153418 152186 153654
rect 152422 153418 188186 153654
rect 188422 153418 224186 153654
rect 224422 153418 260186 153654
rect 260422 153418 296186 153654
rect 296422 153418 332186 153654
rect 332422 153418 368186 153654
rect 368422 153418 404186 153654
rect 404422 153418 440186 153654
rect 440422 153418 476186 153654
rect 476422 153418 512186 153654
rect 512422 153418 548186 153654
rect 548422 153418 589182 153654
rect 589418 153418 590520 153654
rect -6596 153334 590520 153418
rect -6596 153098 -5494 153334
rect -5258 153098 8186 153334
rect 8422 153098 44186 153334
rect 44422 153098 80186 153334
rect 80422 153098 116186 153334
rect 116422 153098 152186 153334
rect 152422 153098 188186 153334
rect 188422 153098 224186 153334
rect 224422 153098 260186 153334
rect 260422 153098 296186 153334
rect 296422 153098 332186 153334
rect 332422 153098 368186 153334
rect 368422 153098 404186 153334
rect 404422 153098 440186 153334
rect 440422 153098 476186 153334
rect 476422 153098 512186 153334
rect 512422 153098 548186 153334
rect 548422 153098 589182 153334
rect 589418 153098 590520 153334
rect -6596 153076 590520 153098
rect -5676 153074 -5076 153076
rect 8004 153074 8604 153076
rect 44004 153074 44604 153076
rect 80004 153074 80604 153076
rect 116004 153074 116604 153076
rect 152004 153074 152604 153076
rect 188004 153074 188604 153076
rect 224004 153074 224604 153076
rect 260004 153074 260604 153076
rect 296004 153074 296604 153076
rect 332004 153074 332604 153076
rect 368004 153074 368604 153076
rect 404004 153074 404604 153076
rect 440004 153074 440604 153076
rect 476004 153074 476604 153076
rect 512004 153074 512604 153076
rect 548004 153074 548604 153076
rect 589000 153074 589600 153076
rect -3836 150076 -3236 150078
rect 4404 150076 5004 150078
rect 40404 150076 41004 150078
rect 76404 150076 77004 150078
rect 112404 150076 113004 150078
rect 148404 150076 149004 150078
rect 184404 150076 185004 150078
rect 220404 150076 221004 150078
rect 256404 150076 257004 150078
rect 292404 150076 293004 150078
rect 328404 150076 329004 150078
rect 364404 150076 365004 150078
rect 400404 150076 401004 150078
rect 436404 150076 437004 150078
rect 472404 150076 473004 150078
rect 508404 150076 509004 150078
rect 544404 150076 545004 150078
rect 580404 150076 581004 150078
rect 587160 150076 587760 150078
rect -4756 150054 588680 150076
rect -4756 149818 -3654 150054
rect -3418 149818 4586 150054
rect 4822 149818 40586 150054
rect 40822 149818 76586 150054
rect 76822 149818 112586 150054
rect 112822 149818 148586 150054
rect 148822 149818 184586 150054
rect 184822 149818 220586 150054
rect 220822 149818 256586 150054
rect 256822 149818 292586 150054
rect 292822 149818 328586 150054
rect 328822 149818 364586 150054
rect 364822 149818 400586 150054
rect 400822 149818 436586 150054
rect 436822 149818 472586 150054
rect 472822 149818 508586 150054
rect 508822 149818 544586 150054
rect 544822 149818 580586 150054
rect 580822 149818 587342 150054
rect 587578 149818 588680 150054
rect -4756 149734 588680 149818
rect -4756 149498 -3654 149734
rect -3418 149498 4586 149734
rect 4822 149498 40586 149734
rect 40822 149498 76586 149734
rect 76822 149498 112586 149734
rect 112822 149498 148586 149734
rect 148822 149498 184586 149734
rect 184822 149498 220586 149734
rect 220822 149498 256586 149734
rect 256822 149498 292586 149734
rect 292822 149498 328586 149734
rect 328822 149498 364586 149734
rect 364822 149498 400586 149734
rect 400822 149498 436586 149734
rect 436822 149498 472586 149734
rect 472822 149498 508586 149734
rect 508822 149498 544586 149734
rect 544822 149498 580586 149734
rect 580822 149498 587342 149734
rect 587578 149498 588680 149734
rect -4756 149476 588680 149498
rect -3836 149474 -3236 149476
rect 4404 149474 5004 149476
rect 40404 149474 41004 149476
rect 76404 149474 77004 149476
rect 112404 149474 113004 149476
rect 148404 149474 149004 149476
rect 184404 149474 185004 149476
rect 220404 149474 221004 149476
rect 256404 149474 257004 149476
rect 292404 149474 293004 149476
rect 328404 149474 329004 149476
rect 364404 149474 365004 149476
rect 400404 149474 401004 149476
rect 436404 149474 437004 149476
rect 472404 149474 473004 149476
rect 508404 149474 509004 149476
rect 544404 149474 545004 149476
rect 580404 149474 581004 149476
rect 587160 149474 587760 149476
rect -1996 146476 -1396 146478
rect 804 146476 1404 146478
rect 36804 146476 37404 146478
rect 72804 146476 73404 146478
rect 108804 146476 109404 146478
rect 144804 146476 145404 146478
rect 180804 146476 181404 146478
rect 216804 146476 217404 146478
rect 252804 146476 253404 146478
rect 288804 146476 289404 146478
rect 324804 146476 325404 146478
rect 360804 146476 361404 146478
rect 396804 146476 397404 146478
rect 432804 146476 433404 146478
rect 468804 146476 469404 146478
rect 504804 146476 505404 146478
rect 540804 146476 541404 146478
rect 576804 146476 577404 146478
rect 585320 146476 585920 146478
rect -2916 146454 586840 146476
rect -2916 146218 -1814 146454
rect -1578 146218 986 146454
rect 1222 146218 36986 146454
rect 37222 146218 72986 146454
rect 73222 146218 108986 146454
rect 109222 146218 144986 146454
rect 145222 146218 180986 146454
rect 181222 146218 216986 146454
rect 217222 146218 252986 146454
rect 253222 146218 288986 146454
rect 289222 146218 324986 146454
rect 325222 146218 360986 146454
rect 361222 146218 396986 146454
rect 397222 146218 432986 146454
rect 433222 146218 468986 146454
rect 469222 146218 504986 146454
rect 505222 146218 540986 146454
rect 541222 146218 576986 146454
rect 577222 146218 585502 146454
rect 585738 146218 586840 146454
rect -2916 146134 586840 146218
rect -2916 145898 -1814 146134
rect -1578 145898 986 146134
rect 1222 145898 36986 146134
rect 37222 145898 72986 146134
rect 73222 145898 108986 146134
rect 109222 145898 144986 146134
rect 145222 145898 180986 146134
rect 181222 145898 216986 146134
rect 217222 145898 252986 146134
rect 253222 145898 288986 146134
rect 289222 145898 324986 146134
rect 325222 145898 360986 146134
rect 361222 145898 396986 146134
rect 397222 145898 432986 146134
rect 433222 145898 468986 146134
rect 469222 145898 504986 146134
rect 505222 145898 540986 146134
rect 541222 145898 576986 146134
rect 577222 145898 585502 146134
rect 585738 145898 586840 146134
rect -2916 145876 586840 145898
rect -1996 145874 -1396 145876
rect 804 145874 1404 145876
rect 36804 145874 37404 145876
rect 72804 145874 73404 145876
rect 108804 145874 109404 145876
rect 144804 145874 145404 145876
rect 180804 145874 181404 145876
rect 216804 145874 217404 145876
rect 252804 145874 253404 145876
rect 288804 145874 289404 145876
rect 324804 145874 325404 145876
rect 360804 145874 361404 145876
rect 396804 145874 397404 145876
rect 432804 145874 433404 145876
rect 468804 145874 469404 145876
rect 504804 145874 505404 145876
rect 540804 145874 541404 145876
rect 576804 145874 577404 145876
rect 585320 145874 585920 145876
rect -8436 139276 -7836 139278
rect 29604 139276 30204 139278
rect 65604 139276 66204 139278
rect 101604 139276 102204 139278
rect 137604 139276 138204 139278
rect 173604 139276 174204 139278
rect 209604 139276 210204 139278
rect 245604 139276 246204 139278
rect 281604 139276 282204 139278
rect 317604 139276 318204 139278
rect 353604 139276 354204 139278
rect 389604 139276 390204 139278
rect 425604 139276 426204 139278
rect 461604 139276 462204 139278
rect 497604 139276 498204 139278
rect 533604 139276 534204 139278
rect 569604 139276 570204 139278
rect 591760 139276 592360 139278
rect -8436 139254 592360 139276
rect -8436 139018 -8254 139254
rect -8018 139018 29786 139254
rect 30022 139018 65786 139254
rect 66022 139018 101786 139254
rect 102022 139018 137786 139254
rect 138022 139018 173786 139254
rect 174022 139018 209786 139254
rect 210022 139018 245786 139254
rect 246022 139018 281786 139254
rect 282022 139018 317786 139254
rect 318022 139018 353786 139254
rect 354022 139018 389786 139254
rect 390022 139018 425786 139254
rect 426022 139018 461786 139254
rect 462022 139018 497786 139254
rect 498022 139018 533786 139254
rect 534022 139018 569786 139254
rect 570022 139018 591942 139254
rect 592178 139018 592360 139254
rect -8436 138934 592360 139018
rect -8436 138698 -8254 138934
rect -8018 138698 29786 138934
rect 30022 138698 65786 138934
rect 66022 138698 101786 138934
rect 102022 138698 137786 138934
rect 138022 138698 173786 138934
rect 174022 138698 209786 138934
rect 210022 138698 245786 138934
rect 246022 138698 281786 138934
rect 282022 138698 317786 138934
rect 318022 138698 353786 138934
rect 354022 138698 389786 138934
rect 390022 138698 425786 138934
rect 426022 138698 461786 138934
rect 462022 138698 497786 138934
rect 498022 138698 533786 138934
rect 534022 138698 569786 138934
rect 570022 138698 591942 138934
rect 592178 138698 592360 138934
rect -8436 138676 592360 138698
rect -8436 138674 -7836 138676
rect 29604 138674 30204 138676
rect 65604 138674 66204 138676
rect 101604 138674 102204 138676
rect 137604 138674 138204 138676
rect 173604 138674 174204 138676
rect 209604 138674 210204 138676
rect 245604 138674 246204 138676
rect 281604 138674 282204 138676
rect 317604 138674 318204 138676
rect 353604 138674 354204 138676
rect 389604 138674 390204 138676
rect 425604 138674 426204 138676
rect 461604 138674 462204 138676
rect 497604 138674 498204 138676
rect 533604 138674 534204 138676
rect 569604 138674 570204 138676
rect 591760 138674 592360 138676
rect -6596 135676 -5996 135678
rect 26004 135676 26604 135678
rect 62004 135676 62604 135678
rect 98004 135676 98604 135678
rect 134004 135676 134604 135678
rect 170004 135676 170604 135678
rect 206004 135676 206604 135678
rect 242004 135676 242604 135678
rect 278004 135676 278604 135678
rect 314004 135676 314604 135678
rect 350004 135676 350604 135678
rect 386004 135676 386604 135678
rect 422004 135676 422604 135678
rect 458004 135676 458604 135678
rect 494004 135676 494604 135678
rect 530004 135676 530604 135678
rect 566004 135676 566604 135678
rect 589920 135676 590520 135678
rect -6596 135654 590520 135676
rect -6596 135418 -6414 135654
rect -6178 135418 26186 135654
rect 26422 135418 62186 135654
rect 62422 135418 98186 135654
rect 98422 135418 134186 135654
rect 134422 135418 170186 135654
rect 170422 135418 206186 135654
rect 206422 135418 242186 135654
rect 242422 135418 278186 135654
rect 278422 135418 314186 135654
rect 314422 135418 350186 135654
rect 350422 135418 386186 135654
rect 386422 135418 422186 135654
rect 422422 135418 458186 135654
rect 458422 135418 494186 135654
rect 494422 135418 530186 135654
rect 530422 135418 566186 135654
rect 566422 135418 590102 135654
rect 590338 135418 590520 135654
rect -6596 135334 590520 135418
rect -6596 135098 -6414 135334
rect -6178 135098 26186 135334
rect 26422 135098 62186 135334
rect 62422 135098 98186 135334
rect 98422 135098 134186 135334
rect 134422 135098 170186 135334
rect 170422 135098 206186 135334
rect 206422 135098 242186 135334
rect 242422 135098 278186 135334
rect 278422 135098 314186 135334
rect 314422 135098 350186 135334
rect 350422 135098 386186 135334
rect 386422 135098 422186 135334
rect 422422 135098 458186 135334
rect 458422 135098 494186 135334
rect 494422 135098 530186 135334
rect 530422 135098 566186 135334
rect 566422 135098 590102 135334
rect 590338 135098 590520 135334
rect -6596 135076 590520 135098
rect -6596 135074 -5996 135076
rect 26004 135074 26604 135076
rect 62004 135074 62604 135076
rect 98004 135074 98604 135076
rect 134004 135074 134604 135076
rect 170004 135074 170604 135076
rect 206004 135074 206604 135076
rect 242004 135074 242604 135076
rect 278004 135074 278604 135076
rect 314004 135074 314604 135076
rect 350004 135074 350604 135076
rect 386004 135074 386604 135076
rect 422004 135074 422604 135076
rect 458004 135074 458604 135076
rect 494004 135074 494604 135076
rect 530004 135074 530604 135076
rect 566004 135074 566604 135076
rect 589920 135074 590520 135076
rect -4756 132076 -4156 132078
rect 22404 132076 23004 132078
rect 58404 132076 59004 132078
rect 94404 132076 95004 132078
rect 130404 132076 131004 132078
rect 166404 132076 167004 132078
rect 202404 132076 203004 132078
rect 238404 132076 239004 132078
rect 274404 132076 275004 132078
rect 310404 132076 311004 132078
rect 346404 132076 347004 132078
rect 382404 132076 383004 132078
rect 418404 132076 419004 132078
rect 454404 132076 455004 132078
rect 490404 132076 491004 132078
rect 526404 132076 527004 132078
rect 562404 132076 563004 132078
rect 588080 132076 588680 132078
rect -4756 132054 588680 132076
rect -4756 131818 -4574 132054
rect -4338 131818 22586 132054
rect 22822 131818 58586 132054
rect 58822 131818 94586 132054
rect 94822 131818 130586 132054
rect 130822 131818 166586 132054
rect 166822 131818 202586 132054
rect 202822 131818 238586 132054
rect 238822 131818 274586 132054
rect 274822 131818 310586 132054
rect 310822 131818 346586 132054
rect 346822 131818 382586 132054
rect 382822 131818 418586 132054
rect 418822 131818 454586 132054
rect 454822 131818 490586 132054
rect 490822 131818 526586 132054
rect 526822 131818 562586 132054
rect 562822 131818 588262 132054
rect 588498 131818 588680 132054
rect -4756 131734 588680 131818
rect -4756 131498 -4574 131734
rect -4338 131498 22586 131734
rect 22822 131498 58586 131734
rect 58822 131498 94586 131734
rect 94822 131498 130586 131734
rect 130822 131498 166586 131734
rect 166822 131498 202586 131734
rect 202822 131498 238586 131734
rect 238822 131498 274586 131734
rect 274822 131498 310586 131734
rect 310822 131498 346586 131734
rect 346822 131498 382586 131734
rect 382822 131498 418586 131734
rect 418822 131498 454586 131734
rect 454822 131498 490586 131734
rect 490822 131498 526586 131734
rect 526822 131498 562586 131734
rect 562822 131498 588262 131734
rect 588498 131498 588680 131734
rect -4756 131476 588680 131498
rect -4756 131474 -4156 131476
rect 22404 131474 23004 131476
rect 58404 131474 59004 131476
rect 94404 131474 95004 131476
rect 130404 131474 131004 131476
rect 166404 131474 167004 131476
rect 202404 131474 203004 131476
rect 238404 131474 239004 131476
rect 274404 131474 275004 131476
rect 310404 131474 311004 131476
rect 346404 131474 347004 131476
rect 382404 131474 383004 131476
rect 418404 131474 419004 131476
rect 454404 131474 455004 131476
rect 490404 131474 491004 131476
rect 526404 131474 527004 131476
rect 562404 131474 563004 131476
rect 588080 131474 588680 131476
rect -2916 128476 -2316 128478
rect 18804 128476 19404 128478
rect 54804 128476 55404 128478
rect 90804 128476 91404 128478
rect 126804 128476 127404 128478
rect 162804 128476 163404 128478
rect 198804 128476 199404 128478
rect 234804 128476 235404 128478
rect 270804 128476 271404 128478
rect 306804 128476 307404 128478
rect 342804 128476 343404 128478
rect 378804 128476 379404 128478
rect 414804 128476 415404 128478
rect 450804 128476 451404 128478
rect 486804 128476 487404 128478
rect 522804 128476 523404 128478
rect 558804 128476 559404 128478
rect 586240 128476 586840 128478
rect -2916 128454 586840 128476
rect -2916 128218 -2734 128454
rect -2498 128218 18986 128454
rect 19222 128218 54986 128454
rect 55222 128218 90986 128454
rect 91222 128218 126986 128454
rect 127222 128218 162986 128454
rect 163222 128218 198986 128454
rect 199222 128218 234986 128454
rect 235222 128218 270986 128454
rect 271222 128218 306986 128454
rect 307222 128218 342986 128454
rect 343222 128218 378986 128454
rect 379222 128218 414986 128454
rect 415222 128218 450986 128454
rect 451222 128218 486986 128454
rect 487222 128218 522986 128454
rect 523222 128218 558986 128454
rect 559222 128218 586422 128454
rect 586658 128218 586840 128454
rect -2916 128134 586840 128218
rect -2916 127898 -2734 128134
rect -2498 127898 18986 128134
rect 19222 127898 54986 128134
rect 55222 127898 90986 128134
rect 91222 127898 126986 128134
rect 127222 127898 162986 128134
rect 163222 127898 198986 128134
rect 199222 127898 234986 128134
rect 235222 127898 270986 128134
rect 271222 127898 306986 128134
rect 307222 127898 342986 128134
rect 343222 127898 378986 128134
rect 379222 127898 414986 128134
rect 415222 127898 450986 128134
rect 451222 127898 486986 128134
rect 487222 127898 522986 128134
rect 523222 127898 558986 128134
rect 559222 127898 586422 128134
rect 586658 127898 586840 128134
rect -2916 127876 586840 127898
rect -2916 127874 -2316 127876
rect 18804 127874 19404 127876
rect 54804 127874 55404 127876
rect 90804 127874 91404 127876
rect 126804 127874 127404 127876
rect 162804 127874 163404 127876
rect 198804 127874 199404 127876
rect 234804 127874 235404 127876
rect 270804 127874 271404 127876
rect 306804 127874 307404 127876
rect 342804 127874 343404 127876
rect 378804 127874 379404 127876
rect 414804 127874 415404 127876
rect 450804 127874 451404 127876
rect 486804 127874 487404 127876
rect 522804 127874 523404 127876
rect 558804 127874 559404 127876
rect 586240 127874 586840 127876
rect -7516 121276 -6916 121278
rect 11604 121276 12204 121278
rect 47604 121276 48204 121278
rect 83604 121276 84204 121278
rect 119604 121276 120204 121278
rect 155604 121276 156204 121278
rect 191604 121276 192204 121278
rect 227604 121276 228204 121278
rect 263604 121276 264204 121278
rect 299604 121276 300204 121278
rect 335604 121276 336204 121278
rect 371604 121276 372204 121278
rect 407604 121276 408204 121278
rect 443604 121276 444204 121278
rect 479604 121276 480204 121278
rect 515604 121276 516204 121278
rect 551604 121276 552204 121278
rect 590840 121276 591440 121278
rect -8436 121254 592360 121276
rect -8436 121018 -7334 121254
rect -7098 121018 11786 121254
rect 12022 121018 47786 121254
rect 48022 121018 83786 121254
rect 84022 121018 119786 121254
rect 120022 121018 155786 121254
rect 156022 121018 191786 121254
rect 192022 121018 227786 121254
rect 228022 121018 263786 121254
rect 264022 121018 299786 121254
rect 300022 121018 335786 121254
rect 336022 121018 371786 121254
rect 372022 121018 407786 121254
rect 408022 121018 443786 121254
rect 444022 121018 479786 121254
rect 480022 121018 515786 121254
rect 516022 121018 551786 121254
rect 552022 121018 591022 121254
rect 591258 121018 592360 121254
rect -8436 120934 592360 121018
rect -8436 120698 -7334 120934
rect -7098 120698 11786 120934
rect 12022 120698 47786 120934
rect 48022 120698 83786 120934
rect 84022 120698 119786 120934
rect 120022 120698 155786 120934
rect 156022 120698 191786 120934
rect 192022 120698 227786 120934
rect 228022 120698 263786 120934
rect 264022 120698 299786 120934
rect 300022 120698 335786 120934
rect 336022 120698 371786 120934
rect 372022 120698 407786 120934
rect 408022 120698 443786 120934
rect 444022 120698 479786 120934
rect 480022 120698 515786 120934
rect 516022 120698 551786 120934
rect 552022 120698 591022 120934
rect 591258 120698 592360 120934
rect -8436 120676 592360 120698
rect -7516 120674 -6916 120676
rect 11604 120674 12204 120676
rect 47604 120674 48204 120676
rect 83604 120674 84204 120676
rect 119604 120674 120204 120676
rect 155604 120674 156204 120676
rect 191604 120674 192204 120676
rect 227604 120674 228204 120676
rect 263604 120674 264204 120676
rect 299604 120674 300204 120676
rect 335604 120674 336204 120676
rect 371604 120674 372204 120676
rect 407604 120674 408204 120676
rect 443604 120674 444204 120676
rect 479604 120674 480204 120676
rect 515604 120674 516204 120676
rect 551604 120674 552204 120676
rect 590840 120674 591440 120676
rect -5676 117676 -5076 117678
rect 8004 117676 8604 117678
rect 44004 117676 44604 117678
rect 80004 117676 80604 117678
rect 116004 117676 116604 117678
rect 152004 117676 152604 117678
rect 188004 117676 188604 117678
rect 224004 117676 224604 117678
rect 260004 117676 260604 117678
rect 296004 117676 296604 117678
rect 332004 117676 332604 117678
rect 368004 117676 368604 117678
rect 404004 117676 404604 117678
rect 440004 117676 440604 117678
rect 476004 117676 476604 117678
rect 512004 117676 512604 117678
rect 548004 117676 548604 117678
rect 589000 117676 589600 117678
rect -6596 117654 590520 117676
rect -6596 117418 -5494 117654
rect -5258 117418 8186 117654
rect 8422 117418 44186 117654
rect 44422 117418 80186 117654
rect 80422 117418 116186 117654
rect 116422 117418 152186 117654
rect 152422 117418 188186 117654
rect 188422 117418 224186 117654
rect 224422 117418 260186 117654
rect 260422 117418 296186 117654
rect 296422 117418 332186 117654
rect 332422 117418 368186 117654
rect 368422 117418 404186 117654
rect 404422 117418 440186 117654
rect 440422 117418 476186 117654
rect 476422 117418 512186 117654
rect 512422 117418 548186 117654
rect 548422 117418 589182 117654
rect 589418 117418 590520 117654
rect -6596 117334 590520 117418
rect -6596 117098 -5494 117334
rect -5258 117098 8186 117334
rect 8422 117098 44186 117334
rect 44422 117098 80186 117334
rect 80422 117098 116186 117334
rect 116422 117098 152186 117334
rect 152422 117098 188186 117334
rect 188422 117098 224186 117334
rect 224422 117098 260186 117334
rect 260422 117098 296186 117334
rect 296422 117098 332186 117334
rect 332422 117098 368186 117334
rect 368422 117098 404186 117334
rect 404422 117098 440186 117334
rect 440422 117098 476186 117334
rect 476422 117098 512186 117334
rect 512422 117098 548186 117334
rect 548422 117098 589182 117334
rect 589418 117098 590520 117334
rect -6596 117076 590520 117098
rect -5676 117074 -5076 117076
rect 8004 117074 8604 117076
rect 44004 117074 44604 117076
rect 80004 117074 80604 117076
rect 116004 117074 116604 117076
rect 152004 117074 152604 117076
rect 188004 117074 188604 117076
rect 224004 117074 224604 117076
rect 260004 117074 260604 117076
rect 296004 117074 296604 117076
rect 332004 117074 332604 117076
rect 368004 117074 368604 117076
rect 404004 117074 404604 117076
rect 440004 117074 440604 117076
rect 476004 117074 476604 117076
rect 512004 117074 512604 117076
rect 548004 117074 548604 117076
rect 589000 117074 589600 117076
rect -3836 114076 -3236 114078
rect 4404 114076 5004 114078
rect 40404 114076 41004 114078
rect 76404 114076 77004 114078
rect 112404 114076 113004 114078
rect 148404 114076 149004 114078
rect 184404 114076 185004 114078
rect 220404 114076 221004 114078
rect 256404 114076 257004 114078
rect 292404 114076 293004 114078
rect 328404 114076 329004 114078
rect 364404 114076 365004 114078
rect 400404 114076 401004 114078
rect 436404 114076 437004 114078
rect 472404 114076 473004 114078
rect 508404 114076 509004 114078
rect 544404 114076 545004 114078
rect 580404 114076 581004 114078
rect 587160 114076 587760 114078
rect -4756 114054 588680 114076
rect -4756 113818 -3654 114054
rect -3418 113818 4586 114054
rect 4822 113818 40586 114054
rect 40822 113818 76586 114054
rect 76822 113818 112586 114054
rect 112822 113818 148586 114054
rect 148822 113818 184586 114054
rect 184822 113818 220586 114054
rect 220822 113818 256586 114054
rect 256822 113818 292586 114054
rect 292822 113818 328586 114054
rect 328822 113818 364586 114054
rect 364822 113818 400586 114054
rect 400822 113818 436586 114054
rect 436822 113818 472586 114054
rect 472822 113818 508586 114054
rect 508822 113818 544586 114054
rect 544822 113818 580586 114054
rect 580822 113818 587342 114054
rect 587578 113818 588680 114054
rect -4756 113734 588680 113818
rect -4756 113498 -3654 113734
rect -3418 113498 4586 113734
rect 4822 113498 40586 113734
rect 40822 113498 76586 113734
rect 76822 113498 112586 113734
rect 112822 113498 148586 113734
rect 148822 113498 184586 113734
rect 184822 113498 220586 113734
rect 220822 113498 256586 113734
rect 256822 113498 292586 113734
rect 292822 113498 328586 113734
rect 328822 113498 364586 113734
rect 364822 113498 400586 113734
rect 400822 113498 436586 113734
rect 436822 113498 472586 113734
rect 472822 113498 508586 113734
rect 508822 113498 544586 113734
rect 544822 113498 580586 113734
rect 580822 113498 587342 113734
rect 587578 113498 588680 113734
rect -4756 113476 588680 113498
rect -3836 113474 -3236 113476
rect 4404 113474 5004 113476
rect 40404 113474 41004 113476
rect 76404 113474 77004 113476
rect 112404 113474 113004 113476
rect 148404 113474 149004 113476
rect 184404 113474 185004 113476
rect 220404 113474 221004 113476
rect 256404 113474 257004 113476
rect 292404 113474 293004 113476
rect 328404 113474 329004 113476
rect 364404 113474 365004 113476
rect 400404 113474 401004 113476
rect 436404 113474 437004 113476
rect 472404 113474 473004 113476
rect 508404 113474 509004 113476
rect 544404 113474 545004 113476
rect 580404 113474 581004 113476
rect 587160 113474 587760 113476
rect -1996 110476 -1396 110478
rect 804 110476 1404 110478
rect 36804 110476 37404 110478
rect 72804 110476 73404 110478
rect 108804 110476 109404 110478
rect 144804 110476 145404 110478
rect 180804 110476 181404 110478
rect 216804 110476 217404 110478
rect 252804 110476 253404 110478
rect 288804 110476 289404 110478
rect 324804 110476 325404 110478
rect 360804 110476 361404 110478
rect 396804 110476 397404 110478
rect 432804 110476 433404 110478
rect 468804 110476 469404 110478
rect 504804 110476 505404 110478
rect 540804 110476 541404 110478
rect 576804 110476 577404 110478
rect 585320 110476 585920 110478
rect -2916 110454 586840 110476
rect -2916 110218 -1814 110454
rect -1578 110218 986 110454
rect 1222 110218 36986 110454
rect 37222 110218 72986 110454
rect 73222 110218 108986 110454
rect 109222 110218 144986 110454
rect 145222 110218 180986 110454
rect 181222 110218 216986 110454
rect 217222 110218 252986 110454
rect 253222 110218 288986 110454
rect 289222 110218 324986 110454
rect 325222 110218 360986 110454
rect 361222 110218 396986 110454
rect 397222 110218 432986 110454
rect 433222 110218 468986 110454
rect 469222 110218 504986 110454
rect 505222 110218 540986 110454
rect 541222 110218 576986 110454
rect 577222 110218 585502 110454
rect 585738 110218 586840 110454
rect -2916 110134 586840 110218
rect -2916 109898 -1814 110134
rect -1578 109898 986 110134
rect 1222 109898 36986 110134
rect 37222 109898 72986 110134
rect 73222 109898 108986 110134
rect 109222 109898 144986 110134
rect 145222 109898 180986 110134
rect 181222 109898 216986 110134
rect 217222 109898 252986 110134
rect 253222 109898 288986 110134
rect 289222 109898 324986 110134
rect 325222 109898 360986 110134
rect 361222 109898 396986 110134
rect 397222 109898 432986 110134
rect 433222 109898 468986 110134
rect 469222 109898 504986 110134
rect 505222 109898 540986 110134
rect 541222 109898 576986 110134
rect 577222 109898 585502 110134
rect 585738 109898 586840 110134
rect -2916 109876 586840 109898
rect -1996 109874 -1396 109876
rect 804 109874 1404 109876
rect 36804 109874 37404 109876
rect 72804 109874 73404 109876
rect 108804 109874 109404 109876
rect 144804 109874 145404 109876
rect 180804 109874 181404 109876
rect 216804 109874 217404 109876
rect 252804 109874 253404 109876
rect 288804 109874 289404 109876
rect 324804 109874 325404 109876
rect 360804 109874 361404 109876
rect 396804 109874 397404 109876
rect 432804 109874 433404 109876
rect 468804 109874 469404 109876
rect 504804 109874 505404 109876
rect 540804 109874 541404 109876
rect 576804 109874 577404 109876
rect 585320 109874 585920 109876
rect -8436 103276 -7836 103278
rect 29604 103276 30204 103278
rect 65604 103276 66204 103278
rect 101604 103276 102204 103278
rect 137604 103276 138204 103278
rect 173604 103276 174204 103278
rect 209604 103276 210204 103278
rect 245604 103276 246204 103278
rect 281604 103276 282204 103278
rect 317604 103276 318204 103278
rect 353604 103276 354204 103278
rect 389604 103276 390204 103278
rect 425604 103276 426204 103278
rect 461604 103276 462204 103278
rect 497604 103276 498204 103278
rect 533604 103276 534204 103278
rect 569604 103276 570204 103278
rect 591760 103276 592360 103278
rect -8436 103254 592360 103276
rect -8436 103018 -8254 103254
rect -8018 103018 29786 103254
rect 30022 103018 65786 103254
rect 66022 103018 101786 103254
rect 102022 103018 137786 103254
rect 138022 103018 173786 103254
rect 174022 103018 209786 103254
rect 210022 103018 245786 103254
rect 246022 103018 281786 103254
rect 282022 103018 317786 103254
rect 318022 103018 353786 103254
rect 354022 103018 389786 103254
rect 390022 103018 425786 103254
rect 426022 103018 461786 103254
rect 462022 103018 497786 103254
rect 498022 103018 533786 103254
rect 534022 103018 569786 103254
rect 570022 103018 591942 103254
rect 592178 103018 592360 103254
rect -8436 102934 592360 103018
rect -8436 102698 -8254 102934
rect -8018 102698 29786 102934
rect 30022 102698 65786 102934
rect 66022 102698 101786 102934
rect 102022 102698 137786 102934
rect 138022 102698 173786 102934
rect 174022 102698 209786 102934
rect 210022 102698 245786 102934
rect 246022 102698 281786 102934
rect 282022 102698 317786 102934
rect 318022 102698 353786 102934
rect 354022 102698 389786 102934
rect 390022 102698 425786 102934
rect 426022 102698 461786 102934
rect 462022 102698 497786 102934
rect 498022 102698 533786 102934
rect 534022 102698 569786 102934
rect 570022 102698 591942 102934
rect 592178 102698 592360 102934
rect -8436 102676 592360 102698
rect -8436 102674 -7836 102676
rect 29604 102674 30204 102676
rect 65604 102674 66204 102676
rect 101604 102674 102204 102676
rect 137604 102674 138204 102676
rect 173604 102674 174204 102676
rect 209604 102674 210204 102676
rect 245604 102674 246204 102676
rect 281604 102674 282204 102676
rect 317604 102674 318204 102676
rect 353604 102674 354204 102676
rect 389604 102674 390204 102676
rect 425604 102674 426204 102676
rect 461604 102674 462204 102676
rect 497604 102674 498204 102676
rect 533604 102674 534204 102676
rect 569604 102674 570204 102676
rect 591760 102674 592360 102676
rect -6596 99676 -5996 99678
rect 26004 99676 26604 99678
rect 62004 99676 62604 99678
rect 98004 99676 98604 99678
rect 134004 99676 134604 99678
rect 170004 99676 170604 99678
rect 206004 99676 206604 99678
rect 242004 99676 242604 99678
rect 278004 99676 278604 99678
rect 314004 99676 314604 99678
rect 350004 99676 350604 99678
rect 386004 99676 386604 99678
rect 422004 99676 422604 99678
rect 458004 99676 458604 99678
rect 494004 99676 494604 99678
rect 530004 99676 530604 99678
rect 566004 99676 566604 99678
rect 589920 99676 590520 99678
rect -6596 99654 590520 99676
rect -6596 99418 -6414 99654
rect -6178 99418 26186 99654
rect 26422 99418 62186 99654
rect 62422 99418 98186 99654
rect 98422 99418 134186 99654
rect 134422 99418 170186 99654
rect 170422 99418 206186 99654
rect 206422 99418 242186 99654
rect 242422 99418 278186 99654
rect 278422 99418 314186 99654
rect 314422 99418 350186 99654
rect 350422 99418 386186 99654
rect 386422 99418 422186 99654
rect 422422 99418 458186 99654
rect 458422 99418 494186 99654
rect 494422 99418 530186 99654
rect 530422 99418 566186 99654
rect 566422 99418 590102 99654
rect 590338 99418 590520 99654
rect -6596 99334 590520 99418
rect -6596 99098 -6414 99334
rect -6178 99098 26186 99334
rect 26422 99098 62186 99334
rect 62422 99098 98186 99334
rect 98422 99098 134186 99334
rect 134422 99098 170186 99334
rect 170422 99098 206186 99334
rect 206422 99098 242186 99334
rect 242422 99098 278186 99334
rect 278422 99098 314186 99334
rect 314422 99098 350186 99334
rect 350422 99098 386186 99334
rect 386422 99098 422186 99334
rect 422422 99098 458186 99334
rect 458422 99098 494186 99334
rect 494422 99098 530186 99334
rect 530422 99098 566186 99334
rect 566422 99098 590102 99334
rect 590338 99098 590520 99334
rect -6596 99076 590520 99098
rect -6596 99074 -5996 99076
rect 26004 99074 26604 99076
rect 62004 99074 62604 99076
rect 98004 99074 98604 99076
rect 134004 99074 134604 99076
rect 170004 99074 170604 99076
rect 206004 99074 206604 99076
rect 242004 99074 242604 99076
rect 278004 99074 278604 99076
rect 314004 99074 314604 99076
rect 350004 99074 350604 99076
rect 386004 99074 386604 99076
rect 422004 99074 422604 99076
rect 458004 99074 458604 99076
rect 494004 99074 494604 99076
rect 530004 99074 530604 99076
rect 566004 99074 566604 99076
rect 589920 99074 590520 99076
rect -4756 96076 -4156 96078
rect 22404 96076 23004 96078
rect 58404 96076 59004 96078
rect 94404 96076 95004 96078
rect 130404 96076 131004 96078
rect 166404 96076 167004 96078
rect 202404 96076 203004 96078
rect 238404 96076 239004 96078
rect 274404 96076 275004 96078
rect 310404 96076 311004 96078
rect 346404 96076 347004 96078
rect 382404 96076 383004 96078
rect 418404 96076 419004 96078
rect 454404 96076 455004 96078
rect 490404 96076 491004 96078
rect 526404 96076 527004 96078
rect 562404 96076 563004 96078
rect 588080 96076 588680 96078
rect -4756 96054 588680 96076
rect -4756 95818 -4574 96054
rect -4338 95818 22586 96054
rect 22822 95818 58586 96054
rect 58822 95818 94586 96054
rect 94822 95818 130586 96054
rect 130822 95818 166586 96054
rect 166822 95818 202586 96054
rect 202822 95818 238586 96054
rect 238822 95818 274586 96054
rect 274822 95818 310586 96054
rect 310822 95818 346586 96054
rect 346822 95818 382586 96054
rect 382822 95818 418586 96054
rect 418822 95818 454586 96054
rect 454822 95818 490586 96054
rect 490822 95818 526586 96054
rect 526822 95818 562586 96054
rect 562822 95818 588262 96054
rect 588498 95818 588680 96054
rect -4756 95734 588680 95818
rect -4756 95498 -4574 95734
rect -4338 95498 22586 95734
rect 22822 95498 58586 95734
rect 58822 95498 94586 95734
rect 94822 95498 130586 95734
rect 130822 95498 166586 95734
rect 166822 95498 202586 95734
rect 202822 95498 238586 95734
rect 238822 95498 274586 95734
rect 274822 95498 310586 95734
rect 310822 95498 346586 95734
rect 346822 95498 382586 95734
rect 382822 95498 418586 95734
rect 418822 95498 454586 95734
rect 454822 95498 490586 95734
rect 490822 95498 526586 95734
rect 526822 95498 562586 95734
rect 562822 95498 588262 95734
rect 588498 95498 588680 95734
rect -4756 95476 588680 95498
rect -4756 95474 -4156 95476
rect 22404 95474 23004 95476
rect 58404 95474 59004 95476
rect 94404 95474 95004 95476
rect 130404 95474 131004 95476
rect 166404 95474 167004 95476
rect 202404 95474 203004 95476
rect 238404 95474 239004 95476
rect 274404 95474 275004 95476
rect 310404 95474 311004 95476
rect 346404 95474 347004 95476
rect 382404 95474 383004 95476
rect 418404 95474 419004 95476
rect 454404 95474 455004 95476
rect 490404 95474 491004 95476
rect 526404 95474 527004 95476
rect 562404 95474 563004 95476
rect 588080 95474 588680 95476
rect -2916 92476 -2316 92478
rect 18804 92476 19404 92478
rect 54804 92476 55404 92478
rect 90804 92476 91404 92478
rect 126804 92476 127404 92478
rect 162804 92476 163404 92478
rect 198804 92476 199404 92478
rect 234804 92476 235404 92478
rect 270804 92476 271404 92478
rect 306804 92476 307404 92478
rect 342804 92476 343404 92478
rect 378804 92476 379404 92478
rect 414804 92476 415404 92478
rect 450804 92476 451404 92478
rect 486804 92476 487404 92478
rect 522804 92476 523404 92478
rect 558804 92476 559404 92478
rect 586240 92476 586840 92478
rect -2916 92454 586840 92476
rect -2916 92218 -2734 92454
rect -2498 92218 18986 92454
rect 19222 92218 54986 92454
rect 55222 92218 90986 92454
rect 91222 92218 126986 92454
rect 127222 92218 162986 92454
rect 163222 92218 198986 92454
rect 199222 92218 234986 92454
rect 235222 92218 270986 92454
rect 271222 92218 306986 92454
rect 307222 92218 342986 92454
rect 343222 92218 378986 92454
rect 379222 92218 414986 92454
rect 415222 92218 450986 92454
rect 451222 92218 486986 92454
rect 487222 92218 522986 92454
rect 523222 92218 558986 92454
rect 559222 92218 586422 92454
rect 586658 92218 586840 92454
rect -2916 92134 586840 92218
rect -2916 91898 -2734 92134
rect -2498 91898 18986 92134
rect 19222 91898 54986 92134
rect 55222 91898 90986 92134
rect 91222 91898 126986 92134
rect 127222 91898 162986 92134
rect 163222 91898 198986 92134
rect 199222 91898 234986 92134
rect 235222 91898 270986 92134
rect 271222 91898 306986 92134
rect 307222 91898 342986 92134
rect 343222 91898 378986 92134
rect 379222 91898 414986 92134
rect 415222 91898 450986 92134
rect 451222 91898 486986 92134
rect 487222 91898 522986 92134
rect 523222 91898 558986 92134
rect 559222 91898 586422 92134
rect 586658 91898 586840 92134
rect -2916 91876 586840 91898
rect -2916 91874 -2316 91876
rect 18804 91874 19404 91876
rect 54804 91874 55404 91876
rect 90804 91874 91404 91876
rect 126804 91874 127404 91876
rect 162804 91874 163404 91876
rect 198804 91874 199404 91876
rect 234804 91874 235404 91876
rect 270804 91874 271404 91876
rect 306804 91874 307404 91876
rect 342804 91874 343404 91876
rect 378804 91874 379404 91876
rect 414804 91874 415404 91876
rect 450804 91874 451404 91876
rect 486804 91874 487404 91876
rect 522804 91874 523404 91876
rect 558804 91874 559404 91876
rect 586240 91874 586840 91876
rect -7516 85276 -6916 85278
rect 11604 85276 12204 85278
rect 47604 85276 48204 85278
rect 83604 85276 84204 85278
rect 119604 85276 120204 85278
rect 155604 85276 156204 85278
rect 191604 85276 192204 85278
rect 227604 85276 228204 85278
rect 263604 85276 264204 85278
rect 299604 85276 300204 85278
rect 335604 85276 336204 85278
rect 371604 85276 372204 85278
rect 407604 85276 408204 85278
rect 443604 85276 444204 85278
rect 479604 85276 480204 85278
rect 515604 85276 516204 85278
rect 551604 85276 552204 85278
rect 590840 85276 591440 85278
rect -8436 85254 592360 85276
rect -8436 85018 -7334 85254
rect -7098 85018 11786 85254
rect 12022 85018 47786 85254
rect 48022 85018 83786 85254
rect 84022 85018 119786 85254
rect 120022 85018 155786 85254
rect 156022 85018 191786 85254
rect 192022 85018 227786 85254
rect 228022 85018 263786 85254
rect 264022 85018 299786 85254
rect 300022 85018 335786 85254
rect 336022 85018 371786 85254
rect 372022 85018 407786 85254
rect 408022 85018 443786 85254
rect 444022 85018 479786 85254
rect 480022 85018 515786 85254
rect 516022 85018 551786 85254
rect 552022 85018 591022 85254
rect 591258 85018 592360 85254
rect -8436 84934 592360 85018
rect -8436 84698 -7334 84934
rect -7098 84698 11786 84934
rect 12022 84698 47786 84934
rect 48022 84698 83786 84934
rect 84022 84698 119786 84934
rect 120022 84698 155786 84934
rect 156022 84698 191786 84934
rect 192022 84698 227786 84934
rect 228022 84698 263786 84934
rect 264022 84698 299786 84934
rect 300022 84698 335786 84934
rect 336022 84698 371786 84934
rect 372022 84698 407786 84934
rect 408022 84698 443786 84934
rect 444022 84698 479786 84934
rect 480022 84698 515786 84934
rect 516022 84698 551786 84934
rect 552022 84698 591022 84934
rect 591258 84698 592360 84934
rect -8436 84676 592360 84698
rect -7516 84674 -6916 84676
rect 11604 84674 12204 84676
rect 47604 84674 48204 84676
rect 83604 84674 84204 84676
rect 119604 84674 120204 84676
rect 155604 84674 156204 84676
rect 191604 84674 192204 84676
rect 227604 84674 228204 84676
rect 263604 84674 264204 84676
rect 299604 84674 300204 84676
rect 335604 84674 336204 84676
rect 371604 84674 372204 84676
rect 407604 84674 408204 84676
rect 443604 84674 444204 84676
rect 479604 84674 480204 84676
rect 515604 84674 516204 84676
rect 551604 84674 552204 84676
rect 590840 84674 591440 84676
rect -5676 81676 -5076 81678
rect 8004 81676 8604 81678
rect 44004 81676 44604 81678
rect 80004 81676 80604 81678
rect 116004 81676 116604 81678
rect 152004 81676 152604 81678
rect 188004 81676 188604 81678
rect 224004 81676 224604 81678
rect 260004 81676 260604 81678
rect 296004 81676 296604 81678
rect 332004 81676 332604 81678
rect 368004 81676 368604 81678
rect 404004 81676 404604 81678
rect 440004 81676 440604 81678
rect 476004 81676 476604 81678
rect 512004 81676 512604 81678
rect 548004 81676 548604 81678
rect 589000 81676 589600 81678
rect -6596 81654 590520 81676
rect -6596 81418 -5494 81654
rect -5258 81418 8186 81654
rect 8422 81418 44186 81654
rect 44422 81418 80186 81654
rect 80422 81418 116186 81654
rect 116422 81418 152186 81654
rect 152422 81418 188186 81654
rect 188422 81418 224186 81654
rect 224422 81418 260186 81654
rect 260422 81418 296186 81654
rect 296422 81418 332186 81654
rect 332422 81418 368186 81654
rect 368422 81418 404186 81654
rect 404422 81418 440186 81654
rect 440422 81418 476186 81654
rect 476422 81418 512186 81654
rect 512422 81418 548186 81654
rect 548422 81418 589182 81654
rect 589418 81418 590520 81654
rect -6596 81334 590520 81418
rect -6596 81098 -5494 81334
rect -5258 81098 8186 81334
rect 8422 81098 44186 81334
rect 44422 81098 80186 81334
rect 80422 81098 116186 81334
rect 116422 81098 152186 81334
rect 152422 81098 188186 81334
rect 188422 81098 224186 81334
rect 224422 81098 260186 81334
rect 260422 81098 296186 81334
rect 296422 81098 332186 81334
rect 332422 81098 368186 81334
rect 368422 81098 404186 81334
rect 404422 81098 440186 81334
rect 440422 81098 476186 81334
rect 476422 81098 512186 81334
rect 512422 81098 548186 81334
rect 548422 81098 589182 81334
rect 589418 81098 590520 81334
rect -6596 81076 590520 81098
rect -5676 81074 -5076 81076
rect 8004 81074 8604 81076
rect 44004 81074 44604 81076
rect 80004 81074 80604 81076
rect 116004 81074 116604 81076
rect 152004 81074 152604 81076
rect 188004 81074 188604 81076
rect 224004 81074 224604 81076
rect 260004 81074 260604 81076
rect 296004 81074 296604 81076
rect 332004 81074 332604 81076
rect 368004 81074 368604 81076
rect 404004 81074 404604 81076
rect 440004 81074 440604 81076
rect 476004 81074 476604 81076
rect 512004 81074 512604 81076
rect 548004 81074 548604 81076
rect 589000 81074 589600 81076
rect -3836 78076 -3236 78078
rect 4404 78076 5004 78078
rect 40404 78076 41004 78078
rect 76404 78076 77004 78078
rect 112404 78076 113004 78078
rect 148404 78076 149004 78078
rect 184404 78076 185004 78078
rect 220404 78076 221004 78078
rect 256404 78076 257004 78078
rect 292404 78076 293004 78078
rect 328404 78076 329004 78078
rect 364404 78076 365004 78078
rect 400404 78076 401004 78078
rect 436404 78076 437004 78078
rect 472404 78076 473004 78078
rect 508404 78076 509004 78078
rect 544404 78076 545004 78078
rect 580404 78076 581004 78078
rect 587160 78076 587760 78078
rect -4756 78054 588680 78076
rect -4756 77818 -3654 78054
rect -3418 77818 4586 78054
rect 4822 77818 40586 78054
rect 40822 77818 76586 78054
rect 76822 77818 112586 78054
rect 112822 77818 148586 78054
rect 148822 77818 184586 78054
rect 184822 77818 220586 78054
rect 220822 77818 256586 78054
rect 256822 77818 292586 78054
rect 292822 77818 328586 78054
rect 328822 77818 364586 78054
rect 364822 77818 400586 78054
rect 400822 77818 436586 78054
rect 436822 77818 472586 78054
rect 472822 77818 508586 78054
rect 508822 77818 544586 78054
rect 544822 77818 580586 78054
rect 580822 77818 587342 78054
rect 587578 77818 588680 78054
rect -4756 77734 588680 77818
rect -4756 77498 -3654 77734
rect -3418 77498 4586 77734
rect 4822 77498 40586 77734
rect 40822 77498 76586 77734
rect 76822 77498 112586 77734
rect 112822 77498 148586 77734
rect 148822 77498 184586 77734
rect 184822 77498 220586 77734
rect 220822 77498 256586 77734
rect 256822 77498 292586 77734
rect 292822 77498 328586 77734
rect 328822 77498 364586 77734
rect 364822 77498 400586 77734
rect 400822 77498 436586 77734
rect 436822 77498 472586 77734
rect 472822 77498 508586 77734
rect 508822 77498 544586 77734
rect 544822 77498 580586 77734
rect 580822 77498 587342 77734
rect 587578 77498 588680 77734
rect -4756 77476 588680 77498
rect -3836 77474 -3236 77476
rect 4404 77474 5004 77476
rect 40404 77474 41004 77476
rect 76404 77474 77004 77476
rect 112404 77474 113004 77476
rect 148404 77474 149004 77476
rect 184404 77474 185004 77476
rect 220404 77474 221004 77476
rect 256404 77474 257004 77476
rect 292404 77474 293004 77476
rect 328404 77474 329004 77476
rect 364404 77474 365004 77476
rect 400404 77474 401004 77476
rect 436404 77474 437004 77476
rect 472404 77474 473004 77476
rect 508404 77474 509004 77476
rect 544404 77474 545004 77476
rect 580404 77474 581004 77476
rect 587160 77474 587760 77476
rect -1996 74476 -1396 74478
rect 804 74476 1404 74478
rect 36804 74476 37404 74478
rect 72804 74476 73404 74478
rect 108804 74476 109404 74478
rect 144804 74476 145404 74478
rect 180804 74476 181404 74478
rect 216804 74476 217404 74478
rect 252804 74476 253404 74478
rect 288804 74476 289404 74478
rect 324804 74476 325404 74478
rect 360804 74476 361404 74478
rect 396804 74476 397404 74478
rect 432804 74476 433404 74478
rect 468804 74476 469404 74478
rect 504804 74476 505404 74478
rect 540804 74476 541404 74478
rect 576804 74476 577404 74478
rect 585320 74476 585920 74478
rect -2916 74454 586840 74476
rect -2916 74218 -1814 74454
rect -1578 74218 986 74454
rect 1222 74218 36986 74454
rect 37222 74218 72986 74454
rect 73222 74218 108986 74454
rect 109222 74218 144986 74454
rect 145222 74218 180986 74454
rect 181222 74218 216986 74454
rect 217222 74218 252986 74454
rect 253222 74218 288986 74454
rect 289222 74218 324986 74454
rect 325222 74218 360986 74454
rect 361222 74218 396986 74454
rect 397222 74218 432986 74454
rect 433222 74218 468986 74454
rect 469222 74218 504986 74454
rect 505222 74218 540986 74454
rect 541222 74218 576986 74454
rect 577222 74218 585502 74454
rect 585738 74218 586840 74454
rect -2916 74134 586840 74218
rect -2916 73898 -1814 74134
rect -1578 73898 986 74134
rect 1222 73898 36986 74134
rect 37222 73898 72986 74134
rect 73222 73898 108986 74134
rect 109222 73898 144986 74134
rect 145222 73898 180986 74134
rect 181222 73898 216986 74134
rect 217222 73898 252986 74134
rect 253222 73898 288986 74134
rect 289222 73898 324986 74134
rect 325222 73898 360986 74134
rect 361222 73898 396986 74134
rect 397222 73898 432986 74134
rect 433222 73898 468986 74134
rect 469222 73898 504986 74134
rect 505222 73898 540986 74134
rect 541222 73898 576986 74134
rect 577222 73898 585502 74134
rect 585738 73898 586840 74134
rect -2916 73876 586840 73898
rect -1996 73874 -1396 73876
rect 804 73874 1404 73876
rect 36804 73874 37404 73876
rect 72804 73874 73404 73876
rect 108804 73874 109404 73876
rect 144804 73874 145404 73876
rect 180804 73874 181404 73876
rect 216804 73874 217404 73876
rect 252804 73874 253404 73876
rect 288804 73874 289404 73876
rect 324804 73874 325404 73876
rect 360804 73874 361404 73876
rect 396804 73874 397404 73876
rect 432804 73874 433404 73876
rect 468804 73874 469404 73876
rect 504804 73874 505404 73876
rect 540804 73874 541404 73876
rect 576804 73874 577404 73876
rect 585320 73874 585920 73876
rect -8436 67276 -7836 67278
rect 29604 67276 30204 67278
rect 65604 67276 66204 67278
rect 101604 67276 102204 67278
rect 137604 67276 138204 67278
rect 173604 67276 174204 67278
rect 209604 67276 210204 67278
rect 245604 67276 246204 67278
rect 281604 67276 282204 67278
rect 317604 67276 318204 67278
rect 353604 67276 354204 67278
rect 389604 67276 390204 67278
rect 425604 67276 426204 67278
rect 461604 67276 462204 67278
rect 497604 67276 498204 67278
rect 533604 67276 534204 67278
rect 569604 67276 570204 67278
rect 591760 67276 592360 67278
rect -8436 67254 592360 67276
rect -8436 67018 -8254 67254
rect -8018 67018 29786 67254
rect 30022 67018 65786 67254
rect 66022 67018 101786 67254
rect 102022 67018 137786 67254
rect 138022 67018 173786 67254
rect 174022 67018 209786 67254
rect 210022 67018 245786 67254
rect 246022 67018 281786 67254
rect 282022 67018 317786 67254
rect 318022 67018 353786 67254
rect 354022 67018 389786 67254
rect 390022 67018 425786 67254
rect 426022 67018 461786 67254
rect 462022 67018 497786 67254
rect 498022 67018 533786 67254
rect 534022 67018 569786 67254
rect 570022 67018 591942 67254
rect 592178 67018 592360 67254
rect -8436 66934 592360 67018
rect -8436 66698 -8254 66934
rect -8018 66698 29786 66934
rect 30022 66698 65786 66934
rect 66022 66698 101786 66934
rect 102022 66698 137786 66934
rect 138022 66698 173786 66934
rect 174022 66698 209786 66934
rect 210022 66698 245786 66934
rect 246022 66698 281786 66934
rect 282022 66698 317786 66934
rect 318022 66698 353786 66934
rect 354022 66698 389786 66934
rect 390022 66698 425786 66934
rect 426022 66698 461786 66934
rect 462022 66698 497786 66934
rect 498022 66698 533786 66934
rect 534022 66698 569786 66934
rect 570022 66698 591942 66934
rect 592178 66698 592360 66934
rect -8436 66676 592360 66698
rect -8436 66674 -7836 66676
rect 29604 66674 30204 66676
rect 65604 66674 66204 66676
rect 101604 66674 102204 66676
rect 137604 66674 138204 66676
rect 173604 66674 174204 66676
rect 209604 66674 210204 66676
rect 245604 66674 246204 66676
rect 281604 66674 282204 66676
rect 317604 66674 318204 66676
rect 353604 66674 354204 66676
rect 389604 66674 390204 66676
rect 425604 66674 426204 66676
rect 461604 66674 462204 66676
rect 497604 66674 498204 66676
rect 533604 66674 534204 66676
rect 569604 66674 570204 66676
rect 591760 66674 592360 66676
rect -6596 63676 -5996 63678
rect 26004 63676 26604 63678
rect 62004 63676 62604 63678
rect 98004 63676 98604 63678
rect 134004 63676 134604 63678
rect 170004 63676 170604 63678
rect 206004 63676 206604 63678
rect 242004 63676 242604 63678
rect 278004 63676 278604 63678
rect 314004 63676 314604 63678
rect 350004 63676 350604 63678
rect 386004 63676 386604 63678
rect 422004 63676 422604 63678
rect 458004 63676 458604 63678
rect 494004 63676 494604 63678
rect 530004 63676 530604 63678
rect 566004 63676 566604 63678
rect 589920 63676 590520 63678
rect -6596 63654 590520 63676
rect -6596 63418 -6414 63654
rect -6178 63418 26186 63654
rect 26422 63418 62186 63654
rect 62422 63418 98186 63654
rect 98422 63418 134186 63654
rect 134422 63418 170186 63654
rect 170422 63418 206186 63654
rect 206422 63418 242186 63654
rect 242422 63418 278186 63654
rect 278422 63418 314186 63654
rect 314422 63418 350186 63654
rect 350422 63418 386186 63654
rect 386422 63418 422186 63654
rect 422422 63418 458186 63654
rect 458422 63418 494186 63654
rect 494422 63418 530186 63654
rect 530422 63418 566186 63654
rect 566422 63418 590102 63654
rect 590338 63418 590520 63654
rect -6596 63334 590520 63418
rect -6596 63098 -6414 63334
rect -6178 63098 26186 63334
rect 26422 63098 62186 63334
rect 62422 63098 98186 63334
rect 98422 63098 134186 63334
rect 134422 63098 170186 63334
rect 170422 63098 206186 63334
rect 206422 63098 242186 63334
rect 242422 63098 278186 63334
rect 278422 63098 314186 63334
rect 314422 63098 350186 63334
rect 350422 63098 386186 63334
rect 386422 63098 422186 63334
rect 422422 63098 458186 63334
rect 458422 63098 494186 63334
rect 494422 63098 530186 63334
rect 530422 63098 566186 63334
rect 566422 63098 590102 63334
rect 590338 63098 590520 63334
rect -6596 63076 590520 63098
rect -6596 63074 -5996 63076
rect 26004 63074 26604 63076
rect 62004 63074 62604 63076
rect 98004 63074 98604 63076
rect 134004 63074 134604 63076
rect 170004 63074 170604 63076
rect 206004 63074 206604 63076
rect 242004 63074 242604 63076
rect 278004 63074 278604 63076
rect 314004 63074 314604 63076
rect 350004 63074 350604 63076
rect 386004 63074 386604 63076
rect 422004 63074 422604 63076
rect 458004 63074 458604 63076
rect 494004 63074 494604 63076
rect 530004 63074 530604 63076
rect 566004 63074 566604 63076
rect 589920 63074 590520 63076
rect -4756 60076 -4156 60078
rect 22404 60076 23004 60078
rect 58404 60076 59004 60078
rect 94404 60076 95004 60078
rect 130404 60076 131004 60078
rect 166404 60076 167004 60078
rect 202404 60076 203004 60078
rect 238404 60076 239004 60078
rect 274404 60076 275004 60078
rect 310404 60076 311004 60078
rect 346404 60076 347004 60078
rect 382404 60076 383004 60078
rect 418404 60076 419004 60078
rect 454404 60076 455004 60078
rect 490404 60076 491004 60078
rect 526404 60076 527004 60078
rect 562404 60076 563004 60078
rect 588080 60076 588680 60078
rect -4756 60054 588680 60076
rect -4756 59818 -4574 60054
rect -4338 59818 22586 60054
rect 22822 59818 58586 60054
rect 58822 59818 94586 60054
rect 94822 59818 130586 60054
rect 130822 59818 166586 60054
rect 166822 59818 202586 60054
rect 202822 59818 238586 60054
rect 238822 59818 274586 60054
rect 274822 59818 310586 60054
rect 310822 59818 346586 60054
rect 346822 59818 382586 60054
rect 382822 59818 418586 60054
rect 418822 59818 454586 60054
rect 454822 59818 490586 60054
rect 490822 59818 526586 60054
rect 526822 59818 562586 60054
rect 562822 59818 588262 60054
rect 588498 59818 588680 60054
rect -4756 59734 588680 59818
rect -4756 59498 -4574 59734
rect -4338 59498 22586 59734
rect 22822 59498 58586 59734
rect 58822 59498 94586 59734
rect 94822 59498 130586 59734
rect 130822 59498 166586 59734
rect 166822 59498 202586 59734
rect 202822 59498 238586 59734
rect 238822 59498 274586 59734
rect 274822 59498 310586 59734
rect 310822 59498 346586 59734
rect 346822 59498 382586 59734
rect 382822 59498 418586 59734
rect 418822 59498 454586 59734
rect 454822 59498 490586 59734
rect 490822 59498 526586 59734
rect 526822 59498 562586 59734
rect 562822 59498 588262 59734
rect 588498 59498 588680 59734
rect -4756 59476 588680 59498
rect -4756 59474 -4156 59476
rect 22404 59474 23004 59476
rect 58404 59474 59004 59476
rect 94404 59474 95004 59476
rect 130404 59474 131004 59476
rect 166404 59474 167004 59476
rect 202404 59474 203004 59476
rect 238404 59474 239004 59476
rect 274404 59474 275004 59476
rect 310404 59474 311004 59476
rect 346404 59474 347004 59476
rect 382404 59474 383004 59476
rect 418404 59474 419004 59476
rect 454404 59474 455004 59476
rect 490404 59474 491004 59476
rect 526404 59474 527004 59476
rect 562404 59474 563004 59476
rect 588080 59474 588680 59476
rect -2916 56476 -2316 56478
rect 18804 56476 19404 56478
rect 54804 56476 55404 56478
rect 90804 56476 91404 56478
rect 126804 56476 127404 56478
rect 162804 56476 163404 56478
rect 198804 56476 199404 56478
rect 234804 56476 235404 56478
rect 270804 56476 271404 56478
rect 306804 56476 307404 56478
rect 342804 56476 343404 56478
rect 378804 56476 379404 56478
rect 414804 56476 415404 56478
rect 450804 56476 451404 56478
rect 486804 56476 487404 56478
rect 522804 56476 523404 56478
rect 558804 56476 559404 56478
rect 586240 56476 586840 56478
rect -2916 56454 586840 56476
rect -2916 56218 -2734 56454
rect -2498 56218 18986 56454
rect 19222 56218 54986 56454
rect 55222 56218 90986 56454
rect 91222 56218 126986 56454
rect 127222 56218 162986 56454
rect 163222 56218 198986 56454
rect 199222 56218 234986 56454
rect 235222 56218 270986 56454
rect 271222 56218 306986 56454
rect 307222 56218 342986 56454
rect 343222 56218 378986 56454
rect 379222 56218 414986 56454
rect 415222 56218 450986 56454
rect 451222 56218 486986 56454
rect 487222 56218 522986 56454
rect 523222 56218 558986 56454
rect 559222 56218 586422 56454
rect 586658 56218 586840 56454
rect -2916 56134 586840 56218
rect -2916 55898 -2734 56134
rect -2498 55898 18986 56134
rect 19222 55898 54986 56134
rect 55222 55898 90986 56134
rect 91222 55898 126986 56134
rect 127222 55898 162986 56134
rect 163222 55898 198986 56134
rect 199222 55898 234986 56134
rect 235222 55898 270986 56134
rect 271222 55898 306986 56134
rect 307222 55898 342986 56134
rect 343222 55898 378986 56134
rect 379222 55898 414986 56134
rect 415222 55898 450986 56134
rect 451222 55898 486986 56134
rect 487222 55898 522986 56134
rect 523222 55898 558986 56134
rect 559222 55898 586422 56134
rect 586658 55898 586840 56134
rect -2916 55876 586840 55898
rect -2916 55874 -2316 55876
rect 18804 55874 19404 55876
rect 54804 55874 55404 55876
rect 90804 55874 91404 55876
rect 126804 55874 127404 55876
rect 162804 55874 163404 55876
rect 198804 55874 199404 55876
rect 234804 55874 235404 55876
rect 270804 55874 271404 55876
rect 306804 55874 307404 55876
rect 342804 55874 343404 55876
rect 378804 55874 379404 55876
rect 414804 55874 415404 55876
rect 450804 55874 451404 55876
rect 486804 55874 487404 55876
rect 522804 55874 523404 55876
rect 558804 55874 559404 55876
rect 586240 55874 586840 55876
rect -7516 49276 -6916 49278
rect 11604 49276 12204 49278
rect 47604 49276 48204 49278
rect 83604 49276 84204 49278
rect 119604 49276 120204 49278
rect 155604 49276 156204 49278
rect 191604 49276 192204 49278
rect 227604 49276 228204 49278
rect 263604 49276 264204 49278
rect 299604 49276 300204 49278
rect 335604 49276 336204 49278
rect 371604 49276 372204 49278
rect 407604 49276 408204 49278
rect 443604 49276 444204 49278
rect 479604 49276 480204 49278
rect 515604 49276 516204 49278
rect 551604 49276 552204 49278
rect 590840 49276 591440 49278
rect -8436 49254 592360 49276
rect -8436 49018 -7334 49254
rect -7098 49018 11786 49254
rect 12022 49018 47786 49254
rect 48022 49018 83786 49254
rect 84022 49018 119786 49254
rect 120022 49018 155786 49254
rect 156022 49018 191786 49254
rect 192022 49018 227786 49254
rect 228022 49018 263786 49254
rect 264022 49018 299786 49254
rect 300022 49018 335786 49254
rect 336022 49018 371786 49254
rect 372022 49018 407786 49254
rect 408022 49018 443786 49254
rect 444022 49018 479786 49254
rect 480022 49018 515786 49254
rect 516022 49018 551786 49254
rect 552022 49018 591022 49254
rect 591258 49018 592360 49254
rect -8436 48934 592360 49018
rect -8436 48698 -7334 48934
rect -7098 48698 11786 48934
rect 12022 48698 47786 48934
rect 48022 48698 83786 48934
rect 84022 48698 119786 48934
rect 120022 48698 155786 48934
rect 156022 48698 191786 48934
rect 192022 48698 227786 48934
rect 228022 48698 263786 48934
rect 264022 48698 299786 48934
rect 300022 48698 335786 48934
rect 336022 48698 371786 48934
rect 372022 48698 407786 48934
rect 408022 48698 443786 48934
rect 444022 48698 479786 48934
rect 480022 48698 515786 48934
rect 516022 48698 551786 48934
rect 552022 48698 591022 48934
rect 591258 48698 592360 48934
rect -8436 48676 592360 48698
rect -7516 48674 -6916 48676
rect 11604 48674 12204 48676
rect 47604 48674 48204 48676
rect 83604 48674 84204 48676
rect 119604 48674 120204 48676
rect 155604 48674 156204 48676
rect 191604 48674 192204 48676
rect 227604 48674 228204 48676
rect 263604 48674 264204 48676
rect 299604 48674 300204 48676
rect 335604 48674 336204 48676
rect 371604 48674 372204 48676
rect 407604 48674 408204 48676
rect 443604 48674 444204 48676
rect 479604 48674 480204 48676
rect 515604 48674 516204 48676
rect 551604 48674 552204 48676
rect 590840 48674 591440 48676
rect -5676 45676 -5076 45678
rect 8004 45676 8604 45678
rect 44004 45676 44604 45678
rect 80004 45676 80604 45678
rect 116004 45676 116604 45678
rect 152004 45676 152604 45678
rect 188004 45676 188604 45678
rect 224004 45676 224604 45678
rect 260004 45676 260604 45678
rect 296004 45676 296604 45678
rect 332004 45676 332604 45678
rect 368004 45676 368604 45678
rect 404004 45676 404604 45678
rect 440004 45676 440604 45678
rect 476004 45676 476604 45678
rect 512004 45676 512604 45678
rect 548004 45676 548604 45678
rect 589000 45676 589600 45678
rect -6596 45654 590520 45676
rect -6596 45418 -5494 45654
rect -5258 45418 8186 45654
rect 8422 45418 44186 45654
rect 44422 45418 80186 45654
rect 80422 45418 116186 45654
rect 116422 45418 152186 45654
rect 152422 45418 188186 45654
rect 188422 45418 224186 45654
rect 224422 45418 260186 45654
rect 260422 45418 296186 45654
rect 296422 45418 332186 45654
rect 332422 45418 368186 45654
rect 368422 45418 404186 45654
rect 404422 45418 440186 45654
rect 440422 45418 476186 45654
rect 476422 45418 512186 45654
rect 512422 45418 548186 45654
rect 548422 45418 589182 45654
rect 589418 45418 590520 45654
rect -6596 45334 590520 45418
rect -6596 45098 -5494 45334
rect -5258 45098 8186 45334
rect 8422 45098 44186 45334
rect 44422 45098 80186 45334
rect 80422 45098 116186 45334
rect 116422 45098 152186 45334
rect 152422 45098 188186 45334
rect 188422 45098 224186 45334
rect 224422 45098 260186 45334
rect 260422 45098 296186 45334
rect 296422 45098 332186 45334
rect 332422 45098 368186 45334
rect 368422 45098 404186 45334
rect 404422 45098 440186 45334
rect 440422 45098 476186 45334
rect 476422 45098 512186 45334
rect 512422 45098 548186 45334
rect 548422 45098 589182 45334
rect 589418 45098 590520 45334
rect -6596 45076 590520 45098
rect -5676 45074 -5076 45076
rect 8004 45074 8604 45076
rect 44004 45074 44604 45076
rect 80004 45074 80604 45076
rect 116004 45074 116604 45076
rect 152004 45074 152604 45076
rect 188004 45074 188604 45076
rect 224004 45074 224604 45076
rect 260004 45074 260604 45076
rect 296004 45074 296604 45076
rect 332004 45074 332604 45076
rect 368004 45074 368604 45076
rect 404004 45074 404604 45076
rect 440004 45074 440604 45076
rect 476004 45074 476604 45076
rect 512004 45074 512604 45076
rect 548004 45074 548604 45076
rect 589000 45074 589600 45076
rect -3836 42076 -3236 42078
rect 4404 42076 5004 42078
rect 40404 42076 41004 42078
rect 76404 42076 77004 42078
rect 112404 42076 113004 42078
rect 148404 42076 149004 42078
rect 184404 42076 185004 42078
rect 220404 42076 221004 42078
rect 256404 42076 257004 42078
rect 292404 42076 293004 42078
rect 328404 42076 329004 42078
rect 364404 42076 365004 42078
rect 400404 42076 401004 42078
rect 436404 42076 437004 42078
rect 472404 42076 473004 42078
rect 508404 42076 509004 42078
rect 544404 42076 545004 42078
rect 580404 42076 581004 42078
rect 587160 42076 587760 42078
rect -4756 42054 588680 42076
rect -4756 41818 -3654 42054
rect -3418 41818 4586 42054
rect 4822 41818 40586 42054
rect 40822 41818 76586 42054
rect 76822 41818 112586 42054
rect 112822 41818 148586 42054
rect 148822 41818 184586 42054
rect 184822 41818 220586 42054
rect 220822 41818 256586 42054
rect 256822 41818 292586 42054
rect 292822 41818 328586 42054
rect 328822 41818 364586 42054
rect 364822 41818 400586 42054
rect 400822 41818 436586 42054
rect 436822 41818 472586 42054
rect 472822 41818 508586 42054
rect 508822 41818 544586 42054
rect 544822 41818 580586 42054
rect 580822 41818 587342 42054
rect 587578 41818 588680 42054
rect -4756 41734 588680 41818
rect -4756 41498 -3654 41734
rect -3418 41498 4586 41734
rect 4822 41498 40586 41734
rect 40822 41498 76586 41734
rect 76822 41498 112586 41734
rect 112822 41498 148586 41734
rect 148822 41498 184586 41734
rect 184822 41498 220586 41734
rect 220822 41498 256586 41734
rect 256822 41498 292586 41734
rect 292822 41498 328586 41734
rect 328822 41498 364586 41734
rect 364822 41498 400586 41734
rect 400822 41498 436586 41734
rect 436822 41498 472586 41734
rect 472822 41498 508586 41734
rect 508822 41498 544586 41734
rect 544822 41498 580586 41734
rect 580822 41498 587342 41734
rect 587578 41498 588680 41734
rect -4756 41476 588680 41498
rect -3836 41474 -3236 41476
rect 4404 41474 5004 41476
rect 40404 41474 41004 41476
rect 76404 41474 77004 41476
rect 112404 41474 113004 41476
rect 148404 41474 149004 41476
rect 184404 41474 185004 41476
rect 220404 41474 221004 41476
rect 256404 41474 257004 41476
rect 292404 41474 293004 41476
rect 328404 41474 329004 41476
rect 364404 41474 365004 41476
rect 400404 41474 401004 41476
rect 436404 41474 437004 41476
rect 472404 41474 473004 41476
rect 508404 41474 509004 41476
rect 544404 41474 545004 41476
rect 580404 41474 581004 41476
rect 587160 41474 587760 41476
rect -1996 38476 -1396 38478
rect 804 38476 1404 38478
rect 36804 38476 37404 38478
rect 72804 38476 73404 38478
rect 108804 38476 109404 38478
rect 144804 38476 145404 38478
rect 180804 38476 181404 38478
rect 216804 38476 217404 38478
rect 252804 38476 253404 38478
rect 288804 38476 289404 38478
rect 324804 38476 325404 38478
rect 360804 38476 361404 38478
rect 396804 38476 397404 38478
rect 432804 38476 433404 38478
rect 468804 38476 469404 38478
rect 504804 38476 505404 38478
rect 540804 38476 541404 38478
rect 576804 38476 577404 38478
rect 585320 38476 585920 38478
rect -2916 38454 586840 38476
rect -2916 38218 -1814 38454
rect -1578 38218 986 38454
rect 1222 38218 36986 38454
rect 37222 38218 72986 38454
rect 73222 38218 108986 38454
rect 109222 38218 144986 38454
rect 145222 38218 180986 38454
rect 181222 38218 216986 38454
rect 217222 38218 252986 38454
rect 253222 38218 288986 38454
rect 289222 38218 324986 38454
rect 325222 38218 360986 38454
rect 361222 38218 396986 38454
rect 397222 38218 432986 38454
rect 433222 38218 468986 38454
rect 469222 38218 504986 38454
rect 505222 38218 540986 38454
rect 541222 38218 576986 38454
rect 577222 38218 585502 38454
rect 585738 38218 586840 38454
rect -2916 38134 586840 38218
rect -2916 37898 -1814 38134
rect -1578 37898 986 38134
rect 1222 37898 36986 38134
rect 37222 37898 72986 38134
rect 73222 37898 108986 38134
rect 109222 37898 144986 38134
rect 145222 37898 180986 38134
rect 181222 37898 216986 38134
rect 217222 37898 252986 38134
rect 253222 37898 288986 38134
rect 289222 37898 324986 38134
rect 325222 37898 360986 38134
rect 361222 37898 396986 38134
rect 397222 37898 432986 38134
rect 433222 37898 468986 38134
rect 469222 37898 504986 38134
rect 505222 37898 540986 38134
rect 541222 37898 576986 38134
rect 577222 37898 585502 38134
rect 585738 37898 586840 38134
rect -2916 37876 586840 37898
rect -1996 37874 -1396 37876
rect 804 37874 1404 37876
rect 36804 37874 37404 37876
rect 72804 37874 73404 37876
rect 108804 37874 109404 37876
rect 144804 37874 145404 37876
rect 180804 37874 181404 37876
rect 216804 37874 217404 37876
rect 252804 37874 253404 37876
rect 288804 37874 289404 37876
rect 324804 37874 325404 37876
rect 360804 37874 361404 37876
rect 396804 37874 397404 37876
rect 432804 37874 433404 37876
rect 468804 37874 469404 37876
rect 504804 37874 505404 37876
rect 540804 37874 541404 37876
rect 576804 37874 577404 37876
rect 585320 37874 585920 37876
rect -8436 31276 -7836 31278
rect 29604 31276 30204 31278
rect 65604 31276 66204 31278
rect 101604 31276 102204 31278
rect 137604 31276 138204 31278
rect 173604 31276 174204 31278
rect 209604 31276 210204 31278
rect 245604 31276 246204 31278
rect 281604 31276 282204 31278
rect 317604 31276 318204 31278
rect 353604 31276 354204 31278
rect 389604 31276 390204 31278
rect 425604 31276 426204 31278
rect 461604 31276 462204 31278
rect 497604 31276 498204 31278
rect 533604 31276 534204 31278
rect 569604 31276 570204 31278
rect 591760 31276 592360 31278
rect -8436 31254 592360 31276
rect -8436 31018 -8254 31254
rect -8018 31018 29786 31254
rect 30022 31018 65786 31254
rect 66022 31018 101786 31254
rect 102022 31018 137786 31254
rect 138022 31018 173786 31254
rect 174022 31018 209786 31254
rect 210022 31018 245786 31254
rect 246022 31018 281786 31254
rect 282022 31018 317786 31254
rect 318022 31018 353786 31254
rect 354022 31018 389786 31254
rect 390022 31018 425786 31254
rect 426022 31018 461786 31254
rect 462022 31018 497786 31254
rect 498022 31018 533786 31254
rect 534022 31018 569786 31254
rect 570022 31018 591942 31254
rect 592178 31018 592360 31254
rect -8436 30934 592360 31018
rect -8436 30698 -8254 30934
rect -8018 30698 29786 30934
rect 30022 30698 65786 30934
rect 66022 30698 101786 30934
rect 102022 30698 137786 30934
rect 138022 30698 173786 30934
rect 174022 30698 209786 30934
rect 210022 30698 245786 30934
rect 246022 30698 281786 30934
rect 282022 30698 317786 30934
rect 318022 30698 353786 30934
rect 354022 30698 389786 30934
rect 390022 30698 425786 30934
rect 426022 30698 461786 30934
rect 462022 30698 497786 30934
rect 498022 30698 533786 30934
rect 534022 30698 569786 30934
rect 570022 30698 591942 30934
rect 592178 30698 592360 30934
rect -8436 30676 592360 30698
rect -8436 30674 -7836 30676
rect 29604 30674 30204 30676
rect 65604 30674 66204 30676
rect 101604 30674 102204 30676
rect 137604 30674 138204 30676
rect 173604 30674 174204 30676
rect 209604 30674 210204 30676
rect 245604 30674 246204 30676
rect 281604 30674 282204 30676
rect 317604 30674 318204 30676
rect 353604 30674 354204 30676
rect 389604 30674 390204 30676
rect 425604 30674 426204 30676
rect 461604 30674 462204 30676
rect 497604 30674 498204 30676
rect 533604 30674 534204 30676
rect 569604 30674 570204 30676
rect 591760 30674 592360 30676
rect -6596 27676 -5996 27678
rect 26004 27676 26604 27678
rect 62004 27676 62604 27678
rect 98004 27676 98604 27678
rect 134004 27676 134604 27678
rect 170004 27676 170604 27678
rect 206004 27676 206604 27678
rect 242004 27676 242604 27678
rect 278004 27676 278604 27678
rect 314004 27676 314604 27678
rect 350004 27676 350604 27678
rect 386004 27676 386604 27678
rect 422004 27676 422604 27678
rect 458004 27676 458604 27678
rect 494004 27676 494604 27678
rect 530004 27676 530604 27678
rect 566004 27676 566604 27678
rect 589920 27676 590520 27678
rect -6596 27654 590520 27676
rect -6596 27418 -6414 27654
rect -6178 27418 26186 27654
rect 26422 27418 62186 27654
rect 62422 27418 98186 27654
rect 98422 27418 134186 27654
rect 134422 27418 170186 27654
rect 170422 27418 206186 27654
rect 206422 27418 242186 27654
rect 242422 27418 278186 27654
rect 278422 27418 314186 27654
rect 314422 27418 350186 27654
rect 350422 27418 386186 27654
rect 386422 27418 422186 27654
rect 422422 27418 458186 27654
rect 458422 27418 494186 27654
rect 494422 27418 530186 27654
rect 530422 27418 566186 27654
rect 566422 27418 590102 27654
rect 590338 27418 590520 27654
rect -6596 27334 590520 27418
rect -6596 27098 -6414 27334
rect -6178 27098 26186 27334
rect 26422 27098 62186 27334
rect 62422 27098 98186 27334
rect 98422 27098 134186 27334
rect 134422 27098 170186 27334
rect 170422 27098 206186 27334
rect 206422 27098 242186 27334
rect 242422 27098 278186 27334
rect 278422 27098 314186 27334
rect 314422 27098 350186 27334
rect 350422 27098 386186 27334
rect 386422 27098 422186 27334
rect 422422 27098 458186 27334
rect 458422 27098 494186 27334
rect 494422 27098 530186 27334
rect 530422 27098 566186 27334
rect 566422 27098 590102 27334
rect 590338 27098 590520 27334
rect -6596 27076 590520 27098
rect -6596 27074 -5996 27076
rect 26004 27074 26604 27076
rect 62004 27074 62604 27076
rect 98004 27074 98604 27076
rect 134004 27074 134604 27076
rect 170004 27074 170604 27076
rect 206004 27074 206604 27076
rect 242004 27074 242604 27076
rect 278004 27074 278604 27076
rect 314004 27074 314604 27076
rect 350004 27074 350604 27076
rect 386004 27074 386604 27076
rect 422004 27074 422604 27076
rect 458004 27074 458604 27076
rect 494004 27074 494604 27076
rect 530004 27074 530604 27076
rect 566004 27074 566604 27076
rect 589920 27074 590520 27076
rect -4756 24076 -4156 24078
rect 22404 24076 23004 24078
rect 58404 24076 59004 24078
rect 94404 24076 95004 24078
rect 130404 24076 131004 24078
rect 166404 24076 167004 24078
rect 202404 24076 203004 24078
rect 238404 24076 239004 24078
rect 274404 24076 275004 24078
rect 310404 24076 311004 24078
rect 346404 24076 347004 24078
rect 382404 24076 383004 24078
rect 418404 24076 419004 24078
rect 454404 24076 455004 24078
rect 490404 24076 491004 24078
rect 526404 24076 527004 24078
rect 562404 24076 563004 24078
rect 588080 24076 588680 24078
rect -4756 24054 588680 24076
rect -4756 23818 -4574 24054
rect -4338 23818 22586 24054
rect 22822 23818 58586 24054
rect 58822 23818 94586 24054
rect 94822 23818 130586 24054
rect 130822 23818 166586 24054
rect 166822 23818 202586 24054
rect 202822 23818 238586 24054
rect 238822 23818 274586 24054
rect 274822 23818 310586 24054
rect 310822 23818 346586 24054
rect 346822 23818 382586 24054
rect 382822 23818 418586 24054
rect 418822 23818 454586 24054
rect 454822 23818 490586 24054
rect 490822 23818 526586 24054
rect 526822 23818 562586 24054
rect 562822 23818 588262 24054
rect 588498 23818 588680 24054
rect -4756 23734 588680 23818
rect -4756 23498 -4574 23734
rect -4338 23498 22586 23734
rect 22822 23498 58586 23734
rect 58822 23498 94586 23734
rect 94822 23498 130586 23734
rect 130822 23498 166586 23734
rect 166822 23498 202586 23734
rect 202822 23498 238586 23734
rect 238822 23498 274586 23734
rect 274822 23498 310586 23734
rect 310822 23498 346586 23734
rect 346822 23498 382586 23734
rect 382822 23498 418586 23734
rect 418822 23498 454586 23734
rect 454822 23498 490586 23734
rect 490822 23498 526586 23734
rect 526822 23498 562586 23734
rect 562822 23498 588262 23734
rect 588498 23498 588680 23734
rect -4756 23476 588680 23498
rect -4756 23474 -4156 23476
rect 22404 23474 23004 23476
rect 58404 23474 59004 23476
rect 94404 23474 95004 23476
rect 130404 23474 131004 23476
rect 166404 23474 167004 23476
rect 202404 23474 203004 23476
rect 238404 23474 239004 23476
rect 274404 23474 275004 23476
rect 310404 23474 311004 23476
rect 346404 23474 347004 23476
rect 382404 23474 383004 23476
rect 418404 23474 419004 23476
rect 454404 23474 455004 23476
rect 490404 23474 491004 23476
rect 526404 23474 527004 23476
rect 562404 23474 563004 23476
rect 588080 23474 588680 23476
rect -2916 20476 -2316 20478
rect 18804 20476 19404 20478
rect 54804 20476 55404 20478
rect 90804 20476 91404 20478
rect 126804 20476 127404 20478
rect 162804 20476 163404 20478
rect 198804 20476 199404 20478
rect 234804 20476 235404 20478
rect 270804 20476 271404 20478
rect 306804 20476 307404 20478
rect 342804 20476 343404 20478
rect 378804 20476 379404 20478
rect 414804 20476 415404 20478
rect 450804 20476 451404 20478
rect 486804 20476 487404 20478
rect 522804 20476 523404 20478
rect 558804 20476 559404 20478
rect 586240 20476 586840 20478
rect -2916 20454 586840 20476
rect -2916 20218 -2734 20454
rect -2498 20218 18986 20454
rect 19222 20218 54986 20454
rect 55222 20218 90986 20454
rect 91222 20218 126986 20454
rect 127222 20218 162986 20454
rect 163222 20218 198986 20454
rect 199222 20218 234986 20454
rect 235222 20218 270986 20454
rect 271222 20218 306986 20454
rect 307222 20218 342986 20454
rect 343222 20218 378986 20454
rect 379222 20218 414986 20454
rect 415222 20218 450986 20454
rect 451222 20218 486986 20454
rect 487222 20218 522986 20454
rect 523222 20218 558986 20454
rect 559222 20218 586422 20454
rect 586658 20218 586840 20454
rect -2916 20134 586840 20218
rect -2916 19898 -2734 20134
rect -2498 19898 18986 20134
rect 19222 19898 54986 20134
rect 55222 19898 90986 20134
rect 91222 19898 126986 20134
rect 127222 19898 162986 20134
rect 163222 19898 198986 20134
rect 199222 19898 234986 20134
rect 235222 19898 270986 20134
rect 271222 19898 306986 20134
rect 307222 19898 342986 20134
rect 343222 19898 378986 20134
rect 379222 19898 414986 20134
rect 415222 19898 450986 20134
rect 451222 19898 486986 20134
rect 487222 19898 522986 20134
rect 523222 19898 558986 20134
rect 559222 19898 586422 20134
rect 586658 19898 586840 20134
rect -2916 19876 586840 19898
rect -2916 19874 -2316 19876
rect 18804 19874 19404 19876
rect 54804 19874 55404 19876
rect 90804 19874 91404 19876
rect 126804 19874 127404 19876
rect 162804 19874 163404 19876
rect 198804 19874 199404 19876
rect 234804 19874 235404 19876
rect 270804 19874 271404 19876
rect 306804 19874 307404 19876
rect 342804 19874 343404 19876
rect 378804 19874 379404 19876
rect 414804 19874 415404 19876
rect 450804 19874 451404 19876
rect 486804 19874 487404 19876
rect 522804 19874 523404 19876
rect 558804 19874 559404 19876
rect 586240 19874 586840 19876
rect -7516 13276 -6916 13278
rect 11604 13276 12204 13278
rect 47604 13276 48204 13278
rect 83604 13276 84204 13278
rect 119604 13276 120204 13278
rect 155604 13276 156204 13278
rect 191604 13276 192204 13278
rect 227604 13276 228204 13278
rect 263604 13276 264204 13278
rect 299604 13276 300204 13278
rect 335604 13276 336204 13278
rect 371604 13276 372204 13278
rect 407604 13276 408204 13278
rect 443604 13276 444204 13278
rect 479604 13276 480204 13278
rect 515604 13276 516204 13278
rect 551604 13276 552204 13278
rect 590840 13276 591440 13278
rect -8436 13254 592360 13276
rect -8436 13018 -7334 13254
rect -7098 13018 11786 13254
rect 12022 13018 47786 13254
rect 48022 13018 83786 13254
rect 84022 13018 119786 13254
rect 120022 13018 155786 13254
rect 156022 13018 191786 13254
rect 192022 13018 227786 13254
rect 228022 13018 263786 13254
rect 264022 13018 299786 13254
rect 300022 13018 335786 13254
rect 336022 13018 371786 13254
rect 372022 13018 407786 13254
rect 408022 13018 443786 13254
rect 444022 13018 479786 13254
rect 480022 13018 515786 13254
rect 516022 13018 551786 13254
rect 552022 13018 591022 13254
rect 591258 13018 592360 13254
rect -8436 12934 592360 13018
rect -8436 12698 -7334 12934
rect -7098 12698 11786 12934
rect 12022 12698 47786 12934
rect 48022 12698 83786 12934
rect 84022 12698 119786 12934
rect 120022 12698 155786 12934
rect 156022 12698 191786 12934
rect 192022 12698 227786 12934
rect 228022 12698 263786 12934
rect 264022 12698 299786 12934
rect 300022 12698 335786 12934
rect 336022 12698 371786 12934
rect 372022 12698 407786 12934
rect 408022 12698 443786 12934
rect 444022 12698 479786 12934
rect 480022 12698 515786 12934
rect 516022 12698 551786 12934
rect 552022 12698 591022 12934
rect 591258 12698 592360 12934
rect -8436 12676 592360 12698
rect -7516 12674 -6916 12676
rect 11604 12674 12204 12676
rect 47604 12674 48204 12676
rect 83604 12674 84204 12676
rect 119604 12674 120204 12676
rect 155604 12674 156204 12676
rect 191604 12674 192204 12676
rect 227604 12674 228204 12676
rect 263604 12674 264204 12676
rect 299604 12674 300204 12676
rect 335604 12674 336204 12676
rect 371604 12674 372204 12676
rect 407604 12674 408204 12676
rect 443604 12674 444204 12676
rect 479604 12674 480204 12676
rect 515604 12674 516204 12676
rect 551604 12674 552204 12676
rect 590840 12674 591440 12676
rect -5676 9676 -5076 9678
rect 8004 9676 8604 9678
rect 44004 9676 44604 9678
rect 80004 9676 80604 9678
rect 116004 9676 116604 9678
rect 152004 9676 152604 9678
rect 188004 9676 188604 9678
rect 224004 9676 224604 9678
rect 260004 9676 260604 9678
rect 296004 9676 296604 9678
rect 332004 9676 332604 9678
rect 368004 9676 368604 9678
rect 404004 9676 404604 9678
rect 440004 9676 440604 9678
rect 476004 9676 476604 9678
rect 512004 9676 512604 9678
rect 548004 9676 548604 9678
rect 589000 9676 589600 9678
rect -6596 9654 590520 9676
rect -6596 9418 -5494 9654
rect -5258 9418 8186 9654
rect 8422 9418 44186 9654
rect 44422 9418 80186 9654
rect 80422 9418 116186 9654
rect 116422 9418 152186 9654
rect 152422 9418 188186 9654
rect 188422 9418 224186 9654
rect 224422 9418 260186 9654
rect 260422 9418 296186 9654
rect 296422 9418 332186 9654
rect 332422 9418 368186 9654
rect 368422 9418 404186 9654
rect 404422 9418 440186 9654
rect 440422 9418 476186 9654
rect 476422 9418 512186 9654
rect 512422 9418 548186 9654
rect 548422 9418 589182 9654
rect 589418 9418 590520 9654
rect -6596 9334 590520 9418
rect -6596 9098 -5494 9334
rect -5258 9098 8186 9334
rect 8422 9098 44186 9334
rect 44422 9098 80186 9334
rect 80422 9098 116186 9334
rect 116422 9098 152186 9334
rect 152422 9098 188186 9334
rect 188422 9098 224186 9334
rect 224422 9098 260186 9334
rect 260422 9098 296186 9334
rect 296422 9098 332186 9334
rect 332422 9098 368186 9334
rect 368422 9098 404186 9334
rect 404422 9098 440186 9334
rect 440422 9098 476186 9334
rect 476422 9098 512186 9334
rect 512422 9098 548186 9334
rect 548422 9098 589182 9334
rect 589418 9098 590520 9334
rect -6596 9076 590520 9098
rect -5676 9074 -5076 9076
rect 8004 9074 8604 9076
rect 44004 9074 44604 9076
rect 80004 9074 80604 9076
rect 116004 9074 116604 9076
rect 152004 9074 152604 9076
rect 188004 9074 188604 9076
rect 224004 9074 224604 9076
rect 260004 9074 260604 9076
rect 296004 9074 296604 9076
rect 332004 9074 332604 9076
rect 368004 9074 368604 9076
rect 404004 9074 404604 9076
rect 440004 9074 440604 9076
rect 476004 9074 476604 9076
rect 512004 9074 512604 9076
rect 548004 9074 548604 9076
rect 589000 9074 589600 9076
rect -3836 6076 -3236 6078
rect 4404 6076 5004 6078
rect 40404 6076 41004 6078
rect 76404 6076 77004 6078
rect 112404 6076 113004 6078
rect 148404 6076 149004 6078
rect 184404 6076 185004 6078
rect 220404 6076 221004 6078
rect 256404 6076 257004 6078
rect 292404 6076 293004 6078
rect 328404 6076 329004 6078
rect 364404 6076 365004 6078
rect 400404 6076 401004 6078
rect 436404 6076 437004 6078
rect 472404 6076 473004 6078
rect 508404 6076 509004 6078
rect 544404 6076 545004 6078
rect 580404 6076 581004 6078
rect 587160 6076 587760 6078
rect -4756 6054 588680 6076
rect -4756 5818 -3654 6054
rect -3418 5818 4586 6054
rect 4822 5818 40586 6054
rect 40822 5818 76586 6054
rect 76822 5818 112586 6054
rect 112822 5818 148586 6054
rect 148822 5818 184586 6054
rect 184822 5818 220586 6054
rect 220822 5818 256586 6054
rect 256822 5818 292586 6054
rect 292822 5818 328586 6054
rect 328822 5818 364586 6054
rect 364822 5818 400586 6054
rect 400822 5818 436586 6054
rect 436822 5818 472586 6054
rect 472822 5818 508586 6054
rect 508822 5818 544586 6054
rect 544822 5818 580586 6054
rect 580822 5818 587342 6054
rect 587578 5818 588680 6054
rect -4756 5734 588680 5818
rect -4756 5498 -3654 5734
rect -3418 5498 4586 5734
rect 4822 5498 40586 5734
rect 40822 5498 76586 5734
rect 76822 5498 112586 5734
rect 112822 5498 148586 5734
rect 148822 5498 184586 5734
rect 184822 5498 220586 5734
rect 220822 5498 256586 5734
rect 256822 5498 292586 5734
rect 292822 5498 328586 5734
rect 328822 5498 364586 5734
rect 364822 5498 400586 5734
rect 400822 5498 436586 5734
rect 436822 5498 472586 5734
rect 472822 5498 508586 5734
rect 508822 5498 544586 5734
rect 544822 5498 580586 5734
rect 580822 5498 587342 5734
rect 587578 5498 588680 5734
rect -4756 5476 588680 5498
rect -3836 5474 -3236 5476
rect 4404 5474 5004 5476
rect 40404 5474 41004 5476
rect 76404 5474 77004 5476
rect 112404 5474 113004 5476
rect 148404 5474 149004 5476
rect 184404 5474 185004 5476
rect 220404 5474 221004 5476
rect 256404 5474 257004 5476
rect 292404 5474 293004 5476
rect 328404 5474 329004 5476
rect 364404 5474 365004 5476
rect 400404 5474 401004 5476
rect 436404 5474 437004 5476
rect 472404 5474 473004 5476
rect 508404 5474 509004 5476
rect 544404 5474 545004 5476
rect 580404 5474 581004 5476
rect 587160 5474 587760 5476
rect -1996 2476 -1396 2478
rect 804 2476 1404 2478
rect 36804 2476 37404 2478
rect 72804 2476 73404 2478
rect 108804 2476 109404 2478
rect 144804 2476 145404 2478
rect 180804 2476 181404 2478
rect 216804 2476 217404 2478
rect 252804 2476 253404 2478
rect 288804 2476 289404 2478
rect 324804 2476 325404 2478
rect 360804 2476 361404 2478
rect 396804 2476 397404 2478
rect 432804 2476 433404 2478
rect 468804 2476 469404 2478
rect 504804 2476 505404 2478
rect 540804 2476 541404 2478
rect 576804 2476 577404 2478
rect 585320 2476 585920 2478
rect -2916 2454 586840 2476
rect -2916 2218 -1814 2454
rect -1578 2218 986 2454
rect 1222 2218 36986 2454
rect 37222 2218 72986 2454
rect 73222 2218 108986 2454
rect 109222 2218 144986 2454
rect 145222 2218 180986 2454
rect 181222 2218 216986 2454
rect 217222 2218 252986 2454
rect 253222 2218 288986 2454
rect 289222 2218 324986 2454
rect 325222 2218 360986 2454
rect 361222 2218 396986 2454
rect 397222 2218 432986 2454
rect 433222 2218 468986 2454
rect 469222 2218 504986 2454
rect 505222 2218 540986 2454
rect 541222 2218 576986 2454
rect 577222 2218 585502 2454
rect 585738 2218 586840 2454
rect -2916 2134 586840 2218
rect -2916 1898 -1814 2134
rect -1578 1898 986 2134
rect 1222 1898 36986 2134
rect 37222 1898 72986 2134
rect 73222 1898 108986 2134
rect 109222 1898 144986 2134
rect 145222 1898 180986 2134
rect 181222 1898 216986 2134
rect 217222 1898 252986 2134
rect 253222 1898 288986 2134
rect 289222 1898 324986 2134
rect 325222 1898 360986 2134
rect 361222 1898 396986 2134
rect 397222 1898 432986 2134
rect 433222 1898 468986 2134
rect 469222 1898 504986 2134
rect 505222 1898 540986 2134
rect 541222 1898 576986 2134
rect 577222 1898 585502 2134
rect 585738 1898 586840 2134
rect -2916 1876 586840 1898
rect -1996 1874 -1396 1876
rect 804 1874 1404 1876
rect 36804 1874 37404 1876
rect 72804 1874 73404 1876
rect 108804 1874 109404 1876
rect 144804 1874 145404 1876
rect 180804 1874 181404 1876
rect 216804 1874 217404 1876
rect 252804 1874 253404 1876
rect 288804 1874 289404 1876
rect 324804 1874 325404 1876
rect 360804 1874 361404 1876
rect 396804 1874 397404 1876
rect 432804 1874 433404 1876
rect 468804 1874 469404 1876
rect 504804 1874 505404 1876
rect 540804 1874 541404 1876
rect 576804 1874 577404 1876
rect 585320 1874 585920 1876
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 180804 -324 181404 -322
rect 216804 -324 217404 -322
rect 252804 -324 253404 -322
rect 288804 -324 289404 -322
rect 324804 -324 325404 -322
rect 360804 -324 361404 -322
rect 396804 -324 397404 -322
rect 432804 -324 433404 -322
rect 468804 -324 469404 -322
rect 504804 -324 505404 -322
rect 540804 -324 541404 -322
rect 576804 -324 577404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 180804 -926 181404 -924
rect 216804 -926 217404 -924
rect 252804 -926 253404 -924
rect 288804 -926 289404 -924
rect 324804 -926 325404 -924
rect 360804 -926 361404 -924
rect 396804 -926 397404 -924
rect 432804 -926 433404 -924
rect 468804 -926 469404 -924
rect 504804 -926 505404 -924
rect 540804 -926 541404 -924
rect 576804 -926 577404 -924
rect 585320 -926 585920 -924
rect -2916 -1244 -2316 -1242
rect 18804 -1244 19404 -1242
rect 54804 -1244 55404 -1242
rect 90804 -1244 91404 -1242
rect 126804 -1244 127404 -1242
rect 162804 -1244 163404 -1242
rect 198804 -1244 199404 -1242
rect 234804 -1244 235404 -1242
rect 270804 -1244 271404 -1242
rect 306804 -1244 307404 -1242
rect 342804 -1244 343404 -1242
rect 378804 -1244 379404 -1242
rect 414804 -1244 415404 -1242
rect 450804 -1244 451404 -1242
rect 486804 -1244 487404 -1242
rect 522804 -1244 523404 -1242
rect 558804 -1244 559404 -1242
rect 586240 -1244 586840 -1242
rect -2916 -1266 586840 -1244
rect -2916 -1502 -2734 -1266
rect -2498 -1502 18986 -1266
rect 19222 -1502 54986 -1266
rect 55222 -1502 90986 -1266
rect 91222 -1502 126986 -1266
rect 127222 -1502 162986 -1266
rect 163222 -1502 198986 -1266
rect 199222 -1502 234986 -1266
rect 235222 -1502 270986 -1266
rect 271222 -1502 306986 -1266
rect 307222 -1502 342986 -1266
rect 343222 -1502 378986 -1266
rect 379222 -1502 414986 -1266
rect 415222 -1502 450986 -1266
rect 451222 -1502 486986 -1266
rect 487222 -1502 522986 -1266
rect 523222 -1502 558986 -1266
rect 559222 -1502 586422 -1266
rect 586658 -1502 586840 -1266
rect -2916 -1586 586840 -1502
rect -2916 -1822 -2734 -1586
rect -2498 -1822 18986 -1586
rect 19222 -1822 54986 -1586
rect 55222 -1822 90986 -1586
rect 91222 -1822 126986 -1586
rect 127222 -1822 162986 -1586
rect 163222 -1822 198986 -1586
rect 199222 -1822 234986 -1586
rect 235222 -1822 270986 -1586
rect 271222 -1822 306986 -1586
rect 307222 -1822 342986 -1586
rect 343222 -1822 378986 -1586
rect 379222 -1822 414986 -1586
rect 415222 -1822 450986 -1586
rect 451222 -1822 486986 -1586
rect 487222 -1822 522986 -1586
rect 523222 -1822 558986 -1586
rect 559222 -1822 586422 -1586
rect 586658 -1822 586840 -1586
rect -2916 -1844 586840 -1822
rect -2916 -1846 -2316 -1844
rect 18804 -1846 19404 -1844
rect 54804 -1846 55404 -1844
rect 90804 -1846 91404 -1844
rect 126804 -1846 127404 -1844
rect 162804 -1846 163404 -1844
rect 198804 -1846 199404 -1844
rect 234804 -1846 235404 -1844
rect 270804 -1846 271404 -1844
rect 306804 -1846 307404 -1844
rect 342804 -1846 343404 -1844
rect 378804 -1846 379404 -1844
rect 414804 -1846 415404 -1844
rect 450804 -1846 451404 -1844
rect 486804 -1846 487404 -1844
rect 522804 -1846 523404 -1844
rect 558804 -1846 559404 -1844
rect 586240 -1846 586840 -1844
rect -3836 -2164 -3236 -2162
rect 4404 -2164 5004 -2162
rect 40404 -2164 41004 -2162
rect 76404 -2164 77004 -2162
rect 112404 -2164 113004 -2162
rect 148404 -2164 149004 -2162
rect 184404 -2164 185004 -2162
rect 220404 -2164 221004 -2162
rect 256404 -2164 257004 -2162
rect 292404 -2164 293004 -2162
rect 328404 -2164 329004 -2162
rect 364404 -2164 365004 -2162
rect 400404 -2164 401004 -2162
rect 436404 -2164 437004 -2162
rect 472404 -2164 473004 -2162
rect 508404 -2164 509004 -2162
rect 544404 -2164 545004 -2162
rect 580404 -2164 581004 -2162
rect 587160 -2164 587760 -2162
rect -3836 -2186 587760 -2164
rect -3836 -2422 -3654 -2186
rect -3418 -2422 4586 -2186
rect 4822 -2422 40586 -2186
rect 40822 -2422 76586 -2186
rect 76822 -2422 112586 -2186
rect 112822 -2422 148586 -2186
rect 148822 -2422 184586 -2186
rect 184822 -2422 220586 -2186
rect 220822 -2422 256586 -2186
rect 256822 -2422 292586 -2186
rect 292822 -2422 328586 -2186
rect 328822 -2422 364586 -2186
rect 364822 -2422 400586 -2186
rect 400822 -2422 436586 -2186
rect 436822 -2422 472586 -2186
rect 472822 -2422 508586 -2186
rect 508822 -2422 544586 -2186
rect 544822 -2422 580586 -2186
rect 580822 -2422 587342 -2186
rect 587578 -2422 587760 -2186
rect -3836 -2506 587760 -2422
rect -3836 -2742 -3654 -2506
rect -3418 -2742 4586 -2506
rect 4822 -2742 40586 -2506
rect 40822 -2742 76586 -2506
rect 76822 -2742 112586 -2506
rect 112822 -2742 148586 -2506
rect 148822 -2742 184586 -2506
rect 184822 -2742 220586 -2506
rect 220822 -2742 256586 -2506
rect 256822 -2742 292586 -2506
rect 292822 -2742 328586 -2506
rect 328822 -2742 364586 -2506
rect 364822 -2742 400586 -2506
rect 400822 -2742 436586 -2506
rect 436822 -2742 472586 -2506
rect 472822 -2742 508586 -2506
rect 508822 -2742 544586 -2506
rect 544822 -2742 580586 -2506
rect 580822 -2742 587342 -2506
rect 587578 -2742 587760 -2506
rect -3836 -2764 587760 -2742
rect -3836 -2766 -3236 -2764
rect 4404 -2766 5004 -2764
rect 40404 -2766 41004 -2764
rect 76404 -2766 77004 -2764
rect 112404 -2766 113004 -2764
rect 148404 -2766 149004 -2764
rect 184404 -2766 185004 -2764
rect 220404 -2766 221004 -2764
rect 256404 -2766 257004 -2764
rect 292404 -2766 293004 -2764
rect 328404 -2766 329004 -2764
rect 364404 -2766 365004 -2764
rect 400404 -2766 401004 -2764
rect 436404 -2766 437004 -2764
rect 472404 -2766 473004 -2764
rect 508404 -2766 509004 -2764
rect 544404 -2766 545004 -2764
rect 580404 -2766 581004 -2764
rect 587160 -2766 587760 -2764
rect -4756 -3084 -4156 -3082
rect 22404 -3084 23004 -3082
rect 58404 -3084 59004 -3082
rect 94404 -3084 95004 -3082
rect 130404 -3084 131004 -3082
rect 166404 -3084 167004 -3082
rect 202404 -3084 203004 -3082
rect 238404 -3084 239004 -3082
rect 274404 -3084 275004 -3082
rect 310404 -3084 311004 -3082
rect 346404 -3084 347004 -3082
rect 382404 -3084 383004 -3082
rect 418404 -3084 419004 -3082
rect 454404 -3084 455004 -3082
rect 490404 -3084 491004 -3082
rect 526404 -3084 527004 -3082
rect 562404 -3084 563004 -3082
rect 588080 -3084 588680 -3082
rect -4756 -3106 588680 -3084
rect -4756 -3342 -4574 -3106
rect -4338 -3342 22586 -3106
rect 22822 -3342 58586 -3106
rect 58822 -3342 94586 -3106
rect 94822 -3342 130586 -3106
rect 130822 -3342 166586 -3106
rect 166822 -3342 202586 -3106
rect 202822 -3342 238586 -3106
rect 238822 -3342 274586 -3106
rect 274822 -3342 310586 -3106
rect 310822 -3342 346586 -3106
rect 346822 -3342 382586 -3106
rect 382822 -3342 418586 -3106
rect 418822 -3342 454586 -3106
rect 454822 -3342 490586 -3106
rect 490822 -3342 526586 -3106
rect 526822 -3342 562586 -3106
rect 562822 -3342 588262 -3106
rect 588498 -3342 588680 -3106
rect -4756 -3426 588680 -3342
rect -4756 -3662 -4574 -3426
rect -4338 -3662 22586 -3426
rect 22822 -3662 58586 -3426
rect 58822 -3662 94586 -3426
rect 94822 -3662 130586 -3426
rect 130822 -3662 166586 -3426
rect 166822 -3662 202586 -3426
rect 202822 -3662 238586 -3426
rect 238822 -3662 274586 -3426
rect 274822 -3662 310586 -3426
rect 310822 -3662 346586 -3426
rect 346822 -3662 382586 -3426
rect 382822 -3662 418586 -3426
rect 418822 -3662 454586 -3426
rect 454822 -3662 490586 -3426
rect 490822 -3662 526586 -3426
rect 526822 -3662 562586 -3426
rect 562822 -3662 588262 -3426
rect 588498 -3662 588680 -3426
rect -4756 -3684 588680 -3662
rect -4756 -3686 -4156 -3684
rect 22404 -3686 23004 -3684
rect 58404 -3686 59004 -3684
rect 94404 -3686 95004 -3684
rect 130404 -3686 131004 -3684
rect 166404 -3686 167004 -3684
rect 202404 -3686 203004 -3684
rect 238404 -3686 239004 -3684
rect 274404 -3686 275004 -3684
rect 310404 -3686 311004 -3684
rect 346404 -3686 347004 -3684
rect 382404 -3686 383004 -3684
rect 418404 -3686 419004 -3684
rect 454404 -3686 455004 -3684
rect 490404 -3686 491004 -3684
rect 526404 -3686 527004 -3684
rect 562404 -3686 563004 -3684
rect 588080 -3686 588680 -3684
rect -5676 -4004 -5076 -4002
rect 8004 -4004 8604 -4002
rect 44004 -4004 44604 -4002
rect 80004 -4004 80604 -4002
rect 116004 -4004 116604 -4002
rect 152004 -4004 152604 -4002
rect 188004 -4004 188604 -4002
rect 224004 -4004 224604 -4002
rect 260004 -4004 260604 -4002
rect 296004 -4004 296604 -4002
rect 332004 -4004 332604 -4002
rect 368004 -4004 368604 -4002
rect 404004 -4004 404604 -4002
rect 440004 -4004 440604 -4002
rect 476004 -4004 476604 -4002
rect 512004 -4004 512604 -4002
rect 548004 -4004 548604 -4002
rect 589000 -4004 589600 -4002
rect -5676 -4026 589600 -4004
rect -5676 -4262 -5494 -4026
rect -5258 -4262 8186 -4026
rect 8422 -4262 44186 -4026
rect 44422 -4262 80186 -4026
rect 80422 -4262 116186 -4026
rect 116422 -4262 152186 -4026
rect 152422 -4262 188186 -4026
rect 188422 -4262 224186 -4026
rect 224422 -4262 260186 -4026
rect 260422 -4262 296186 -4026
rect 296422 -4262 332186 -4026
rect 332422 -4262 368186 -4026
rect 368422 -4262 404186 -4026
rect 404422 -4262 440186 -4026
rect 440422 -4262 476186 -4026
rect 476422 -4262 512186 -4026
rect 512422 -4262 548186 -4026
rect 548422 -4262 589182 -4026
rect 589418 -4262 589600 -4026
rect -5676 -4346 589600 -4262
rect -5676 -4582 -5494 -4346
rect -5258 -4582 8186 -4346
rect 8422 -4582 44186 -4346
rect 44422 -4582 80186 -4346
rect 80422 -4582 116186 -4346
rect 116422 -4582 152186 -4346
rect 152422 -4582 188186 -4346
rect 188422 -4582 224186 -4346
rect 224422 -4582 260186 -4346
rect 260422 -4582 296186 -4346
rect 296422 -4582 332186 -4346
rect 332422 -4582 368186 -4346
rect 368422 -4582 404186 -4346
rect 404422 -4582 440186 -4346
rect 440422 -4582 476186 -4346
rect 476422 -4582 512186 -4346
rect 512422 -4582 548186 -4346
rect 548422 -4582 589182 -4346
rect 589418 -4582 589600 -4346
rect -5676 -4604 589600 -4582
rect -5676 -4606 -5076 -4604
rect 8004 -4606 8604 -4604
rect 44004 -4606 44604 -4604
rect 80004 -4606 80604 -4604
rect 116004 -4606 116604 -4604
rect 152004 -4606 152604 -4604
rect 188004 -4606 188604 -4604
rect 224004 -4606 224604 -4604
rect 260004 -4606 260604 -4604
rect 296004 -4606 296604 -4604
rect 332004 -4606 332604 -4604
rect 368004 -4606 368604 -4604
rect 404004 -4606 404604 -4604
rect 440004 -4606 440604 -4604
rect 476004 -4606 476604 -4604
rect 512004 -4606 512604 -4604
rect 548004 -4606 548604 -4604
rect 589000 -4606 589600 -4604
rect -6596 -4924 -5996 -4922
rect 26004 -4924 26604 -4922
rect 62004 -4924 62604 -4922
rect 98004 -4924 98604 -4922
rect 134004 -4924 134604 -4922
rect 170004 -4924 170604 -4922
rect 206004 -4924 206604 -4922
rect 242004 -4924 242604 -4922
rect 278004 -4924 278604 -4922
rect 314004 -4924 314604 -4922
rect 350004 -4924 350604 -4922
rect 386004 -4924 386604 -4922
rect 422004 -4924 422604 -4922
rect 458004 -4924 458604 -4922
rect 494004 -4924 494604 -4922
rect 530004 -4924 530604 -4922
rect 566004 -4924 566604 -4922
rect 589920 -4924 590520 -4922
rect -6596 -4946 590520 -4924
rect -6596 -5182 -6414 -4946
rect -6178 -5182 26186 -4946
rect 26422 -5182 62186 -4946
rect 62422 -5182 98186 -4946
rect 98422 -5182 134186 -4946
rect 134422 -5182 170186 -4946
rect 170422 -5182 206186 -4946
rect 206422 -5182 242186 -4946
rect 242422 -5182 278186 -4946
rect 278422 -5182 314186 -4946
rect 314422 -5182 350186 -4946
rect 350422 -5182 386186 -4946
rect 386422 -5182 422186 -4946
rect 422422 -5182 458186 -4946
rect 458422 -5182 494186 -4946
rect 494422 -5182 530186 -4946
rect 530422 -5182 566186 -4946
rect 566422 -5182 590102 -4946
rect 590338 -5182 590520 -4946
rect -6596 -5266 590520 -5182
rect -6596 -5502 -6414 -5266
rect -6178 -5502 26186 -5266
rect 26422 -5502 62186 -5266
rect 62422 -5502 98186 -5266
rect 98422 -5502 134186 -5266
rect 134422 -5502 170186 -5266
rect 170422 -5502 206186 -5266
rect 206422 -5502 242186 -5266
rect 242422 -5502 278186 -5266
rect 278422 -5502 314186 -5266
rect 314422 -5502 350186 -5266
rect 350422 -5502 386186 -5266
rect 386422 -5502 422186 -5266
rect 422422 -5502 458186 -5266
rect 458422 -5502 494186 -5266
rect 494422 -5502 530186 -5266
rect 530422 -5502 566186 -5266
rect 566422 -5502 590102 -5266
rect 590338 -5502 590520 -5266
rect -6596 -5524 590520 -5502
rect -6596 -5526 -5996 -5524
rect 26004 -5526 26604 -5524
rect 62004 -5526 62604 -5524
rect 98004 -5526 98604 -5524
rect 134004 -5526 134604 -5524
rect 170004 -5526 170604 -5524
rect 206004 -5526 206604 -5524
rect 242004 -5526 242604 -5524
rect 278004 -5526 278604 -5524
rect 314004 -5526 314604 -5524
rect 350004 -5526 350604 -5524
rect 386004 -5526 386604 -5524
rect 422004 -5526 422604 -5524
rect 458004 -5526 458604 -5524
rect 494004 -5526 494604 -5524
rect 530004 -5526 530604 -5524
rect 566004 -5526 566604 -5524
rect 589920 -5526 590520 -5524
rect -7516 -5844 -6916 -5842
rect 11604 -5844 12204 -5842
rect 47604 -5844 48204 -5842
rect 83604 -5844 84204 -5842
rect 119604 -5844 120204 -5842
rect 155604 -5844 156204 -5842
rect 191604 -5844 192204 -5842
rect 227604 -5844 228204 -5842
rect 263604 -5844 264204 -5842
rect 299604 -5844 300204 -5842
rect 335604 -5844 336204 -5842
rect 371604 -5844 372204 -5842
rect 407604 -5844 408204 -5842
rect 443604 -5844 444204 -5842
rect 479604 -5844 480204 -5842
rect 515604 -5844 516204 -5842
rect 551604 -5844 552204 -5842
rect 590840 -5844 591440 -5842
rect -7516 -5866 591440 -5844
rect -7516 -6102 -7334 -5866
rect -7098 -6102 11786 -5866
rect 12022 -6102 47786 -5866
rect 48022 -6102 83786 -5866
rect 84022 -6102 119786 -5866
rect 120022 -6102 155786 -5866
rect 156022 -6102 191786 -5866
rect 192022 -6102 227786 -5866
rect 228022 -6102 263786 -5866
rect 264022 -6102 299786 -5866
rect 300022 -6102 335786 -5866
rect 336022 -6102 371786 -5866
rect 372022 -6102 407786 -5866
rect 408022 -6102 443786 -5866
rect 444022 -6102 479786 -5866
rect 480022 -6102 515786 -5866
rect 516022 -6102 551786 -5866
rect 552022 -6102 591022 -5866
rect 591258 -6102 591440 -5866
rect -7516 -6186 591440 -6102
rect -7516 -6422 -7334 -6186
rect -7098 -6422 11786 -6186
rect 12022 -6422 47786 -6186
rect 48022 -6422 83786 -6186
rect 84022 -6422 119786 -6186
rect 120022 -6422 155786 -6186
rect 156022 -6422 191786 -6186
rect 192022 -6422 227786 -6186
rect 228022 -6422 263786 -6186
rect 264022 -6422 299786 -6186
rect 300022 -6422 335786 -6186
rect 336022 -6422 371786 -6186
rect 372022 -6422 407786 -6186
rect 408022 -6422 443786 -6186
rect 444022 -6422 479786 -6186
rect 480022 -6422 515786 -6186
rect 516022 -6422 551786 -6186
rect 552022 -6422 591022 -6186
rect 591258 -6422 591440 -6186
rect -7516 -6444 591440 -6422
rect -7516 -6446 -6916 -6444
rect 11604 -6446 12204 -6444
rect 47604 -6446 48204 -6444
rect 83604 -6446 84204 -6444
rect 119604 -6446 120204 -6444
rect 155604 -6446 156204 -6444
rect 191604 -6446 192204 -6444
rect 227604 -6446 228204 -6444
rect 263604 -6446 264204 -6444
rect 299604 -6446 300204 -6444
rect 335604 -6446 336204 -6444
rect 371604 -6446 372204 -6444
rect 407604 -6446 408204 -6444
rect 443604 -6446 444204 -6444
rect 479604 -6446 480204 -6444
rect 515604 -6446 516204 -6444
rect 551604 -6446 552204 -6444
rect 590840 -6446 591440 -6444
rect -8436 -6764 -7836 -6762
rect 29604 -6764 30204 -6762
rect 65604 -6764 66204 -6762
rect 101604 -6764 102204 -6762
rect 137604 -6764 138204 -6762
rect 173604 -6764 174204 -6762
rect 209604 -6764 210204 -6762
rect 245604 -6764 246204 -6762
rect 281604 -6764 282204 -6762
rect 317604 -6764 318204 -6762
rect 353604 -6764 354204 -6762
rect 389604 -6764 390204 -6762
rect 425604 -6764 426204 -6762
rect 461604 -6764 462204 -6762
rect 497604 -6764 498204 -6762
rect 533604 -6764 534204 -6762
rect 569604 -6764 570204 -6762
rect 591760 -6764 592360 -6762
rect -8436 -6786 592360 -6764
rect -8436 -7022 -8254 -6786
rect -8018 -7022 29786 -6786
rect 30022 -7022 65786 -6786
rect 66022 -7022 101786 -6786
rect 102022 -7022 137786 -6786
rect 138022 -7022 173786 -6786
rect 174022 -7022 209786 -6786
rect 210022 -7022 245786 -6786
rect 246022 -7022 281786 -6786
rect 282022 -7022 317786 -6786
rect 318022 -7022 353786 -6786
rect 354022 -7022 389786 -6786
rect 390022 -7022 425786 -6786
rect 426022 -7022 461786 -6786
rect 462022 -7022 497786 -6786
rect 498022 -7022 533786 -6786
rect 534022 -7022 569786 -6786
rect 570022 -7022 591942 -6786
rect 592178 -7022 592360 -6786
rect -8436 -7106 592360 -7022
rect -8436 -7342 -8254 -7106
rect -8018 -7342 29786 -7106
rect 30022 -7342 65786 -7106
rect 66022 -7342 101786 -7106
rect 102022 -7342 137786 -7106
rect 138022 -7342 173786 -7106
rect 174022 -7342 209786 -7106
rect 210022 -7342 245786 -7106
rect 246022 -7342 281786 -7106
rect 282022 -7342 317786 -7106
rect 318022 -7342 353786 -7106
rect 354022 -7342 389786 -7106
rect 390022 -7342 425786 -7106
rect 426022 -7342 461786 -7106
rect 462022 -7342 497786 -7106
rect 498022 -7342 533786 -7106
rect 534022 -7342 569786 -7106
rect 570022 -7342 591942 -7106
rect 592178 -7342 592360 -7106
rect -8436 -7364 592360 -7342
rect -8436 -7366 -7836 -7364
rect 29604 -7366 30204 -7364
rect 65604 -7366 66204 -7364
rect 101604 -7366 102204 -7364
rect 137604 -7366 138204 -7364
rect 173604 -7366 174204 -7364
rect 209604 -7366 210204 -7364
rect 245604 -7366 246204 -7364
rect 281604 -7366 282204 -7364
rect 317604 -7366 318204 -7364
rect 353604 -7366 354204 -7364
rect 389604 -7366 390204 -7364
rect 425604 -7366 426204 -7364
rect 461604 -7366 462204 -7364
rect 497604 -7366 498204 -7364
rect 533604 -7366 534204 -7364
rect 569604 -7366 570204 -7364
rect 591760 -7366 592360 -7364
use user_proj_aes  mprj
timestamp 1607420573
transform 1 0 170000 0 1 220000
box 0 0 200000 300000
<< labels >>
rlabel metal3 s 583600 5796 584800 6036 6 analog_io[0]
port 0 nsew default bidirectional
rlabel metal3 s 583600 474996 584800 475236 6 analog_io[10]
port 1 nsew default bidirectional
rlabel metal3 s 583600 521916 584800 522156 6 analog_io[11]
port 2 nsew default bidirectional
rlabel metal3 s 583600 568836 584800 569076 6 analog_io[12]
port 3 nsew default bidirectional
rlabel metal3 s 583600 615756 584800 615996 6 analog_io[13]
port 4 nsew default bidirectional
rlabel metal3 s 583600 662676 584800 662916 6 analog_io[14]
port 5 nsew default bidirectional
rlabel metal2 s 575818 703600 575930 704800 6 analog_io[15]
port 6 nsew default bidirectional
rlabel metal2 s 510958 703600 511070 704800 6 analog_io[16]
port 7 nsew default bidirectional
rlabel metal2 s 446098 703600 446210 704800 6 analog_io[17]
port 8 nsew default bidirectional
rlabel metal2 s 381146 703600 381258 704800 6 analog_io[18]
port 9 nsew default bidirectional
rlabel metal2 s 316286 703600 316398 704800 6 analog_io[19]
port 10 nsew default bidirectional
rlabel metal3 s 583600 52716 584800 52956 6 analog_io[1]
port 11 nsew default bidirectional
rlabel metal2 s 251426 703600 251538 704800 6 analog_io[20]
port 12 nsew default bidirectional
rlabel metal2 s 186474 703600 186586 704800 6 analog_io[21]
port 13 nsew default bidirectional
rlabel metal2 s 121614 703600 121726 704800 6 analog_io[22]
port 14 nsew default bidirectional
rlabel metal2 s 56754 703600 56866 704800 6 analog_io[23]
port 15 nsew default bidirectional
rlabel metal3 s -800 696540 400 696780 4 analog_io[24]
port 16 nsew default bidirectional
rlabel metal3 s -800 639012 400 639252 4 analog_io[25]
port 17 nsew default bidirectional
rlabel metal3 s -800 581620 400 581860 4 analog_io[26]
port 18 nsew default bidirectional
rlabel metal3 s -800 524092 400 524332 4 analog_io[27]
port 19 nsew default bidirectional
rlabel metal3 s -800 466700 400 466940 4 analog_io[28]
port 20 nsew default bidirectional
rlabel metal3 s -800 409172 400 409412 4 analog_io[29]
port 21 nsew default bidirectional
rlabel metal3 s 583600 99636 584800 99876 6 analog_io[2]
port 22 nsew default bidirectional
rlabel metal3 s -800 351780 400 352020 4 analog_io[30]
port 23 nsew default bidirectional
rlabel metal3 s 583600 146556 584800 146796 6 analog_io[3]
port 24 nsew default bidirectional
rlabel metal3 s 583600 193476 584800 193716 6 analog_io[4]
port 25 nsew default bidirectional
rlabel metal3 s 583600 240396 584800 240636 6 analog_io[5]
port 26 nsew default bidirectional
rlabel metal3 s 583600 287316 584800 287556 6 analog_io[6]
port 27 nsew default bidirectional
rlabel metal3 s 583600 334236 584800 334476 6 analog_io[7]
port 28 nsew default bidirectional
rlabel metal3 s 583600 381156 584800 381396 6 analog_io[8]
port 29 nsew default bidirectional
rlabel metal3 s 583600 428076 584800 428316 6 analog_io[9]
port 30 nsew default bidirectional
rlabel metal3 s 583600 17492 584800 17732 6 io_in[0]
port 31 nsew default input
rlabel metal3 s 583600 486692 584800 486932 6 io_in[10]
port 32 nsew default input
rlabel metal3 s 583600 533748 584800 533988 6 io_in[11]
port 33 nsew default input
rlabel metal3 s 583600 580668 584800 580908 6 io_in[12]
port 34 nsew default input
rlabel metal3 s 583600 627588 584800 627828 6 io_in[13]
port 35 nsew default input
rlabel metal3 s 583600 674508 584800 674748 6 io_in[14]
port 36 nsew default input
rlabel metal2 s 559626 703600 559738 704800 6 io_in[15]
port 37 nsew default input
rlabel metal2 s 494766 703600 494878 704800 6 io_in[16]
port 38 nsew default input
rlabel metal2 s 429814 703600 429926 704800 6 io_in[17]
port 39 nsew default input
rlabel metal2 s 364954 703600 365066 704800 6 io_in[18]
port 40 nsew default input
rlabel metal2 s 300094 703600 300206 704800 6 io_in[19]
port 41 nsew default input
rlabel metal3 s 583600 64412 584800 64652 6 io_in[1]
port 42 nsew default input
rlabel metal2 s 235142 703600 235254 704800 6 io_in[20]
port 43 nsew default input
rlabel metal2 s 170282 703600 170394 704800 6 io_in[21]
port 44 nsew default input
rlabel metal2 s 105422 703600 105534 704800 6 io_in[22]
port 45 nsew default input
rlabel metal2 s 40470 703600 40582 704800 6 io_in[23]
port 46 nsew default input
rlabel metal3 s -800 682124 400 682364 4 io_in[24]
port 47 nsew default input
rlabel metal3 s -800 624732 400 624972 4 io_in[25]
port 48 nsew default input
rlabel metal3 s -800 567204 400 567444 4 io_in[26]
port 49 nsew default input
rlabel metal3 s -800 509812 400 510052 4 io_in[27]
port 50 nsew default input
rlabel metal3 s -800 452284 400 452524 4 io_in[28]
port 51 nsew default input
rlabel metal3 s -800 394892 400 395132 4 io_in[29]
port 52 nsew default input
rlabel metal3 s 583600 111332 584800 111572 6 io_in[2]
port 53 nsew default input
rlabel metal3 s -800 337364 400 337604 4 io_in[30]
port 54 nsew default input
rlabel metal3 s -800 294252 400 294492 4 io_in[31]
port 55 nsew default input
rlabel metal3 s -800 251140 400 251380 4 io_in[32]
port 56 nsew default input
rlabel metal3 s -800 208028 400 208268 4 io_in[33]
port 57 nsew default input
rlabel metal3 s -800 164916 400 165156 4 io_in[34]
port 58 nsew default input
rlabel metal3 s -800 121940 400 122180 4 io_in[35]
port 59 nsew default input
rlabel metal3 s -800 78828 400 79068 4 io_in[36]
port 60 nsew default input
rlabel metal3 s -800 35716 400 35956 4 io_in[37]
port 61 nsew default input
rlabel metal3 s 583600 158252 584800 158492 6 io_in[3]
port 62 nsew default input
rlabel metal3 s 583600 205172 584800 205412 6 io_in[4]
port 63 nsew default input
rlabel metal3 s 583600 252092 584800 252332 6 io_in[5]
port 64 nsew default input
rlabel metal3 s 583600 299012 584800 299252 6 io_in[6]
port 65 nsew default input
rlabel metal3 s 583600 345932 584800 346172 6 io_in[7]
port 66 nsew default input
rlabel metal3 s 583600 392852 584800 393092 6 io_in[8]
port 67 nsew default input
rlabel metal3 s 583600 439772 584800 440012 6 io_in[9]
port 68 nsew default input
rlabel metal3 s 583600 40884 584800 41124 6 io_oeb[0]
port 69 nsew default tristate
rlabel metal3 s 583600 510220 584800 510460 6 io_oeb[10]
port 70 nsew default tristate
rlabel metal3 s 583600 557140 584800 557380 6 io_oeb[11]
port 71 nsew default tristate
rlabel metal3 s 583600 604060 584800 604300 6 io_oeb[12]
port 72 nsew default tristate
rlabel metal3 s 583600 650980 584800 651220 6 io_oeb[13]
port 73 nsew default tristate
rlabel metal3 s 583600 697900 584800 698140 6 io_oeb[14]
port 74 nsew default tristate
rlabel metal2 s 527150 703600 527262 704800 6 io_oeb[15]
port 75 nsew default tristate
rlabel metal2 s 462290 703600 462402 704800 6 io_oeb[16]
port 76 nsew default tristate
rlabel metal2 s 397430 703600 397542 704800 6 io_oeb[17]
port 77 nsew default tristate
rlabel metal2 s 332478 703600 332590 704800 6 io_oeb[18]
port 78 nsew default tristate
rlabel metal2 s 267618 703600 267730 704800 6 io_oeb[19]
port 79 nsew default tristate
rlabel metal3 s 583600 87804 584800 88044 6 io_oeb[1]
port 80 nsew default tristate
rlabel metal2 s 202758 703600 202870 704800 6 io_oeb[20]
port 81 nsew default tristate
rlabel metal2 s 137806 703600 137918 704800 6 io_oeb[21]
port 82 nsew default tristate
rlabel metal2 s 72946 703600 73058 704800 6 io_oeb[22]
port 83 nsew default tristate
rlabel metal2 s 8086 703600 8198 704800 6 io_oeb[23]
port 84 nsew default tristate
rlabel metal3 s -800 653428 400 653668 4 io_oeb[24]
port 85 nsew default tristate
rlabel metal3 s -800 595900 400 596140 4 io_oeb[25]
port 86 nsew default tristate
rlabel metal3 s -800 538508 400 538748 4 io_oeb[26]
port 87 nsew default tristate
rlabel metal3 s -800 480980 400 481220 4 io_oeb[27]
port 88 nsew default tristate
rlabel metal3 s -800 423588 400 423828 4 io_oeb[28]
port 89 nsew default tristate
rlabel metal3 s -800 366060 400 366300 4 io_oeb[29]
port 90 nsew default tristate
rlabel metal3 s 583600 134724 584800 134964 6 io_oeb[2]
port 91 nsew default tristate
rlabel metal3 s -800 308668 400 308908 4 io_oeb[30]
port 92 nsew default tristate
rlabel metal3 s -800 265556 400 265796 4 io_oeb[31]
port 93 nsew default tristate
rlabel metal3 s -800 222444 400 222684 4 io_oeb[32]
port 94 nsew default tristate
rlabel metal3 s -800 179332 400 179572 4 io_oeb[33]
port 95 nsew default tristate
rlabel metal3 s -800 136220 400 136460 4 io_oeb[34]
port 96 nsew default tristate
rlabel metal3 s -800 93108 400 93348 4 io_oeb[35]
port 97 nsew default tristate
rlabel metal3 s -800 49996 400 50236 4 io_oeb[36]
port 98 nsew default tristate
rlabel metal3 s -800 7020 400 7260 4 io_oeb[37]
port 99 nsew default tristate
rlabel metal3 s 583600 181780 584800 182020 6 io_oeb[3]
port 100 nsew default tristate
rlabel metal3 s 583600 228700 584800 228940 6 io_oeb[4]
port 101 nsew default tristate
rlabel metal3 s 583600 275620 584800 275860 6 io_oeb[5]
port 102 nsew default tristate
rlabel metal3 s 583600 322540 584800 322780 6 io_oeb[6]
port 103 nsew default tristate
rlabel metal3 s 583600 369460 584800 369700 6 io_oeb[7]
port 104 nsew default tristate
rlabel metal3 s 583600 416380 584800 416620 6 io_oeb[8]
port 105 nsew default tristate
rlabel metal3 s 583600 463300 584800 463540 6 io_oeb[9]
port 106 nsew default tristate
rlabel metal3 s 583600 29188 584800 29428 6 io_out[0]
port 107 nsew default tristate
rlabel metal3 s 583600 498524 584800 498764 6 io_out[10]
port 108 nsew default tristate
rlabel metal3 s 583600 545444 584800 545684 6 io_out[11]
port 109 nsew default tristate
rlabel metal3 s 583600 592364 584800 592604 6 io_out[12]
port 110 nsew default tristate
rlabel metal3 s 583600 639284 584800 639524 6 io_out[13]
port 111 nsew default tristate
rlabel metal3 s 583600 686204 584800 686444 6 io_out[14]
port 112 nsew default tristate
rlabel metal2 s 543434 703600 543546 704800 6 io_out[15]
port 113 nsew default tristate
rlabel metal2 s 478482 703600 478594 704800 6 io_out[16]
port 114 nsew default tristate
rlabel metal2 s 413622 703600 413734 704800 6 io_out[17]
port 115 nsew default tristate
rlabel metal2 s 348762 703600 348874 704800 6 io_out[18]
port 116 nsew default tristate
rlabel metal2 s 283810 703600 283922 704800 6 io_out[19]
port 117 nsew default tristate
rlabel metal3 s 583600 76108 584800 76348 6 io_out[1]
port 118 nsew default tristate
rlabel metal2 s 218950 703600 219062 704800 6 io_out[20]
port 119 nsew default tristate
rlabel metal2 s 154090 703600 154202 704800 6 io_out[21]
port 120 nsew default tristate
rlabel metal2 s 89138 703600 89250 704800 6 io_out[22]
port 121 nsew default tristate
rlabel metal2 s 24278 703600 24390 704800 6 io_out[23]
port 122 nsew default tristate
rlabel metal3 s -800 667844 400 668084 4 io_out[24]
port 123 nsew default tristate
rlabel metal3 s -800 610316 400 610556 4 io_out[25]
port 124 nsew default tristate
rlabel metal3 s -800 552924 400 553164 4 io_out[26]
port 125 nsew default tristate
rlabel metal3 s -800 495396 400 495636 4 io_out[27]
port 126 nsew default tristate
rlabel metal3 s -800 437868 400 438108 4 io_out[28]
port 127 nsew default tristate
rlabel metal3 s -800 380476 400 380716 4 io_out[29]
port 128 nsew default tristate
rlabel metal3 s 583600 123028 584800 123268 6 io_out[2]
port 129 nsew default tristate
rlabel metal3 s -800 322948 400 323188 4 io_out[30]
port 130 nsew default tristate
rlabel metal3 s -800 279972 400 280212 4 io_out[31]
port 131 nsew default tristate
rlabel metal3 s -800 236860 400 237100 4 io_out[32]
port 132 nsew default tristate
rlabel metal3 s -800 193748 400 193988 4 io_out[33]
port 133 nsew default tristate
rlabel metal3 s -800 150636 400 150876 4 io_out[34]
port 134 nsew default tristate
rlabel metal3 s -800 107524 400 107764 4 io_out[35]
port 135 nsew default tristate
rlabel metal3 s -800 64412 400 64652 4 io_out[36]
port 136 nsew default tristate
rlabel metal3 s -800 21300 400 21540 4 io_out[37]
port 137 nsew default tristate
rlabel metal3 s 583600 169948 584800 170188 6 io_out[3]
port 138 nsew default tristate
rlabel metal3 s 583600 216868 584800 217108 6 io_out[4]
port 139 nsew default tristate
rlabel metal3 s 583600 263788 584800 264028 6 io_out[5]
port 140 nsew default tristate
rlabel metal3 s 583600 310708 584800 310948 6 io_out[6]
port 141 nsew default tristate
rlabel metal3 s 583600 357764 584800 358004 6 io_out[7]
port 142 nsew default tristate
rlabel metal3 s 583600 404684 584800 404924 6 io_out[8]
port 143 nsew default tristate
rlabel metal3 s 583600 451604 584800 451844 6 io_out[9]
port 144 nsew default tristate
rlabel metal2 s 126582 -800 126694 400 8 la_data_in[0]
port 145 nsew default input
rlabel metal2 s 483450 -800 483562 400 8 la_data_in[100]
port 146 nsew default input
rlabel metal2 s 486946 -800 487058 400 8 la_data_in[101]
port 147 nsew default input
rlabel metal2 s 490534 -800 490646 400 8 la_data_in[102]
port 148 nsew default input
rlabel metal2 s 494122 -800 494234 400 8 la_data_in[103]
port 149 nsew default input
rlabel metal2 s 497710 -800 497822 400 8 la_data_in[104]
port 150 nsew default input
rlabel metal2 s 501206 -800 501318 400 8 la_data_in[105]
port 151 nsew default input
rlabel metal2 s 504794 -800 504906 400 8 la_data_in[106]
port 152 nsew default input
rlabel metal2 s 508382 -800 508494 400 8 la_data_in[107]
port 153 nsew default input
rlabel metal2 s 511970 -800 512082 400 8 la_data_in[108]
port 154 nsew default input
rlabel metal2 s 515558 -800 515670 400 8 la_data_in[109]
port 155 nsew default input
rlabel metal2 s 162278 -800 162390 400 8 la_data_in[10]
port 156 nsew default input
rlabel metal2 s 519054 -800 519166 400 8 la_data_in[110]
port 157 nsew default input
rlabel metal2 s 522642 -800 522754 400 8 la_data_in[111]
port 158 nsew default input
rlabel metal2 s 526230 -800 526342 400 8 la_data_in[112]
port 159 nsew default input
rlabel metal2 s 529818 -800 529930 400 8 la_data_in[113]
port 160 nsew default input
rlabel metal2 s 533406 -800 533518 400 8 la_data_in[114]
port 161 nsew default input
rlabel metal2 s 536902 -800 537014 400 8 la_data_in[115]
port 162 nsew default input
rlabel metal2 s 540490 -800 540602 400 8 la_data_in[116]
port 163 nsew default input
rlabel metal2 s 544078 -800 544190 400 8 la_data_in[117]
port 164 nsew default input
rlabel metal2 s 547666 -800 547778 400 8 la_data_in[118]
port 165 nsew default input
rlabel metal2 s 551162 -800 551274 400 8 la_data_in[119]
port 166 nsew default input
rlabel metal2 s 165866 -800 165978 400 8 la_data_in[11]
port 167 nsew default input
rlabel metal2 s 554750 -800 554862 400 8 la_data_in[120]
port 168 nsew default input
rlabel metal2 s 558338 -800 558450 400 8 la_data_in[121]
port 169 nsew default input
rlabel metal2 s 561926 -800 562038 400 8 la_data_in[122]
port 170 nsew default input
rlabel metal2 s 565514 -800 565626 400 8 la_data_in[123]
port 171 nsew default input
rlabel metal2 s 569010 -800 569122 400 8 la_data_in[124]
port 172 nsew default input
rlabel metal2 s 572598 -800 572710 400 8 la_data_in[125]
port 173 nsew default input
rlabel metal2 s 576186 -800 576298 400 8 la_data_in[126]
port 174 nsew default input
rlabel metal2 s 579774 -800 579886 400 8 la_data_in[127]
port 175 nsew default input
rlabel metal2 s 169362 -800 169474 400 8 la_data_in[12]
port 176 nsew default input
rlabel metal2 s 172950 -800 173062 400 8 la_data_in[13]
port 177 nsew default input
rlabel metal2 s 176538 -800 176650 400 8 la_data_in[14]
port 178 nsew default input
rlabel metal2 s 180126 -800 180238 400 8 la_data_in[15]
port 179 nsew default input
rlabel metal2 s 183714 -800 183826 400 8 la_data_in[16]
port 180 nsew default input
rlabel metal2 s 187210 -800 187322 400 8 la_data_in[17]
port 181 nsew default input
rlabel metal2 s 190798 -800 190910 400 8 la_data_in[18]
port 182 nsew default input
rlabel metal2 s 194386 -800 194498 400 8 la_data_in[19]
port 183 nsew default input
rlabel metal2 s 130170 -800 130282 400 8 la_data_in[1]
port 184 nsew default input
rlabel metal2 s 197974 -800 198086 400 8 la_data_in[20]
port 185 nsew default input
rlabel metal2 s 201470 -800 201582 400 8 la_data_in[21]
port 186 nsew default input
rlabel metal2 s 205058 -800 205170 400 8 la_data_in[22]
port 187 nsew default input
rlabel metal2 s 208646 -800 208758 400 8 la_data_in[23]
port 188 nsew default input
rlabel metal2 s 212234 -800 212346 400 8 la_data_in[24]
port 189 nsew default input
rlabel metal2 s 215822 -800 215934 400 8 la_data_in[25]
port 190 nsew default input
rlabel metal2 s 219318 -800 219430 400 8 la_data_in[26]
port 191 nsew default input
rlabel metal2 s 222906 -800 223018 400 8 la_data_in[27]
port 192 nsew default input
rlabel metal2 s 226494 -800 226606 400 8 la_data_in[28]
port 193 nsew default input
rlabel metal2 s 230082 -800 230194 400 8 la_data_in[29]
port 194 nsew default input
rlabel metal2 s 133758 -800 133870 400 8 la_data_in[2]
port 195 nsew default input
rlabel metal2 s 233670 -800 233782 400 8 la_data_in[30]
port 196 nsew default input
rlabel metal2 s 237166 -800 237278 400 8 la_data_in[31]
port 197 nsew default input
rlabel metal2 s 240754 -800 240866 400 8 la_data_in[32]
port 198 nsew default input
rlabel metal2 s 244342 -800 244454 400 8 la_data_in[33]
port 199 nsew default input
rlabel metal2 s 247930 -800 248042 400 8 la_data_in[34]
port 200 nsew default input
rlabel metal2 s 251426 -800 251538 400 8 la_data_in[35]
port 201 nsew default input
rlabel metal2 s 255014 -800 255126 400 8 la_data_in[36]
port 202 nsew default input
rlabel metal2 s 258602 -800 258714 400 8 la_data_in[37]
port 203 nsew default input
rlabel metal2 s 262190 -800 262302 400 8 la_data_in[38]
port 204 nsew default input
rlabel metal2 s 265778 -800 265890 400 8 la_data_in[39]
port 205 nsew default input
rlabel metal2 s 137254 -800 137366 400 8 la_data_in[3]
port 206 nsew default input
rlabel metal2 s 269274 -800 269386 400 8 la_data_in[40]
port 207 nsew default input
rlabel metal2 s 272862 -800 272974 400 8 la_data_in[41]
port 208 nsew default input
rlabel metal2 s 276450 -800 276562 400 8 la_data_in[42]
port 209 nsew default input
rlabel metal2 s 280038 -800 280150 400 8 la_data_in[43]
port 210 nsew default input
rlabel metal2 s 283626 -800 283738 400 8 la_data_in[44]
port 211 nsew default input
rlabel metal2 s 287122 -800 287234 400 8 la_data_in[45]
port 212 nsew default input
rlabel metal2 s 290710 -800 290822 400 8 la_data_in[46]
port 213 nsew default input
rlabel metal2 s 294298 -800 294410 400 8 la_data_in[47]
port 214 nsew default input
rlabel metal2 s 297886 -800 297998 400 8 la_data_in[48]
port 215 nsew default input
rlabel metal2 s 301382 -800 301494 400 8 la_data_in[49]
port 216 nsew default input
rlabel metal2 s 140842 -800 140954 400 8 la_data_in[4]
port 217 nsew default input
rlabel metal2 s 304970 -800 305082 400 8 la_data_in[50]
port 218 nsew default input
rlabel metal2 s 308558 -800 308670 400 8 la_data_in[51]
port 219 nsew default input
rlabel metal2 s 312146 -800 312258 400 8 la_data_in[52]
port 220 nsew default input
rlabel metal2 s 315734 -800 315846 400 8 la_data_in[53]
port 221 nsew default input
rlabel metal2 s 319230 -800 319342 400 8 la_data_in[54]
port 222 nsew default input
rlabel metal2 s 322818 -800 322930 400 8 la_data_in[55]
port 223 nsew default input
rlabel metal2 s 326406 -800 326518 400 8 la_data_in[56]
port 224 nsew default input
rlabel metal2 s 329994 -800 330106 400 8 la_data_in[57]
port 225 nsew default input
rlabel metal2 s 333582 -800 333694 400 8 la_data_in[58]
port 226 nsew default input
rlabel metal2 s 337078 -800 337190 400 8 la_data_in[59]
port 227 nsew default input
rlabel metal2 s 144430 -800 144542 400 8 la_data_in[5]
port 228 nsew default input
rlabel metal2 s 340666 -800 340778 400 8 la_data_in[60]
port 229 nsew default input
rlabel metal2 s 344254 -800 344366 400 8 la_data_in[61]
port 230 nsew default input
rlabel metal2 s 347842 -800 347954 400 8 la_data_in[62]
port 231 nsew default input
rlabel metal2 s 351338 -800 351450 400 8 la_data_in[63]
port 232 nsew default input
rlabel metal2 s 354926 -800 355038 400 8 la_data_in[64]
port 233 nsew default input
rlabel metal2 s 358514 -800 358626 400 8 la_data_in[65]
port 234 nsew default input
rlabel metal2 s 362102 -800 362214 400 8 la_data_in[66]
port 235 nsew default input
rlabel metal2 s 365690 -800 365802 400 8 la_data_in[67]
port 236 nsew default input
rlabel metal2 s 369186 -800 369298 400 8 la_data_in[68]
port 237 nsew default input
rlabel metal2 s 372774 -800 372886 400 8 la_data_in[69]
port 238 nsew default input
rlabel metal2 s 148018 -800 148130 400 8 la_data_in[6]
port 239 nsew default input
rlabel metal2 s 376362 -800 376474 400 8 la_data_in[70]
port 240 nsew default input
rlabel metal2 s 379950 -800 380062 400 8 la_data_in[71]
port 241 nsew default input
rlabel metal2 s 383538 -800 383650 400 8 la_data_in[72]
port 242 nsew default input
rlabel metal2 s 387034 -800 387146 400 8 la_data_in[73]
port 243 nsew default input
rlabel metal2 s 390622 -800 390734 400 8 la_data_in[74]
port 244 nsew default input
rlabel metal2 s 394210 -800 394322 400 8 la_data_in[75]
port 245 nsew default input
rlabel metal2 s 397798 -800 397910 400 8 la_data_in[76]
port 246 nsew default input
rlabel metal2 s 401294 -800 401406 400 8 la_data_in[77]
port 247 nsew default input
rlabel metal2 s 404882 -800 404994 400 8 la_data_in[78]
port 248 nsew default input
rlabel metal2 s 408470 -800 408582 400 8 la_data_in[79]
port 249 nsew default input
rlabel metal2 s 151514 -800 151626 400 8 la_data_in[7]
port 250 nsew default input
rlabel metal2 s 412058 -800 412170 400 8 la_data_in[80]
port 251 nsew default input
rlabel metal2 s 415646 -800 415758 400 8 la_data_in[81]
port 252 nsew default input
rlabel metal2 s 419142 -800 419254 400 8 la_data_in[82]
port 253 nsew default input
rlabel metal2 s 422730 -800 422842 400 8 la_data_in[83]
port 254 nsew default input
rlabel metal2 s 426318 -800 426430 400 8 la_data_in[84]
port 255 nsew default input
rlabel metal2 s 429906 -800 430018 400 8 la_data_in[85]
port 256 nsew default input
rlabel metal2 s 433494 -800 433606 400 8 la_data_in[86]
port 257 nsew default input
rlabel metal2 s 436990 -800 437102 400 8 la_data_in[87]
port 258 nsew default input
rlabel metal2 s 440578 -800 440690 400 8 la_data_in[88]
port 259 nsew default input
rlabel metal2 s 444166 -800 444278 400 8 la_data_in[89]
port 260 nsew default input
rlabel metal2 s 155102 -800 155214 400 8 la_data_in[8]
port 261 nsew default input
rlabel metal2 s 447754 -800 447866 400 8 la_data_in[90]
port 262 nsew default input
rlabel metal2 s 451250 -800 451362 400 8 la_data_in[91]
port 263 nsew default input
rlabel metal2 s 454838 -800 454950 400 8 la_data_in[92]
port 264 nsew default input
rlabel metal2 s 458426 -800 458538 400 8 la_data_in[93]
port 265 nsew default input
rlabel metal2 s 462014 -800 462126 400 8 la_data_in[94]
port 266 nsew default input
rlabel metal2 s 465602 -800 465714 400 8 la_data_in[95]
port 267 nsew default input
rlabel metal2 s 469098 -800 469210 400 8 la_data_in[96]
port 268 nsew default input
rlabel metal2 s 472686 -800 472798 400 8 la_data_in[97]
port 269 nsew default input
rlabel metal2 s 476274 -800 476386 400 8 la_data_in[98]
port 270 nsew default input
rlabel metal2 s 479862 -800 479974 400 8 la_data_in[99]
port 271 nsew default input
rlabel metal2 s 158690 -800 158802 400 8 la_data_in[9]
port 272 nsew default input
rlabel metal2 s 127778 -800 127890 400 8 la_data_out[0]
port 273 nsew default tristate
rlabel metal2 s 484554 -800 484666 400 8 la_data_out[100]
port 274 nsew default tristate
rlabel metal2 s 488142 -800 488254 400 8 la_data_out[101]
port 275 nsew default tristate
rlabel metal2 s 491730 -800 491842 400 8 la_data_out[102]
port 276 nsew default tristate
rlabel metal2 s 495318 -800 495430 400 8 la_data_out[103]
port 277 nsew default tristate
rlabel metal2 s 498906 -800 499018 400 8 la_data_out[104]
port 278 nsew default tristate
rlabel metal2 s 502402 -800 502514 400 8 la_data_out[105]
port 279 nsew default tristate
rlabel metal2 s 505990 -800 506102 400 8 la_data_out[106]
port 280 nsew default tristate
rlabel metal2 s 509578 -800 509690 400 8 la_data_out[107]
port 281 nsew default tristate
rlabel metal2 s 513166 -800 513278 400 8 la_data_out[108]
port 282 nsew default tristate
rlabel metal2 s 516754 -800 516866 400 8 la_data_out[109]
port 283 nsew default tristate
rlabel metal2 s 163474 -800 163586 400 8 la_data_out[10]
port 284 nsew default tristate
rlabel metal2 s 520250 -800 520362 400 8 la_data_out[110]
port 285 nsew default tristate
rlabel metal2 s 523838 -800 523950 400 8 la_data_out[111]
port 286 nsew default tristate
rlabel metal2 s 527426 -800 527538 400 8 la_data_out[112]
port 287 nsew default tristate
rlabel metal2 s 531014 -800 531126 400 8 la_data_out[113]
port 288 nsew default tristate
rlabel metal2 s 534510 -800 534622 400 8 la_data_out[114]
port 289 nsew default tristate
rlabel metal2 s 538098 -800 538210 400 8 la_data_out[115]
port 290 nsew default tristate
rlabel metal2 s 541686 -800 541798 400 8 la_data_out[116]
port 291 nsew default tristate
rlabel metal2 s 545274 -800 545386 400 8 la_data_out[117]
port 292 nsew default tristate
rlabel metal2 s 548862 -800 548974 400 8 la_data_out[118]
port 293 nsew default tristate
rlabel metal2 s 552358 -800 552470 400 8 la_data_out[119]
port 294 nsew default tristate
rlabel metal2 s 167062 -800 167174 400 8 la_data_out[11]
port 295 nsew default tristate
rlabel metal2 s 555946 -800 556058 400 8 la_data_out[120]
port 296 nsew default tristate
rlabel metal2 s 559534 -800 559646 400 8 la_data_out[121]
port 297 nsew default tristate
rlabel metal2 s 563122 -800 563234 400 8 la_data_out[122]
port 298 nsew default tristate
rlabel metal2 s 566710 -800 566822 400 8 la_data_out[123]
port 299 nsew default tristate
rlabel metal2 s 570206 -800 570318 400 8 la_data_out[124]
port 300 nsew default tristate
rlabel metal2 s 573794 -800 573906 400 8 la_data_out[125]
port 301 nsew default tristate
rlabel metal2 s 577382 -800 577494 400 8 la_data_out[126]
port 302 nsew default tristate
rlabel metal2 s 580970 -800 581082 400 8 la_data_out[127]
port 303 nsew default tristate
rlabel metal2 s 170558 -800 170670 400 8 la_data_out[12]
port 304 nsew default tristate
rlabel metal2 s 174146 -800 174258 400 8 la_data_out[13]
port 305 nsew default tristate
rlabel metal2 s 177734 -800 177846 400 8 la_data_out[14]
port 306 nsew default tristate
rlabel metal2 s 181322 -800 181434 400 8 la_data_out[15]
port 307 nsew default tristate
rlabel metal2 s 184818 -800 184930 400 8 la_data_out[16]
port 308 nsew default tristate
rlabel metal2 s 188406 -800 188518 400 8 la_data_out[17]
port 309 nsew default tristate
rlabel metal2 s 191994 -800 192106 400 8 la_data_out[18]
port 310 nsew default tristate
rlabel metal2 s 195582 -800 195694 400 8 la_data_out[19]
port 311 nsew default tristate
rlabel metal2 s 131366 -800 131478 400 8 la_data_out[1]
port 312 nsew default tristate
rlabel metal2 s 199170 -800 199282 400 8 la_data_out[20]
port 313 nsew default tristate
rlabel metal2 s 202666 -800 202778 400 8 la_data_out[21]
port 314 nsew default tristate
rlabel metal2 s 206254 -800 206366 400 8 la_data_out[22]
port 315 nsew default tristate
rlabel metal2 s 209842 -800 209954 400 8 la_data_out[23]
port 316 nsew default tristate
rlabel metal2 s 213430 -800 213542 400 8 la_data_out[24]
port 317 nsew default tristate
rlabel metal2 s 217018 -800 217130 400 8 la_data_out[25]
port 318 nsew default tristate
rlabel metal2 s 220514 -800 220626 400 8 la_data_out[26]
port 319 nsew default tristate
rlabel metal2 s 224102 -800 224214 400 8 la_data_out[27]
port 320 nsew default tristate
rlabel metal2 s 227690 -800 227802 400 8 la_data_out[28]
port 321 nsew default tristate
rlabel metal2 s 231278 -800 231390 400 8 la_data_out[29]
port 322 nsew default tristate
rlabel metal2 s 134862 -800 134974 400 8 la_data_out[2]
port 323 nsew default tristate
rlabel metal2 s 234774 -800 234886 400 8 la_data_out[30]
port 324 nsew default tristate
rlabel metal2 s 238362 -800 238474 400 8 la_data_out[31]
port 325 nsew default tristate
rlabel metal2 s 241950 -800 242062 400 8 la_data_out[32]
port 326 nsew default tristate
rlabel metal2 s 245538 -800 245650 400 8 la_data_out[33]
port 327 nsew default tristate
rlabel metal2 s 249126 -800 249238 400 8 la_data_out[34]
port 328 nsew default tristate
rlabel metal2 s 252622 -800 252734 400 8 la_data_out[35]
port 329 nsew default tristate
rlabel metal2 s 256210 -800 256322 400 8 la_data_out[36]
port 330 nsew default tristate
rlabel metal2 s 259798 -800 259910 400 8 la_data_out[37]
port 331 nsew default tristate
rlabel metal2 s 263386 -800 263498 400 8 la_data_out[38]
port 332 nsew default tristate
rlabel metal2 s 266974 -800 267086 400 8 la_data_out[39]
port 333 nsew default tristate
rlabel metal2 s 138450 -800 138562 400 8 la_data_out[3]
port 334 nsew default tristate
rlabel metal2 s 270470 -800 270582 400 8 la_data_out[40]
port 335 nsew default tristate
rlabel metal2 s 274058 -800 274170 400 8 la_data_out[41]
port 336 nsew default tristate
rlabel metal2 s 277646 -800 277758 400 8 la_data_out[42]
port 337 nsew default tristate
rlabel metal2 s 281234 -800 281346 400 8 la_data_out[43]
port 338 nsew default tristate
rlabel metal2 s 284730 -800 284842 400 8 la_data_out[44]
port 339 nsew default tristate
rlabel metal2 s 288318 -800 288430 400 8 la_data_out[45]
port 340 nsew default tristate
rlabel metal2 s 291906 -800 292018 400 8 la_data_out[46]
port 341 nsew default tristate
rlabel metal2 s 295494 -800 295606 400 8 la_data_out[47]
port 342 nsew default tristate
rlabel metal2 s 299082 -800 299194 400 8 la_data_out[48]
port 343 nsew default tristate
rlabel metal2 s 302578 -800 302690 400 8 la_data_out[49]
port 344 nsew default tristate
rlabel metal2 s 142038 -800 142150 400 8 la_data_out[4]
port 345 nsew default tristate
rlabel metal2 s 306166 -800 306278 400 8 la_data_out[50]
port 346 nsew default tristate
rlabel metal2 s 309754 -800 309866 400 8 la_data_out[51]
port 347 nsew default tristate
rlabel metal2 s 313342 -800 313454 400 8 la_data_out[52]
port 348 nsew default tristate
rlabel metal2 s 316930 -800 317042 400 8 la_data_out[53]
port 349 nsew default tristate
rlabel metal2 s 320426 -800 320538 400 8 la_data_out[54]
port 350 nsew default tristate
rlabel metal2 s 324014 -800 324126 400 8 la_data_out[55]
port 351 nsew default tristate
rlabel metal2 s 327602 -800 327714 400 8 la_data_out[56]
port 352 nsew default tristate
rlabel metal2 s 331190 -800 331302 400 8 la_data_out[57]
port 353 nsew default tristate
rlabel metal2 s 334686 -800 334798 400 8 la_data_out[58]
port 354 nsew default tristate
rlabel metal2 s 338274 -800 338386 400 8 la_data_out[59]
port 355 nsew default tristate
rlabel metal2 s 145626 -800 145738 400 8 la_data_out[5]
port 356 nsew default tristate
rlabel metal2 s 341862 -800 341974 400 8 la_data_out[60]
port 357 nsew default tristate
rlabel metal2 s 345450 -800 345562 400 8 la_data_out[61]
port 358 nsew default tristate
rlabel metal2 s 349038 -800 349150 400 8 la_data_out[62]
port 359 nsew default tristate
rlabel metal2 s 352534 -800 352646 400 8 la_data_out[63]
port 360 nsew default tristate
rlabel metal2 s 356122 -800 356234 400 8 la_data_out[64]
port 361 nsew default tristate
rlabel metal2 s 359710 -800 359822 400 8 la_data_out[65]
port 362 nsew default tristate
rlabel metal2 s 363298 -800 363410 400 8 la_data_out[66]
port 363 nsew default tristate
rlabel metal2 s 366886 -800 366998 400 8 la_data_out[67]
port 364 nsew default tristate
rlabel metal2 s 370382 -800 370494 400 8 la_data_out[68]
port 365 nsew default tristate
rlabel metal2 s 373970 -800 374082 400 8 la_data_out[69]
port 366 nsew default tristate
rlabel metal2 s 149214 -800 149326 400 8 la_data_out[6]
port 367 nsew default tristate
rlabel metal2 s 377558 -800 377670 400 8 la_data_out[70]
port 368 nsew default tristate
rlabel metal2 s 381146 -800 381258 400 8 la_data_out[71]
port 369 nsew default tristate
rlabel metal2 s 384642 -800 384754 400 8 la_data_out[72]
port 370 nsew default tristate
rlabel metal2 s 388230 -800 388342 400 8 la_data_out[73]
port 371 nsew default tristate
rlabel metal2 s 391818 -800 391930 400 8 la_data_out[74]
port 372 nsew default tristate
rlabel metal2 s 395406 -800 395518 400 8 la_data_out[75]
port 373 nsew default tristate
rlabel metal2 s 398994 -800 399106 400 8 la_data_out[76]
port 374 nsew default tristate
rlabel metal2 s 402490 -800 402602 400 8 la_data_out[77]
port 375 nsew default tristate
rlabel metal2 s 406078 -800 406190 400 8 la_data_out[78]
port 376 nsew default tristate
rlabel metal2 s 409666 -800 409778 400 8 la_data_out[79]
port 377 nsew default tristate
rlabel metal2 s 152710 -800 152822 400 8 la_data_out[7]
port 378 nsew default tristate
rlabel metal2 s 413254 -800 413366 400 8 la_data_out[80]
port 379 nsew default tristate
rlabel metal2 s 416842 -800 416954 400 8 la_data_out[81]
port 380 nsew default tristate
rlabel metal2 s 420338 -800 420450 400 8 la_data_out[82]
port 381 nsew default tristate
rlabel metal2 s 423926 -800 424038 400 8 la_data_out[83]
port 382 nsew default tristate
rlabel metal2 s 427514 -800 427626 400 8 la_data_out[84]
port 383 nsew default tristate
rlabel metal2 s 431102 -800 431214 400 8 la_data_out[85]
port 384 nsew default tristate
rlabel metal2 s 434598 -800 434710 400 8 la_data_out[86]
port 385 nsew default tristate
rlabel metal2 s 438186 -800 438298 400 8 la_data_out[87]
port 386 nsew default tristate
rlabel metal2 s 441774 -800 441886 400 8 la_data_out[88]
port 387 nsew default tristate
rlabel metal2 s 445362 -800 445474 400 8 la_data_out[89]
port 388 nsew default tristate
rlabel metal2 s 156298 -800 156410 400 8 la_data_out[8]
port 389 nsew default tristate
rlabel metal2 s 448950 -800 449062 400 8 la_data_out[90]
port 390 nsew default tristate
rlabel metal2 s 452446 -800 452558 400 8 la_data_out[91]
port 391 nsew default tristate
rlabel metal2 s 456034 -800 456146 400 8 la_data_out[92]
port 392 nsew default tristate
rlabel metal2 s 459622 -800 459734 400 8 la_data_out[93]
port 393 nsew default tristate
rlabel metal2 s 463210 -800 463322 400 8 la_data_out[94]
port 394 nsew default tristate
rlabel metal2 s 466798 -800 466910 400 8 la_data_out[95]
port 395 nsew default tristate
rlabel metal2 s 470294 -800 470406 400 8 la_data_out[96]
port 396 nsew default tristate
rlabel metal2 s 473882 -800 473994 400 8 la_data_out[97]
port 397 nsew default tristate
rlabel metal2 s 477470 -800 477582 400 8 la_data_out[98]
port 398 nsew default tristate
rlabel metal2 s 481058 -800 481170 400 8 la_data_out[99]
port 399 nsew default tristate
rlabel metal2 s 159886 -800 159998 400 8 la_data_out[9]
port 400 nsew default tristate
rlabel metal2 s 128974 -800 129086 400 8 la_oen[0]
port 401 nsew default input
rlabel metal2 s 485750 -800 485862 400 8 la_oen[100]
port 402 nsew default input
rlabel metal2 s 489338 -800 489450 400 8 la_oen[101]
port 403 nsew default input
rlabel metal2 s 492926 -800 493038 400 8 la_oen[102]
port 404 nsew default input
rlabel metal2 s 496514 -800 496626 400 8 la_oen[103]
port 405 nsew default input
rlabel metal2 s 500102 -800 500214 400 8 la_oen[104]
port 406 nsew default input
rlabel metal2 s 503598 -800 503710 400 8 la_oen[105]
port 407 nsew default input
rlabel metal2 s 507186 -800 507298 400 8 la_oen[106]
port 408 nsew default input
rlabel metal2 s 510774 -800 510886 400 8 la_oen[107]
port 409 nsew default input
rlabel metal2 s 514362 -800 514474 400 8 la_oen[108]
port 410 nsew default input
rlabel metal2 s 517858 -800 517970 400 8 la_oen[109]
port 411 nsew default input
rlabel metal2 s 164670 -800 164782 400 8 la_oen[10]
port 412 nsew default input
rlabel metal2 s 521446 -800 521558 400 8 la_oen[110]
port 413 nsew default input
rlabel metal2 s 525034 -800 525146 400 8 la_oen[111]
port 414 nsew default input
rlabel metal2 s 528622 -800 528734 400 8 la_oen[112]
port 415 nsew default input
rlabel metal2 s 532210 -800 532322 400 8 la_oen[113]
port 416 nsew default input
rlabel metal2 s 535706 -800 535818 400 8 la_oen[114]
port 417 nsew default input
rlabel metal2 s 539294 -800 539406 400 8 la_oen[115]
port 418 nsew default input
rlabel metal2 s 542882 -800 542994 400 8 la_oen[116]
port 419 nsew default input
rlabel metal2 s 546470 -800 546582 400 8 la_oen[117]
port 420 nsew default input
rlabel metal2 s 550058 -800 550170 400 8 la_oen[118]
port 421 nsew default input
rlabel metal2 s 553554 -800 553666 400 8 la_oen[119]
port 422 nsew default input
rlabel metal2 s 168166 -800 168278 400 8 la_oen[11]
port 423 nsew default input
rlabel metal2 s 557142 -800 557254 400 8 la_oen[120]
port 424 nsew default input
rlabel metal2 s 560730 -800 560842 400 8 la_oen[121]
port 425 nsew default input
rlabel metal2 s 564318 -800 564430 400 8 la_oen[122]
port 426 nsew default input
rlabel metal2 s 567814 -800 567926 400 8 la_oen[123]
port 427 nsew default input
rlabel metal2 s 571402 -800 571514 400 8 la_oen[124]
port 428 nsew default input
rlabel metal2 s 574990 -800 575102 400 8 la_oen[125]
port 429 nsew default input
rlabel metal2 s 578578 -800 578690 400 8 la_oen[126]
port 430 nsew default input
rlabel metal2 s 582166 -800 582278 400 8 la_oen[127]
port 431 nsew default input
rlabel metal2 s 171754 -800 171866 400 8 la_oen[12]
port 432 nsew default input
rlabel metal2 s 175342 -800 175454 400 8 la_oen[13]
port 433 nsew default input
rlabel metal2 s 178930 -800 179042 400 8 la_oen[14]
port 434 nsew default input
rlabel metal2 s 182518 -800 182630 400 8 la_oen[15]
port 435 nsew default input
rlabel metal2 s 186014 -800 186126 400 8 la_oen[16]
port 436 nsew default input
rlabel metal2 s 189602 -800 189714 400 8 la_oen[17]
port 437 nsew default input
rlabel metal2 s 193190 -800 193302 400 8 la_oen[18]
port 438 nsew default input
rlabel metal2 s 196778 -800 196890 400 8 la_oen[19]
port 439 nsew default input
rlabel metal2 s 132562 -800 132674 400 8 la_oen[1]
port 440 nsew default input
rlabel metal2 s 200366 -800 200478 400 8 la_oen[20]
port 441 nsew default input
rlabel metal2 s 203862 -800 203974 400 8 la_oen[21]
port 442 nsew default input
rlabel metal2 s 207450 -800 207562 400 8 la_oen[22]
port 443 nsew default input
rlabel metal2 s 211038 -800 211150 400 8 la_oen[23]
port 444 nsew default input
rlabel metal2 s 214626 -800 214738 400 8 la_oen[24]
port 445 nsew default input
rlabel metal2 s 218122 -800 218234 400 8 la_oen[25]
port 446 nsew default input
rlabel metal2 s 221710 -800 221822 400 8 la_oen[26]
port 447 nsew default input
rlabel metal2 s 225298 -800 225410 400 8 la_oen[27]
port 448 nsew default input
rlabel metal2 s 228886 -800 228998 400 8 la_oen[28]
port 449 nsew default input
rlabel metal2 s 232474 -800 232586 400 8 la_oen[29]
port 450 nsew default input
rlabel metal2 s 136058 -800 136170 400 8 la_oen[2]
port 451 nsew default input
rlabel metal2 s 235970 -800 236082 400 8 la_oen[30]
port 452 nsew default input
rlabel metal2 s 239558 -800 239670 400 8 la_oen[31]
port 453 nsew default input
rlabel metal2 s 243146 -800 243258 400 8 la_oen[32]
port 454 nsew default input
rlabel metal2 s 246734 -800 246846 400 8 la_oen[33]
port 455 nsew default input
rlabel metal2 s 250322 -800 250434 400 8 la_oen[34]
port 456 nsew default input
rlabel metal2 s 253818 -800 253930 400 8 la_oen[35]
port 457 nsew default input
rlabel metal2 s 257406 -800 257518 400 8 la_oen[36]
port 458 nsew default input
rlabel metal2 s 260994 -800 261106 400 8 la_oen[37]
port 459 nsew default input
rlabel metal2 s 264582 -800 264694 400 8 la_oen[38]
port 460 nsew default input
rlabel metal2 s 268078 -800 268190 400 8 la_oen[39]
port 461 nsew default input
rlabel metal2 s 139646 -800 139758 400 8 la_oen[3]
port 462 nsew default input
rlabel metal2 s 271666 -800 271778 400 8 la_oen[40]
port 463 nsew default input
rlabel metal2 s 275254 -800 275366 400 8 la_oen[41]
port 464 nsew default input
rlabel metal2 s 278842 -800 278954 400 8 la_oen[42]
port 465 nsew default input
rlabel metal2 s 282430 -800 282542 400 8 la_oen[43]
port 466 nsew default input
rlabel metal2 s 285926 -800 286038 400 8 la_oen[44]
port 467 nsew default input
rlabel metal2 s 289514 -800 289626 400 8 la_oen[45]
port 468 nsew default input
rlabel metal2 s 293102 -800 293214 400 8 la_oen[46]
port 469 nsew default input
rlabel metal2 s 296690 -800 296802 400 8 la_oen[47]
port 470 nsew default input
rlabel metal2 s 300278 -800 300390 400 8 la_oen[48]
port 471 nsew default input
rlabel metal2 s 303774 -800 303886 400 8 la_oen[49]
port 472 nsew default input
rlabel metal2 s 143234 -800 143346 400 8 la_oen[4]
port 473 nsew default input
rlabel metal2 s 307362 -800 307474 400 8 la_oen[50]
port 474 nsew default input
rlabel metal2 s 310950 -800 311062 400 8 la_oen[51]
port 475 nsew default input
rlabel metal2 s 314538 -800 314650 400 8 la_oen[52]
port 476 nsew default input
rlabel metal2 s 318034 -800 318146 400 8 la_oen[53]
port 477 nsew default input
rlabel metal2 s 321622 -800 321734 400 8 la_oen[54]
port 478 nsew default input
rlabel metal2 s 325210 -800 325322 400 8 la_oen[55]
port 479 nsew default input
rlabel metal2 s 328798 -800 328910 400 8 la_oen[56]
port 480 nsew default input
rlabel metal2 s 332386 -800 332498 400 8 la_oen[57]
port 481 nsew default input
rlabel metal2 s 335882 -800 335994 400 8 la_oen[58]
port 482 nsew default input
rlabel metal2 s 339470 -800 339582 400 8 la_oen[59]
port 483 nsew default input
rlabel metal2 s 146822 -800 146934 400 8 la_oen[5]
port 484 nsew default input
rlabel metal2 s 343058 -800 343170 400 8 la_oen[60]
port 485 nsew default input
rlabel metal2 s 346646 -800 346758 400 8 la_oen[61]
port 486 nsew default input
rlabel metal2 s 350234 -800 350346 400 8 la_oen[62]
port 487 nsew default input
rlabel metal2 s 353730 -800 353842 400 8 la_oen[63]
port 488 nsew default input
rlabel metal2 s 357318 -800 357430 400 8 la_oen[64]
port 489 nsew default input
rlabel metal2 s 360906 -800 361018 400 8 la_oen[65]
port 490 nsew default input
rlabel metal2 s 364494 -800 364606 400 8 la_oen[66]
port 491 nsew default input
rlabel metal2 s 367990 -800 368102 400 8 la_oen[67]
port 492 nsew default input
rlabel metal2 s 371578 -800 371690 400 8 la_oen[68]
port 493 nsew default input
rlabel metal2 s 375166 -800 375278 400 8 la_oen[69]
port 494 nsew default input
rlabel metal2 s 150410 -800 150522 400 8 la_oen[6]
port 495 nsew default input
rlabel metal2 s 378754 -800 378866 400 8 la_oen[70]
port 496 nsew default input
rlabel metal2 s 382342 -800 382454 400 8 la_oen[71]
port 497 nsew default input
rlabel metal2 s 385838 -800 385950 400 8 la_oen[72]
port 498 nsew default input
rlabel metal2 s 389426 -800 389538 400 8 la_oen[73]
port 499 nsew default input
rlabel metal2 s 393014 -800 393126 400 8 la_oen[74]
port 500 nsew default input
rlabel metal2 s 396602 -800 396714 400 8 la_oen[75]
port 501 nsew default input
rlabel metal2 s 400190 -800 400302 400 8 la_oen[76]
port 502 nsew default input
rlabel metal2 s 403686 -800 403798 400 8 la_oen[77]
port 503 nsew default input
rlabel metal2 s 407274 -800 407386 400 8 la_oen[78]
port 504 nsew default input
rlabel metal2 s 410862 -800 410974 400 8 la_oen[79]
port 505 nsew default input
rlabel metal2 s 153906 -800 154018 400 8 la_oen[7]
port 506 nsew default input
rlabel metal2 s 414450 -800 414562 400 8 la_oen[80]
port 507 nsew default input
rlabel metal2 s 417946 -800 418058 400 8 la_oen[81]
port 508 nsew default input
rlabel metal2 s 421534 -800 421646 400 8 la_oen[82]
port 509 nsew default input
rlabel metal2 s 425122 -800 425234 400 8 la_oen[83]
port 510 nsew default input
rlabel metal2 s 428710 -800 428822 400 8 la_oen[84]
port 511 nsew default input
rlabel metal2 s 432298 -800 432410 400 8 la_oen[85]
port 512 nsew default input
rlabel metal2 s 435794 -800 435906 400 8 la_oen[86]
port 513 nsew default input
rlabel metal2 s 439382 -800 439494 400 8 la_oen[87]
port 514 nsew default input
rlabel metal2 s 442970 -800 443082 400 8 la_oen[88]
port 515 nsew default input
rlabel metal2 s 446558 -800 446670 400 8 la_oen[89]
port 516 nsew default input
rlabel metal2 s 157494 -800 157606 400 8 la_oen[8]
port 517 nsew default input
rlabel metal2 s 450146 -800 450258 400 8 la_oen[90]
port 518 nsew default input
rlabel metal2 s 453642 -800 453754 400 8 la_oen[91]
port 519 nsew default input
rlabel metal2 s 457230 -800 457342 400 8 la_oen[92]
port 520 nsew default input
rlabel metal2 s 460818 -800 460930 400 8 la_oen[93]
port 521 nsew default input
rlabel metal2 s 464406 -800 464518 400 8 la_oen[94]
port 522 nsew default input
rlabel metal2 s 467902 -800 468014 400 8 la_oen[95]
port 523 nsew default input
rlabel metal2 s 471490 -800 471602 400 8 la_oen[96]
port 524 nsew default input
rlabel metal2 s 475078 -800 475190 400 8 la_oen[97]
port 525 nsew default input
rlabel metal2 s 478666 -800 478778 400 8 la_oen[98]
port 526 nsew default input
rlabel metal2 s 482254 -800 482366 400 8 la_oen[99]
port 527 nsew default input
rlabel metal2 s 161082 -800 161194 400 8 la_oen[9]
port 528 nsew default input
rlabel metal2 s 583362 -800 583474 400 8 user_clock2
port 529 nsew default input
rlabel metal2 s 542 -800 654 400 8 wb_clk_i
port 530 nsew default input
rlabel metal2 s 1646 -800 1758 400 8 wb_rst_i
port 531 nsew default input
rlabel metal2 s 2842 -800 2954 400 8 wbs_ack_o
port 532 nsew default tristate
rlabel metal2 s 7626 -800 7738 400 8 wbs_adr_i[0]
port 533 nsew default input
rlabel metal2 s 48106 -800 48218 400 8 wbs_adr_i[10]
port 534 nsew default input
rlabel metal2 s 51602 -800 51714 400 8 wbs_adr_i[11]
port 535 nsew default input
rlabel metal2 s 55190 -800 55302 400 8 wbs_adr_i[12]
port 536 nsew default input
rlabel metal2 s 58778 -800 58890 400 8 wbs_adr_i[13]
port 537 nsew default input
rlabel metal2 s 62366 -800 62478 400 8 wbs_adr_i[14]
port 538 nsew default input
rlabel metal2 s 65954 -800 66066 400 8 wbs_adr_i[15]
port 539 nsew default input
rlabel metal2 s 69450 -800 69562 400 8 wbs_adr_i[16]
port 540 nsew default input
rlabel metal2 s 73038 -800 73150 400 8 wbs_adr_i[17]
port 541 nsew default input
rlabel metal2 s 76626 -800 76738 400 8 wbs_adr_i[18]
port 542 nsew default input
rlabel metal2 s 80214 -800 80326 400 8 wbs_adr_i[19]
port 543 nsew default input
rlabel metal2 s 12410 -800 12522 400 8 wbs_adr_i[1]
port 544 nsew default input
rlabel metal2 s 83802 -800 83914 400 8 wbs_adr_i[20]
port 545 nsew default input
rlabel metal2 s 87298 -800 87410 400 8 wbs_adr_i[21]
port 546 nsew default input
rlabel metal2 s 90886 -800 90998 400 8 wbs_adr_i[22]
port 547 nsew default input
rlabel metal2 s 94474 -800 94586 400 8 wbs_adr_i[23]
port 548 nsew default input
rlabel metal2 s 98062 -800 98174 400 8 wbs_adr_i[24]
port 549 nsew default input
rlabel metal2 s 101558 -800 101670 400 8 wbs_adr_i[25]
port 550 nsew default input
rlabel metal2 s 105146 -800 105258 400 8 wbs_adr_i[26]
port 551 nsew default input
rlabel metal2 s 108734 -800 108846 400 8 wbs_adr_i[27]
port 552 nsew default input
rlabel metal2 s 112322 -800 112434 400 8 wbs_adr_i[28]
port 553 nsew default input
rlabel metal2 s 115910 -800 116022 400 8 wbs_adr_i[29]
port 554 nsew default input
rlabel metal2 s 17194 -800 17306 400 8 wbs_adr_i[2]
port 555 nsew default input
rlabel metal2 s 119406 -800 119518 400 8 wbs_adr_i[30]
port 556 nsew default input
rlabel metal2 s 122994 -800 123106 400 8 wbs_adr_i[31]
port 557 nsew default input
rlabel metal2 s 21886 -800 21998 400 8 wbs_adr_i[3]
port 558 nsew default input
rlabel metal2 s 26670 -800 26782 400 8 wbs_adr_i[4]
port 559 nsew default input
rlabel metal2 s 30258 -800 30370 400 8 wbs_adr_i[5]
port 560 nsew default input
rlabel metal2 s 33846 -800 33958 400 8 wbs_adr_i[6]
port 561 nsew default input
rlabel metal2 s 37342 -800 37454 400 8 wbs_adr_i[7]
port 562 nsew default input
rlabel metal2 s 40930 -800 41042 400 8 wbs_adr_i[8]
port 563 nsew default input
rlabel metal2 s 44518 -800 44630 400 8 wbs_adr_i[9]
port 564 nsew default input
rlabel metal2 s 4038 -800 4150 400 8 wbs_cyc_i
port 565 nsew default input
rlabel metal2 s 8822 -800 8934 400 8 wbs_dat_i[0]
port 566 nsew default input
rlabel metal2 s 49302 -800 49414 400 8 wbs_dat_i[10]
port 567 nsew default input
rlabel metal2 s 52798 -800 52910 400 8 wbs_dat_i[11]
port 568 nsew default input
rlabel metal2 s 56386 -800 56498 400 8 wbs_dat_i[12]
port 569 nsew default input
rlabel metal2 s 59974 -800 60086 400 8 wbs_dat_i[13]
port 570 nsew default input
rlabel metal2 s 63562 -800 63674 400 8 wbs_dat_i[14]
port 571 nsew default input
rlabel metal2 s 67150 -800 67262 400 8 wbs_dat_i[15]
port 572 nsew default input
rlabel metal2 s 70646 -800 70758 400 8 wbs_dat_i[16]
port 573 nsew default input
rlabel metal2 s 74234 -800 74346 400 8 wbs_dat_i[17]
port 574 nsew default input
rlabel metal2 s 77822 -800 77934 400 8 wbs_dat_i[18]
port 575 nsew default input
rlabel metal2 s 81410 -800 81522 400 8 wbs_dat_i[19]
port 576 nsew default input
rlabel metal2 s 13606 -800 13718 400 8 wbs_dat_i[1]
port 577 nsew default input
rlabel metal2 s 84906 -800 85018 400 8 wbs_dat_i[20]
port 578 nsew default input
rlabel metal2 s 88494 -800 88606 400 8 wbs_dat_i[21]
port 579 nsew default input
rlabel metal2 s 92082 -800 92194 400 8 wbs_dat_i[22]
port 580 nsew default input
rlabel metal2 s 95670 -800 95782 400 8 wbs_dat_i[23]
port 581 nsew default input
rlabel metal2 s 99258 -800 99370 400 8 wbs_dat_i[24]
port 582 nsew default input
rlabel metal2 s 102754 -800 102866 400 8 wbs_dat_i[25]
port 583 nsew default input
rlabel metal2 s 106342 -800 106454 400 8 wbs_dat_i[26]
port 584 nsew default input
rlabel metal2 s 109930 -800 110042 400 8 wbs_dat_i[27]
port 585 nsew default input
rlabel metal2 s 113518 -800 113630 400 8 wbs_dat_i[28]
port 586 nsew default input
rlabel metal2 s 117106 -800 117218 400 8 wbs_dat_i[29]
port 587 nsew default input
rlabel metal2 s 18298 -800 18410 400 8 wbs_dat_i[2]
port 588 nsew default input
rlabel metal2 s 120602 -800 120714 400 8 wbs_dat_i[30]
port 589 nsew default input
rlabel metal2 s 124190 -800 124302 400 8 wbs_dat_i[31]
port 590 nsew default input
rlabel metal2 s 23082 -800 23194 400 8 wbs_dat_i[3]
port 591 nsew default input
rlabel metal2 s 27866 -800 27978 400 8 wbs_dat_i[4]
port 592 nsew default input
rlabel metal2 s 31454 -800 31566 400 8 wbs_dat_i[5]
port 593 nsew default input
rlabel metal2 s 34950 -800 35062 400 8 wbs_dat_i[6]
port 594 nsew default input
rlabel metal2 s 38538 -800 38650 400 8 wbs_dat_i[7]
port 595 nsew default input
rlabel metal2 s 42126 -800 42238 400 8 wbs_dat_i[8]
port 596 nsew default input
rlabel metal2 s 45714 -800 45826 400 8 wbs_dat_i[9]
port 597 nsew default input
rlabel metal2 s 10018 -800 10130 400 8 wbs_dat_o[0]
port 598 nsew default tristate
rlabel metal2 s 50498 -800 50610 400 8 wbs_dat_o[10]
port 599 nsew default tristate
rlabel metal2 s 53994 -800 54106 400 8 wbs_dat_o[11]
port 600 nsew default tristate
rlabel metal2 s 57582 -800 57694 400 8 wbs_dat_o[12]
port 601 nsew default tristate
rlabel metal2 s 61170 -800 61282 400 8 wbs_dat_o[13]
port 602 nsew default tristate
rlabel metal2 s 64758 -800 64870 400 8 wbs_dat_o[14]
port 603 nsew default tristate
rlabel metal2 s 68254 -800 68366 400 8 wbs_dat_o[15]
port 604 nsew default tristate
rlabel metal2 s 71842 -800 71954 400 8 wbs_dat_o[16]
port 605 nsew default tristate
rlabel metal2 s 75430 -800 75542 400 8 wbs_dat_o[17]
port 606 nsew default tristate
rlabel metal2 s 79018 -800 79130 400 8 wbs_dat_o[18]
port 607 nsew default tristate
rlabel metal2 s 82606 -800 82718 400 8 wbs_dat_o[19]
port 608 nsew default tristate
rlabel metal2 s 14802 -800 14914 400 8 wbs_dat_o[1]
port 609 nsew default tristate
rlabel metal2 s 86102 -800 86214 400 8 wbs_dat_o[20]
port 610 nsew default tristate
rlabel metal2 s 89690 -800 89802 400 8 wbs_dat_o[21]
port 611 nsew default tristate
rlabel metal2 s 93278 -800 93390 400 8 wbs_dat_o[22]
port 612 nsew default tristate
rlabel metal2 s 96866 -800 96978 400 8 wbs_dat_o[23]
port 613 nsew default tristate
rlabel metal2 s 100454 -800 100566 400 8 wbs_dat_o[24]
port 614 nsew default tristate
rlabel metal2 s 103950 -800 104062 400 8 wbs_dat_o[25]
port 615 nsew default tristate
rlabel metal2 s 107538 -800 107650 400 8 wbs_dat_o[26]
port 616 nsew default tristate
rlabel metal2 s 111126 -800 111238 400 8 wbs_dat_o[27]
port 617 nsew default tristate
rlabel metal2 s 114714 -800 114826 400 8 wbs_dat_o[28]
port 618 nsew default tristate
rlabel metal2 s 118210 -800 118322 400 8 wbs_dat_o[29]
port 619 nsew default tristate
rlabel metal2 s 19494 -800 19606 400 8 wbs_dat_o[2]
port 620 nsew default tristate
rlabel metal2 s 121798 -800 121910 400 8 wbs_dat_o[30]
port 621 nsew default tristate
rlabel metal2 s 125386 -800 125498 400 8 wbs_dat_o[31]
port 622 nsew default tristate
rlabel metal2 s 24278 -800 24390 400 8 wbs_dat_o[3]
port 623 nsew default tristate
rlabel metal2 s 29062 -800 29174 400 8 wbs_dat_o[4]
port 624 nsew default tristate
rlabel metal2 s 32650 -800 32762 400 8 wbs_dat_o[5]
port 625 nsew default tristate
rlabel metal2 s 36146 -800 36258 400 8 wbs_dat_o[6]
port 626 nsew default tristate
rlabel metal2 s 39734 -800 39846 400 8 wbs_dat_o[7]
port 627 nsew default tristate
rlabel metal2 s 43322 -800 43434 400 8 wbs_dat_o[8]
port 628 nsew default tristate
rlabel metal2 s 46910 -800 47022 400 8 wbs_dat_o[9]
port 629 nsew default tristate
rlabel metal2 s 11214 -800 11326 400 8 wbs_sel_i[0]
port 630 nsew default input
rlabel metal2 s 15998 -800 16110 400 8 wbs_sel_i[1]
port 631 nsew default input
rlabel metal2 s 20690 -800 20802 400 8 wbs_sel_i[2]
port 632 nsew default input
rlabel metal2 s 25474 -800 25586 400 8 wbs_sel_i[3]
port 633 nsew default input
rlabel metal2 s 5234 -800 5346 400 8 wbs_stb_i
port 634 nsew default input
rlabel metal2 s 6430 -800 6542 400 8 wbs_we_i
port 635 nsew default input
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 636 nsew default input
rlabel metal5 s -2916 -1844 586840 -1244 8 vssd1
port 637 nsew default input
rlabel metal5 s -3836 -2764 587760 -2164 8 vccd2
port 638 nsew default input
rlabel metal5 s -4756 -3684 588680 -3084 8 vssd2
port 639 nsew default input
rlabel metal5 s -5676 -4604 589600 -4004 8 vdda1
port 640 nsew default input
rlabel metal5 s -6596 -5524 590520 -4924 8 vssa1
port 641 nsew default input
rlabel metal5 s -7516 -6444 591440 -5844 8 vdda2
port 642 nsew default input
rlabel metal5 s -8436 -7364 592360 -6764 8 vssa2
port 643 nsew default input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
